magic
tech sky130A
magscale 1 2
timestamp 1679151745
<< nwell >>
rect -1410 6040 5250 10790
<< pwell >>
rect -5213 8647 -2017 11585
rect 6517 8647 9713 11585
rect 1191 4501 2631 5921
rect 1191 2981 2631 4401
rect 200 1460 3630 2880
rect -60 -60 3886 1360
<< nmos >>
rect 1387 4711 1487 5711
rect 1545 4711 1645 5711
rect 1703 4711 1803 5711
rect 1861 4711 1961 5711
rect 2019 4711 2119 5711
rect 2177 4711 2277 5711
rect 2335 4711 2435 5711
rect 1387 3191 1487 4191
rect 1545 3191 1645 4191
rect 1703 3191 1803 4191
rect 1861 3191 1961 4191
rect 2019 3191 2119 4191
rect 2177 3191 2277 4191
rect 2335 3191 2435 4191
rect 396 1670 596 2670
rect 654 1670 854 2670
rect 912 1670 1112 2670
rect 1170 1670 1370 2670
rect 1428 1670 1628 2670
rect 1686 1670 1886 2670
rect 1944 1670 2144 2670
rect 2202 1670 2402 2670
rect 2460 1670 2660 2670
rect 2718 1670 2918 2670
rect 2976 1670 3176 2670
rect 3234 1670 3434 2670
rect 136 150 336 1150
rect 394 150 594 1150
rect 652 150 852 1150
rect 910 150 1110 1150
rect 1168 150 1368 1150
rect 1426 150 1626 1150
rect 1684 150 1884 1150
rect 1942 150 2142 1150
rect 2200 150 2400 1150
rect 2458 150 2658 1150
rect 2716 150 2916 1150
rect 2974 150 3174 1150
rect 3232 150 3432 1150
rect 3490 150 3690 1150
<< pmos >>
rect -1214 9489 -1114 10489
rect -1056 9489 -956 10489
rect -898 9489 -798 10489
rect -740 9489 -640 10489
rect -582 9489 -482 10489
rect -424 9489 -324 10489
rect -266 9489 -166 10489
rect -108 9489 -8 10489
rect 50 9489 150 10489
rect 208 9489 308 10489
rect 366 9489 466 10489
rect 524 9489 624 10489
rect 682 9489 782 10489
rect 840 9489 940 10489
rect 998 9489 1098 10489
rect 1156 9489 1256 10489
rect 1314 9489 1414 10489
rect 1472 9489 1572 10489
rect 1630 9489 1730 10489
rect 1788 9489 1888 10489
rect 1946 9489 2046 10489
rect 2104 9489 2204 10489
rect 2262 9489 2362 10489
rect 2420 9489 2520 10489
rect 2578 9489 2678 10489
rect 2736 9489 2836 10489
rect 2894 9489 2994 10489
rect 3052 9489 3152 10489
rect 3210 9489 3310 10489
rect 3368 9489 3468 10489
rect 3526 9489 3626 10489
rect 3684 9489 3784 10489
rect 3842 9489 3942 10489
rect 4000 9489 4100 10489
rect 4158 9489 4258 10489
rect 4316 9489 4416 10489
rect 4474 9489 4574 10489
rect 4632 9489 4732 10489
rect 4790 9489 4890 10489
rect 4948 9489 5048 10489
rect 286 7819 386 8819
rect 444 7819 544 8819
rect 602 7819 702 8819
rect 760 7819 860 8819
rect 918 7819 1018 8819
rect 1076 7819 1176 8819
rect 1234 7819 1334 8819
rect 1392 7819 1492 8819
rect 1550 7819 1650 8819
rect 1708 7819 1808 8819
rect 1866 7819 1966 8819
rect 2024 7819 2124 8819
rect 2182 7819 2282 8819
rect 2340 7819 2440 8819
rect 2498 7819 2598 8819
rect 2656 7819 2756 8819
rect 2814 7819 2914 8819
rect 2972 7819 3072 8819
rect 3130 7819 3230 8819
rect 3288 7819 3388 8819
rect 3446 7819 3546 8819
rect 286 6279 386 7279
rect 444 6279 544 7279
rect 602 6279 702 7279
rect 760 6279 860 7279
rect 918 6279 1018 7279
rect 1076 6279 1176 7279
rect 1234 6279 1334 7279
rect 1392 6279 1492 7279
rect 1550 6279 1650 7279
rect 1708 6279 1808 7279
rect 1866 6279 1966 7279
rect 2024 6279 2124 7279
rect 2182 6279 2282 7279
rect 2340 6279 2440 7279
rect 2498 6279 2598 7279
rect 2656 6279 2756 7279
rect 2814 6279 2914 7279
rect 2972 6279 3072 7279
rect 3130 6279 3230 7279
rect 3288 6279 3388 7279
rect 3446 6279 3546 7279
<< ndiff >>
rect 1329 5699 1387 5711
rect 1329 4723 1341 5699
rect 1375 4723 1387 5699
rect 1329 4711 1387 4723
rect 1487 5699 1545 5711
rect 1487 4723 1499 5699
rect 1533 4723 1545 5699
rect 1487 4711 1545 4723
rect 1645 5699 1703 5711
rect 1645 4723 1657 5699
rect 1691 4723 1703 5699
rect 1645 4711 1703 4723
rect 1803 5699 1861 5711
rect 1803 4723 1815 5699
rect 1849 4723 1861 5699
rect 1803 4711 1861 4723
rect 1961 5699 2019 5711
rect 1961 4723 1973 5699
rect 2007 4723 2019 5699
rect 1961 4711 2019 4723
rect 2119 5699 2177 5711
rect 2119 4723 2131 5699
rect 2165 4723 2177 5699
rect 2119 4711 2177 4723
rect 2277 5699 2335 5711
rect 2277 4723 2289 5699
rect 2323 4723 2335 5699
rect 2277 4711 2335 4723
rect 2435 5699 2493 5711
rect 2435 4723 2447 5699
rect 2481 4723 2493 5699
rect 2435 4711 2493 4723
rect 1329 4179 1387 4191
rect 1329 3203 1341 4179
rect 1375 3203 1387 4179
rect 1329 3191 1387 3203
rect 1487 4179 1545 4191
rect 1487 3203 1499 4179
rect 1533 3203 1545 4179
rect 1487 3191 1545 3203
rect 1645 4179 1703 4191
rect 1645 3203 1657 4179
rect 1691 3203 1703 4179
rect 1645 3191 1703 3203
rect 1803 4179 1861 4191
rect 1803 3203 1815 4179
rect 1849 3203 1861 4179
rect 1803 3191 1861 3203
rect 1961 4179 2019 4191
rect 1961 3203 1973 4179
rect 2007 3203 2019 4179
rect 1961 3191 2019 3203
rect 2119 4179 2177 4191
rect 2119 3203 2131 4179
rect 2165 3203 2177 4179
rect 2119 3191 2177 3203
rect 2277 4179 2335 4191
rect 2277 3203 2289 4179
rect 2323 3203 2335 4179
rect 2277 3191 2335 3203
rect 2435 4179 2493 4191
rect 2435 3203 2447 4179
rect 2481 3203 2493 4179
rect 2435 3191 2493 3203
rect 338 2658 396 2670
rect 338 1682 350 2658
rect 384 1682 396 2658
rect 338 1670 396 1682
rect 596 2658 654 2670
rect 596 1682 608 2658
rect 642 1682 654 2658
rect 596 1670 654 1682
rect 854 2658 912 2670
rect 854 1682 866 2658
rect 900 1682 912 2658
rect 854 1670 912 1682
rect 1112 2658 1170 2670
rect 1112 1682 1124 2658
rect 1158 1682 1170 2658
rect 1112 1670 1170 1682
rect 1370 2658 1428 2670
rect 1370 1682 1382 2658
rect 1416 1682 1428 2658
rect 1370 1670 1428 1682
rect 1628 2658 1686 2670
rect 1628 1682 1640 2658
rect 1674 1682 1686 2658
rect 1628 1670 1686 1682
rect 1886 2658 1944 2670
rect 1886 1682 1898 2658
rect 1932 1682 1944 2658
rect 1886 1670 1944 1682
rect 2144 2658 2202 2670
rect 2144 1682 2156 2658
rect 2190 1682 2202 2658
rect 2144 1670 2202 1682
rect 2402 2658 2460 2670
rect 2402 1682 2414 2658
rect 2448 1682 2460 2658
rect 2402 1670 2460 1682
rect 2660 2658 2718 2670
rect 2660 1682 2672 2658
rect 2706 1682 2718 2658
rect 2660 1670 2718 1682
rect 2918 2658 2976 2670
rect 2918 1682 2930 2658
rect 2964 1682 2976 2658
rect 2918 1670 2976 1682
rect 3176 2658 3234 2670
rect 3176 1682 3188 2658
rect 3222 1682 3234 2658
rect 3176 1670 3234 1682
rect 3434 2658 3492 2670
rect 3434 1682 3446 2658
rect 3480 1682 3492 2658
rect 3434 1670 3492 1682
rect 78 1138 136 1150
rect 78 162 90 1138
rect 124 162 136 1138
rect 78 150 136 162
rect 336 1138 394 1150
rect 336 162 348 1138
rect 382 162 394 1138
rect 336 150 394 162
rect 594 1138 652 1150
rect 594 162 606 1138
rect 640 162 652 1138
rect 594 150 652 162
rect 852 1138 910 1150
rect 852 162 864 1138
rect 898 162 910 1138
rect 852 150 910 162
rect 1110 1138 1168 1150
rect 1110 162 1122 1138
rect 1156 162 1168 1138
rect 1110 150 1168 162
rect 1368 1138 1426 1150
rect 1368 162 1380 1138
rect 1414 162 1426 1138
rect 1368 150 1426 162
rect 1626 1138 1684 1150
rect 1626 162 1638 1138
rect 1672 162 1684 1138
rect 1626 150 1684 162
rect 1884 1138 1942 1150
rect 1884 162 1896 1138
rect 1930 162 1942 1138
rect 1884 150 1942 162
rect 2142 1138 2200 1150
rect 2142 162 2154 1138
rect 2188 162 2200 1138
rect 2142 150 2200 162
rect 2400 1138 2458 1150
rect 2400 162 2412 1138
rect 2446 162 2458 1138
rect 2400 150 2458 162
rect 2658 1138 2716 1150
rect 2658 162 2670 1138
rect 2704 162 2716 1138
rect 2658 150 2716 162
rect 2916 1138 2974 1150
rect 2916 162 2928 1138
rect 2962 162 2974 1138
rect 2916 150 2974 162
rect 3174 1138 3232 1150
rect 3174 162 3186 1138
rect 3220 162 3232 1138
rect 3174 150 3232 162
rect 3432 1138 3490 1150
rect 3432 162 3444 1138
rect 3478 162 3490 1138
rect 3432 150 3490 162
rect 3690 1138 3748 1150
rect 3690 162 3702 1138
rect 3736 162 3748 1138
rect 3690 150 3748 162
<< pdiff >>
rect -1272 10477 -1214 10489
rect -1272 9501 -1260 10477
rect -1226 9501 -1214 10477
rect -1272 9489 -1214 9501
rect -1114 10477 -1056 10489
rect -1114 9501 -1102 10477
rect -1068 9501 -1056 10477
rect -1114 9489 -1056 9501
rect -956 10477 -898 10489
rect -956 9501 -944 10477
rect -910 9501 -898 10477
rect -956 9489 -898 9501
rect -798 10477 -740 10489
rect -798 9501 -786 10477
rect -752 9501 -740 10477
rect -798 9489 -740 9501
rect -640 10477 -582 10489
rect -640 9501 -628 10477
rect -594 9501 -582 10477
rect -640 9489 -582 9501
rect -482 10477 -424 10489
rect -482 9501 -470 10477
rect -436 9501 -424 10477
rect -482 9489 -424 9501
rect -324 10477 -266 10489
rect -324 9501 -312 10477
rect -278 9501 -266 10477
rect -324 9489 -266 9501
rect -166 10477 -108 10489
rect -166 9501 -154 10477
rect -120 9501 -108 10477
rect -166 9489 -108 9501
rect -8 10477 50 10489
rect -8 9501 4 10477
rect 38 9501 50 10477
rect -8 9489 50 9501
rect 150 10477 208 10489
rect 150 9501 162 10477
rect 196 9501 208 10477
rect 150 9489 208 9501
rect 308 10477 366 10489
rect 308 9501 320 10477
rect 354 9501 366 10477
rect 308 9489 366 9501
rect 466 10477 524 10489
rect 466 9501 478 10477
rect 512 9501 524 10477
rect 466 9489 524 9501
rect 624 10477 682 10489
rect 624 9501 636 10477
rect 670 9501 682 10477
rect 624 9489 682 9501
rect 782 10477 840 10489
rect 782 9501 794 10477
rect 828 9501 840 10477
rect 782 9489 840 9501
rect 940 10477 998 10489
rect 940 9501 952 10477
rect 986 9501 998 10477
rect 940 9489 998 9501
rect 1098 10477 1156 10489
rect 1098 9501 1110 10477
rect 1144 9501 1156 10477
rect 1098 9489 1156 9501
rect 1256 10477 1314 10489
rect 1256 9501 1268 10477
rect 1302 9501 1314 10477
rect 1256 9489 1314 9501
rect 1414 10477 1472 10489
rect 1414 9501 1426 10477
rect 1460 9501 1472 10477
rect 1414 9489 1472 9501
rect 1572 10477 1630 10489
rect 1572 9501 1584 10477
rect 1618 9501 1630 10477
rect 1572 9489 1630 9501
rect 1730 10477 1788 10489
rect 1730 9501 1742 10477
rect 1776 9501 1788 10477
rect 1730 9489 1788 9501
rect 1888 10477 1946 10489
rect 1888 9501 1900 10477
rect 1934 9501 1946 10477
rect 1888 9489 1946 9501
rect 2046 10477 2104 10489
rect 2046 9501 2058 10477
rect 2092 9501 2104 10477
rect 2046 9489 2104 9501
rect 2204 10477 2262 10489
rect 2204 9501 2216 10477
rect 2250 9501 2262 10477
rect 2204 9489 2262 9501
rect 2362 10477 2420 10489
rect 2362 9501 2374 10477
rect 2408 9501 2420 10477
rect 2362 9489 2420 9501
rect 2520 10477 2578 10489
rect 2520 9501 2532 10477
rect 2566 9501 2578 10477
rect 2520 9489 2578 9501
rect 2678 10477 2736 10489
rect 2678 9501 2690 10477
rect 2724 9501 2736 10477
rect 2678 9489 2736 9501
rect 2836 10477 2894 10489
rect 2836 9501 2848 10477
rect 2882 9501 2894 10477
rect 2836 9489 2894 9501
rect 2994 10477 3052 10489
rect 2994 9501 3006 10477
rect 3040 9501 3052 10477
rect 2994 9489 3052 9501
rect 3152 10477 3210 10489
rect 3152 9501 3164 10477
rect 3198 9501 3210 10477
rect 3152 9489 3210 9501
rect 3310 10477 3368 10489
rect 3310 9501 3322 10477
rect 3356 9501 3368 10477
rect 3310 9489 3368 9501
rect 3468 10477 3526 10489
rect 3468 9501 3480 10477
rect 3514 9501 3526 10477
rect 3468 9489 3526 9501
rect 3626 10477 3684 10489
rect 3626 9501 3638 10477
rect 3672 9501 3684 10477
rect 3626 9489 3684 9501
rect 3784 10477 3842 10489
rect 3784 9501 3796 10477
rect 3830 9501 3842 10477
rect 3784 9489 3842 9501
rect 3942 10477 4000 10489
rect 3942 9501 3954 10477
rect 3988 9501 4000 10477
rect 3942 9489 4000 9501
rect 4100 10477 4158 10489
rect 4100 9501 4112 10477
rect 4146 9501 4158 10477
rect 4100 9489 4158 9501
rect 4258 10477 4316 10489
rect 4258 9501 4270 10477
rect 4304 9501 4316 10477
rect 4258 9489 4316 9501
rect 4416 10477 4474 10489
rect 4416 9501 4428 10477
rect 4462 9501 4474 10477
rect 4416 9489 4474 9501
rect 4574 10477 4632 10489
rect 4574 9501 4586 10477
rect 4620 9501 4632 10477
rect 4574 9489 4632 9501
rect 4732 10477 4790 10489
rect 4732 9501 4744 10477
rect 4778 9501 4790 10477
rect 4732 9489 4790 9501
rect 4890 10477 4948 10489
rect 4890 9501 4902 10477
rect 4936 9501 4948 10477
rect 4890 9489 4948 9501
rect 5048 10477 5106 10489
rect 5048 9501 5060 10477
rect 5094 9501 5106 10477
rect 5048 9489 5106 9501
rect 228 8807 286 8819
rect 228 7831 240 8807
rect 274 7831 286 8807
rect 228 7819 286 7831
rect 386 8807 444 8819
rect 386 7831 398 8807
rect 432 7831 444 8807
rect 386 7819 444 7831
rect 544 8807 602 8819
rect 544 7831 556 8807
rect 590 7831 602 8807
rect 544 7819 602 7831
rect 702 8807 760 8819
rect 702 7831 714 8807
rect 748 7831 760 8807
rect 702 7819 760 7831
rect 860 8807 918 8819
rect 860 7831 872 8807
rect 906 7831 918 8807
rect 860 7819 918 7831
rect 1018 8807 1076 8819
rect 1018 7831 1030 8807
rect 1064 7831 1076 8807
rect 1018 7819 1076 7831
rect 1176 8807 1234 8819
rect 1176 7831 1188 8807
rect 1222 7831 1234 8807
rect 1176 7819 1234 7831
rect 1334 8807 1392 8819
rect 1334 7831 1346 8807
rect 1380 7831 1392 8807
rect 1334 7819 1392 7831
rect 1492 8807 1550 8819
rect 1492 7831 1504 8807
rect 1538 7831 1550 8807
rect 1492 7819 1550 7831
rect 1650 8807 1708 8819
rect 1650 7831 1662 8807
rect 1696 7831 1708 8807
rect 1650 7819 1708 7831
rect 1808 8807 1866 8819
rect 1808 7831 1820 8807
rect 1854 7831 1866 8807
rect 1808 7819 1866 7831
rect 1966 8807 2024 8819
rect 1966 7831 1978 8807
rect 2012 7831 2024 8807
rect 1966 7819 2024 7831
rect 2124 8807 2182 8819
rect 2124 7831 2136 8807
rect 2170 7831 2182 8807
rect 2124 7819 2182 7831
rect 2282 8807 2340 8819
rect 2282 7831 2294 8807
rect 2328 7831 2340 8807
rect 2282 7819 2340 7831
rect 2440 8807 2498 8819
rect 2440 7831 2452 8807
rect 2486 7831 2498 8807
rect 2440 7819 2498 7831
rect 2598 8807 2656 8819
rect 2598 7831 2610 8807
rect 2644 7831 2656 8807
rect 2598 7819 2656 7831
rect 2756 8807 2814 8819
rect 2756 7831 2768 8807
rect 2802 7831 2814 8807
rect 2756 7819 2814 7831
rect 2914 8807 2972 8819
rect 2914 7831 2926 8807
rect 2960 7831 2972 8807
rect 2914 7819 2972 7831
rect 3072 8807 3130 8819
rect 3072 7831 3084 8807
rect 3118 7831 3130 8807
rect 3072 7819 3130 7831
rect 3230 8807 3288 8819
rect 3230 7831 3242 8807
rect 3276 7831 3288 8807
rect 3230 7819 3288 7831
rect 3388 8807 3446 8819
rect 3388 7831 3400 8807
rect 3434 7831 3446 8807
rect 3388 7819 3446 7831
rect 3546 8807 3604 8819
rect 3546 7831 3558 8807
rect 3592 7831 3604 8807
rect 3546 7819 3604 7831
rect 228 7267 286 7279
rect 228 6291 240 7267
rect 274 6291 286 7267
rect 228 6279 286 6291
rect 386 7267 444 7279
rect 386 6291 398 7267
rect 432 6291 444 7267
rect 386 6279 444 6291
rect 544 7267 602 7279
rect 544 6291 556 7267
rect 590 6291 602 7267
rect 544 6279 602 6291
rect 702 7267 760 7279
rect 702 6291 714 7267
rect 748 6291 760 7267
rect 702 6279 760 6291
rect 860 7267 918 7279
rect 860 6291 872 7267
rect 906 6291 918 7267
rect 860 6279 918 6291
rect 1018 7267 1076 7279
rect 1018 6291 1030 7267
rect 1064 6291 1076 7267
rect 1018 6279 1076 6291
rect 1176 7267 1234 7279
rect 1176 6291 1188 7267
rect 1222 6291 1234 7267
rect 1176 6279 1234 6291
rect 1334 7267 1392 7279
rect 1334 6291 1346 7267
rect 1380 6291 1392 7267
rect 1334 6279 1392 6291
rect 1492 7267 1550 7279
rect 1492 6291 1504 7267
rect 1538 6291 1550 7267
rect 1492 6279 1550 6291
rect 1650 7267 1708 7279
rect 1650 6291 1662 7267
rect 1696 6291 1708 7267
rect 1650 6279 1708 6291
rect 1808 7267 1866 7279
rect 1808 6291 1820 7267
rect 1854 6291 1866 7267
rect 1808 6279 1866 6291
rect 1966 7267 2024 7279
rect 1966 6291 1978 7267
rect 2012 6291 2024 7267
rect 1966 6279 2024 6291
rect 2124 7267 2182 7279
rect 2124 6291 2136 7267
rect 2170 6291 2182 7267
rect 2124 6279 2182 6291
rect 2282 7267 2340 7279
rect 2282 6291 2294 7267
rect 2328 6291 2340 7267
rect 2282 6279 2340 6291
rect 2440 7267 2498 7279
rect 2440 6291 2452 7267
rect 2486 6291 2498 7267
rect 2440 6279 2498 6291
rect 2598 7267 2656 7279
rect 2598 6291 2610 7267
rect 2644 6291 2656 7267
rect 2598 6279 2656 6291
rect 2756 7267 2814 7279
rect 2756 6291 2768 7267
rect 2802 6291 2814 7267
rect 2756 6279 2814 6291
rect 2914 7267 2972 7279
rect 2914 6291 2926 7267
rect 2960 6291 2972 7267
rect 2914 6279 2972 6291
rect 3072 7267 3130 7279
rect 3072 6291 3084 7267
rect 3118 6291 3130 7267
rect 3072 6279 3130 6291
rect 3230 7267 3288 7279
rect 3230 6291 3242 7267
rect 3276 6291 3288 7267
rect 3230 6279 3288 6291
rect 3388 7267 3446 7279
rect 3388 6291 3400 7267
rect 3434 6291 3446 7267
rect 3388 6279 3446 6291
rect 3546 7267 3604 7279
rect 3546 6291 3558 7267
rect 3592 6291 3604 7267
rect 3546 6279 3604 6291
<< ndiffc >>
rect 1341 4723 1375 5699
rect 1499 4723 1533 5699
rect 1657 4723 1691 5699
rect 1815 4723 1849 5699
rect 1973 4723 2007 5699
rect 2131 4723 2165 5699
rect 2289 4723 2323 5699
rect 2447 4723 2481 5699
rect 1341 3203 1375 4179
rect 1499 3203 1533 4179
rect 1657 3203 1691 4179
rect 1815 3203 1849 4179
rect 1973 3203 2007 4179
rect 2131 3203 2165 4179
rect 2289 3203 2323 4179
rect 2447 3203 2481 4179
rect 350 1682 384 2658
rect 608 1682 642 2658
rect 866 1682 900 2658
rect 1124 1682 1158 2658
rect 1382 1682 1416 2658
rect 1640 1682 1674 2658
rect 1898 1682 1932 2658
rect 2156 1682 2190 2658
rect 2414 1682 2448 2658
rect 2672 1682 2706 2658
rect 2930 1682 2964 2658
rect 3188 1682 3222 2658
rect 3446 1682 3480 2658
rect 90 162 124 1138
rect 348 162 382 1138
rect 606 162 640 1138
rect 864 162 898 1138
rect 1122 162 1156 1138
rect 1380 162 1414 1138
rect 1638 162 1672 1138
rect 1896 162 1930 1138
rect 2154 162 2188 1138
rect 2412 162 2446 1138
rect 2670 162 2704 1138
rect 2928 162 2962 1138
rect 3186 162 3220 1138
rect 3444 162 3478 1138
rect 3702 162 3736 1138
<< pdiffc >>
rect -1260 9501 -1226 10477
rect -1102 9501 -1068 10477
rect -944 9501 -910 10477
rect -786 9501 -752 10477
rect -628 9501 -594 10477
rect -470 9501 -436 10477
rect -312 9501 -278 10477
rect -154 9501 -120 10477
rect 4 9501 38 10477
rect 162 9501 196 10477
rect 320 9501 354 10477
rect 478 9501 512 10477
rect 636 9501 670 10477
rect 794 9501 828 10477
rect 952 9501 986 10477
rect 1110 9501 1144 10477
rect 1268 9501 1302 10477
rect 1426 9501 1460 10477
rect 1584 9501 1618 10477
rect 1742 9501 1776 10477
rect 1900 9501 1934 10477
rect 2058 9501 2092 10477
rect 2216 9501 2250 10477
rect 2374 9501 2408 10477
rect 2532 9501 2566 10477
rect 2690 9501 2724 10477
rect 2848 9501 2882 10477
rect 3006 9501 3040 10477
rect 3164 9501 3198 10477
rect 3322 9501 3356 10477
rect 3480 9501 3514 10477
rect 3638 9501 3672 10477
rect 3796 9501 3830 10477
rect 3954 9501 3988 10477
rect 4112 9501 4146 10477
rect 4270 9501 4304 10477
rect 4428 9501 4462 10477
rect 4586 9501 4620 10477
rect 4744 9501 4778 10477
rect 4902 9501 4936 10477
rect 5060 9501 5094 10477
rect 240 7831 274 8807
rect 398 7831 432 8807
rect 556 7831 590 8807
rect 714 7831 748 8807
rect 872 7831 906 8807
rect 1030 7831 1064 8807
rect 1188 7831 1222 8807
rect 1346 7831 1380 8807
rect 1504 7831 1538 8807
rect 1662 7831 1696 8807
rect 1820 7831 1854 8807
rect 1978 7831 2012 8807
rect 2136 7831 2170 8807
rect 2294 7831 2328 8807
rect 2452 7831 2486 8807
rect 2610 7831 2644 8807
rect 2768 7831 2802 8807
rect 2926 7831 2960 8807
rect 3084 7831 3118 8807
rect 3242 7831 3276 8807
rect 3400 7831 3434 8807
rect 3558 7831 3592 8807
rect 240 6291 274 7267
rect 398 6291 432 7267
rect 556 6291 590 7267
rect 714 6291 748 7267
rect 872 6291 906 7267
rect 1030 6291 1064 7267
rect 1188 6291 1222 7267
rect 1346 6291 1380 7267
rect 1504 6291 1538 7267
rect 1662 6291 1696 7267
rect 1820 6291 1854 7267
rect 1978 6291 2012 7267
rect 2136 6291 2170 7267
rect 2294 6291 2328 7267
rect 2452 6291 2486 7267
rect 2610 6291 2644 7267
rect 2768 6291 2802 7267
rect 2926 6291 2960 7267
rect 3084 6291 3118 7267
rect 3242 6291 3276 7267
rect 3400 6291 3434 7267
rect 3558 6291 3592 7267
<< psubdiff >>
rect -5177 11515 -5081 11549
rect -2149 11515 -2053 11549
rect -5177 11453 -5143 11515
rect -2087 11453 -2053 11515
rect -5177 10177 -5143 10239
rect 6553 11515 6649 11549
rect 9581 11515 9677 11549
rect 6553 11453 6587 11515
rect -2087 10177 -2053 10239
rect -5177 10143 -5081 10177
rect -2149 10143 -2053 10177
rect -5177 10055 -5081 10089
rect -2149 10055 -2053 10089
rect -5177 9993 -5143 10055
rect -2087 9993 -2053 10055
rect -5177 8717 -5143 8779
rect 9643 11453 9677 11515
rect 6553 10177 6587 10239
rect 9643 10177 9677 10239
rect 6553 10143 6649 10177
rect 9581 10143 9677 10177
rect 6553 10055 6649 10089
rect 9581 10055 9677 10089
rect 6553 9993 6587 10055
rect -2087 8717 -2053 8779
rect -5177 8683 -5081 8717
rect -2149 8683 -2053 8717
rect -4610 8220 -4480 8244
rect -4610 8036 -4480 8060
rect -2940 8230 -2810 8254
rect -2940 8046 -2810 8070
rect 9643 9993 9677 10055
rect 6553 8717 6587 8779
rect 9643 8717 9677 8779
rect 6553 8683 6649 8717
rect 9581 8683 9677 8717
rect 7010 8360 7120 8384
rect 7010 8206 7120 8230
rect 8890 8350 9000 8374
rect 8890 8196 9000 8220
rect 1227 5851 1323 5885
rect 2499 5851 2595 5885
rect 1227 5789 1261 5851
rect 2561 5789 2595 5851
rect 1227 4571 1261 4633
rect 2561 4571 2595 4633
rect 1227 4537 1323 4571
rect 2499 4537 2595 4571
rect 1227 4331 1323 4365
rect 2499 4331 2595 4365
rect 1227 4269 1261 4331
rect 2561 4269 2595 4331
rect 1227 3051 1261 3113
rect 2561 3051 2595 3113
rect 1227 3017 1323 3051
rect 2499 3017 2595 3051
rect 236 2810 332 2844
rect 3498 2810 3594 2844
rect 236 2748 270 2810
rect 3560 2748 3594 2810
rect 236 1530 270 1592
rect 3560 1530 3594 1592
rect 236 1496 332 1530
rect 3498 1496 3594 1530
rect -24 1290 72 1324
rect 3754 1290 3850 1324
rect -24 1228 10 1290
rect 3816 1228 3850 1290
rect -24 10 10 72
rect 3816 10 3850 72
rect -24 -24 72 10
rect 3754 -24 3850 10
<< nsubdiff >>
rect -1374 10638 -1278 10672
rect 5112 10638 5208 10672
rect -1374 10576 -1340 10638
rect 5174 10576 5208 10638
rect -1374 9340 -1340 9402
rect 5174 9340 5208 9402
rect -1374 9306 -1278 9340
rect 5112 9306 5208 9340
rect 126 8968 222 9002
rect 3610 8968 3706 9002
rect 126 8906 160 8968
rect 3672 8906 3706 8968
rect 126 7670 160 7732
rect 3672 7670 3706 7732
rect 126 7636 222 7670
rect 3610 7636 3706 7670
rect 126 7428 222 7462
rect 3610 7428 3706 7462
rect 126 7366 160 7428
rect 3672 7366 3706 7428
rect 126 6130 160 6192
rect 3672 6130 3706 6192
rect 126 6096 222 6130
rect 3610 6096 3706 6130
<< psubdiffcont >>
rect -5081 11515 -2149 11549
rect -5177 10239 -5143 11453
rect -2087 10239 -2053 11453
rect 6649 11515 9581 11549
rect -5081 10143 -2149 10177
rect -5081 10055 -2149 10089
rect -5177 8779 -5143 9993
rect -2087 8779 -2053 9993
rect 6553 10239 6587 11453
rect 9643 10239 9677 11453
rect 6649 10143 9581 10177
rect 6649 10055 9581 10089
rect -5081 8683 -2149 8717
rect -4610 8060 -4480 8220
rect -2940 8070 -2810 8230
rect 6553 8779 6587 9993
rect 9643 8779 9677 9993
rect 6649 8683 9581 8717
rect 7010 8230 7120 8360
rect 8890 8220 9000 8350
rect 1323 5851 2499 5885
rect 1227 4633 1261 5789
rect 2561 4633 2595 5789
rect 1323 4537 2499 4571
rect 1323 4331 2499 4365
rect 1227 3113 1261 4269
rect 2561 3113 2595 4269
rect 1323 3017 2499 3051
rect 332 2810 3498 2844
rect 236 1592 270 2748
rect 3560 1592 3594 2748
rect 332 1496 3498 1530
rect 72 1290 3754 1324
rect -24 72 10 1228
rect 3816 72 3850 1228
rect 72 -24 3754 10
<< nsubdiffcont >>
rect -1278 10638 5112 10672
rect -1374 9402 -1340 10576
rect 5174 9402 5208 10576
rect -1278 9306 5112 9340
rect 222 8968 3610 9002
rect 126 7732 160 8906
rect 3672 7732 3706 8906
rect 222 7636 3610 7670
rect 222 7428 3610 7462
rect 126 6192 160 7366
rect 3672 6192 3706 7366
rect 222 6096 3610 6130
<< poly >>
rect -1214 10570 -1114 10586
rect -1214 10536 -1198 10570
rect -1130 10536 -1114 10570
rect -1214 10489 -1114 10536
rect -1056 10570 -956 10586
rect -1056 10536 -1040 10570
rect -972 10536 -956 10570
rect -1056 10489 -956 10536
rect -898 10570 -798 10586
rect -898 10536 -882 10570
rect -814 10536 -798 10570
rect -898 10489 -798 10536
rect -740 10570 -640 10586
rect -740 10536 -724 10570
rect -656 10536 -640 10570
rect -740 10489 -640 10536
rect -582 10570 -482 10586
rect -582 10536 -566 10570
rect -498 10536 -482 10570
rect -582 10489 -482 10536
rect -424 10570 -324 10586
rect -424 10536 -408 10570
rect -340 10536 -324 10570
rect -424 10489 -324 10536
rect -266 10570 -166 10586
rect -266 10536 -250 10570
rect -182 10536 -166 10570
rect -266 10489 -166 10536
rect -108 10570 -8 10586
rect -108 10536 -92 10570
rect -24 10536 -8 10570
rect -108 10489 -8 10536
rect 50 10570 150 10586
rect 50 10536 66 10570
rect 134 10536 150 10570
rect 50 10489 150 10536
rect 208 10570 308 10586
rect 208 10536 224 10570
rect 292 10536 308 10570
rect 208 10489 308 10536
rect 366 10570 466 10586
rect 366 10536 382 10570
rect 450 10536 466 10570
rect 366 10489 466 10536
rect 524 10570 624 10586
rect 524 10536 540 10570
rect 608 10536 624 10570
rect 524 10489 624 10536
rect 682 10570 782 10586
rect 682 10536 698 10570
rect 766 10536 782 10570
rect 682 10489 782 10536
rect 840 10570 940 10586
rect 840 10536 856 10570
rect 924 10536 940 10570
rect 840 10489 940 10536
rect 998 10570 1098 10586
rect 998 10536 1014 10570
rect 1082 10536 1098 10570
rect 998 10489 1098 10536
rect 1156 10570 1256 10586
rect 1156 10536 1172 10570
rect 1240 10536 1256 10570
rect 1156 10489 1256 10536
rect 1314 10570 1414 10586
rect 1314 10536 1330 10570
rect 1398 10536 1414 10570
rect 1314 10489 1414 10536
rect 1472 10570 1572 10586
rect 1472 10536 1488 10570
rect 1556 10536 1572 10570
rect 1472 10489 1572 10536
rect 1630 10570 1730 10586
rect 1630 10536 1646 10570
rect 1714 10536 1730 10570
rect 1630 10489 1730 10536
rect 1788 10570 1888 10586
rect 1788 10536 1804 10570
rect 1872 10536 1888 10570
rect 1788 10489 1888 10536
rect 1946 10570 2046 10586
rect 1946 10536 1962 10570
rect 2030 10536 2046 10570
rect 1946 10489 2046 10536
rect 2104 10570 2204 10586
rect 2104 10536 2120 10570
rect 2188 10536 2204 10570
rect 2104 10489 2204 10536
rect 2262 10570 2362 10586
rect 2262 10536 2278 10570
rect 2346 10536 2362 10570
rect 2262 10489 2362 10536
rect 2420 10570 2520 10586
rect 2420 10536 2436 10570
rect 2504 10536 2520 10570
rect 2420 10489 2520 10536
rect 2578 10570 2678 10586
rect 2578 10536 2594 10570
rect 2662 10536 2678 10570
rect 2578 10489 2678 10536
rect 2736 10570 2836 10586
rect 2736 10536 2752 10570
rect 2820 10536 2836 10570
rect 2736 10489 2836 10536
rect 2894 10570 2994 10586
rect 2894 10536 2910 10570
rect 2978 10536 2994 10570
rect 2894 10489 2994 10536
rect 3052 10570 3152 10586
rect 3052 10536 3068 10570
rect 3136 10536 3152 10570
rect 3052 10489 3152 10536
rect 3210 10570 3310 10586
rect 3210 10536 3226 10570
rect 3294 10536 3310 10570
rect 3210 10489 3310 10536
rect 3368 10570 3468 10586
rect 3368 10536 3384 10570
rect 3452 10536 3468 10570
rect 3368 10489 3468 10536
rect 3526 10570 3626 10586
rect 3526 10536 3542 10570
rect 3610 10536 3626 10570
rect 3526 10489 3626 10536
rect 3684 10570 3784 10586
rect 3684 10536 3700 10570
rect 3768 10536 3784 10570
rect 3684 10489 3784 10536
rect 3842 10570 3942 10586
rect 3842 10536 3858 10570
rect 3926 10536 3942 10570
rect 3842 10489 3942 10536
rect 4000 10570 4100 10586
rect 4000 10536 4016 10570
rect 4084 10536 4100 10570
rect 4000 10489 4100 10536
rect 4158 10570 4258 10586
rect 4158 10536 4174 10570
rect 4242 10536 4258 10570
rect 4158 10489 4258 10536
rect 4316 10570 4416 10586
rect 4316 10536 4332 10570
rect 4400 10536 4416 10570
rect 4316 10489 4416 10536
rect 4474 10570 4574 10586
rect 4474 10536 4490 10570
rect 4558 10536 4574 10570
rect 4474 10489 4574 10536
rect 4632 10570 4732 10586
rect 4632 10536 4648 10570
rect 4716 10536 4732 10570
rect 4632 10489 4732 10536
rect 4790 10570 4890 10586
rect 4790 10536 4806 10570
rect 4874 10536 4890 10570
rect 4790 10489 4890 10536
rect 4948 10570 5048 10586
rect 4948 10536 4964 10570
rect 5032 10536 5048 10570
rect 4948 10489 5048 10536
rect -1214 9442 -1114 9489
rect -1214 9408 -1198 9442
rect -1130 9408 -1114 9442
rect -1214 9392 -1114 9408
rect -1056 9442 -956 9489
rect -1056 9408 -1040 9442
rect -972 9408 -956 9442
rect -1056 9392 -956 9408
rect -898 9442 -798 9489
rect -898 9408 -882 9442
rect -814 9408 -798 9442
rect -898 9392 -798 9408
rect -740 9442 -640 9489
rect -740 9408 -724 9442
rect -656 9408 -640 9442
rect -740 9392 -640 9408
rect -582 9442 -482 9489
rect -582 9408 -566 9442
rect -498 9408 -482 9442
rect -582 9392 -482 9408
rect -424 9442 -324 9489
rect -424 9408 -408 9442
rect -340 9408 -324 9442
rect -424 9392 -324 9408
rect -266 9442 -166 9489
rect -266 9408 -250 9442
rect -182 9408 -166 9442
rect -266 9392 -166 9408
rect -108 9442 -8 9489
rect -108 9408 -92 9442
rect -24 9408 -8 9442
rect -108 9392 -8 9408
rect 50 9442 150 9489
rect 50 9408 66 9442
rect 134 9408 150 9442
rect 50 9392 150 9408
rect 208 9442 308 9489
rect 208 9408 224 9442
rect 292 9408 308 9442
rect 208 9392 308 9408
rect 366 9442 466 9489
rect 366 9408 382 9442
rect 450 9408 466 9442
rect 366 9392 466 9408
rect 524 9442 624 9489
rect 524 9408 540 9442
rect 608 9408 624 9442
rect 524 9392 624 9408
rect 682 9442 782 9489
rect 682 9408 698 9442
rect 766 9408 782 9442
rect 682 9392 782 9408
rect 840 9442 940 9489
rect 840 9408 856 9442
rect 924 9408 940 9442
rect 840 9392 940 9408
rect 998 9442 1098 9489
rect 998 9408 1014 9442
rect 1082 9408 1098 9442
rect 998 9392 1098 9408
rect 1156 9442 1256 9489
rect 1156 9408 1172 9442
rect 1240 9408 1256 9442
rect 1156 9392 1256 9408
rect 1314 9442 1414 9489
rect 1314 9408 1330 9442
rect 1398 9408 1414 9442
rect 1314 9392 1414 9408
rect 1472 9442 1572 9489
rect 1472 9408 1488 9442
rect 1556 9408 1572 9442
rect 1472 9392 1572 9408
rect 1630 9442 1730 9489
rect 1630 9408 1646 9442
rect 1714 9408 1730 9442
rect 1630 9392 1730 9408
rect 1788 9442 1888 9489
rect 1788 9408 1804 9442
rect 1872 9408 1888 9442
rect 1788 9392 1888 9408
rect 1946 9442 2046 9489
rect 1946 9408 1962 9442
rect 2030 9408 2046 9442
rect 1946 9392 2046 9408
rect 2104 9442 2204 9489
rect 2104 9408 2120 9442
rect 2188 9408 2204 9442
rect 2104 9392 2204 9408
rect 2262 9442 2362 9489
rect 2262 9408 2278 9442
rect 2346 9408 2362 9442
rect 2262 9392 2362 9408
rect 2420 9442 2520 9489
rect 2420 9408 2436 9442
rect 2504 9408 2520 9442
rect 2420 9392 2520 9408
rect 2578 9442 2678 9489
rect 2578 9408 2594 9442
rect 2662 9408 2678 9442
rect 2578 9392 2678 9408
rect 2736 9442 2836 9489
rect 2736 9408 2752 9442
rect 2820 9408 2836 9442
rect 2736 9392 2836 9408
rect 2894 9442 2994 9489
rect 2894 9408 2910 9442
rect 2978 9408 2994 9442
rect 2894 9392 2994 9408
rect 3052 9442 3152 9489
rect 3052 9408 3068 9442
rect 3136 9408 3152 9442
rect 3052 9392 3152 9408
rect 3210 9442 3310 9489
rect 3210 9408 3226 9442
rect 3294 9408 3310 9442
rect 3210 9392 3310 9408
rect 3368 9442 3468 9489
rect 3368 9408 3384 9442
rect 3452 9408 3468 9442
rect 3368 9392 3468 9408
rect 3526 9442 3626 9489
rect 3526 9408 3542 9442
rect 3610 9408 3626 9442
rect 3526 9392 3626 9408
rect 3684 9442 3784 9489
rect 3684 9408 3700 9442
rect 3768 9408 3784 9442
rect 3684 9392 3784 9408
rect 3842 9442 3942 9489
rect 3842 9408 3858 9442
rect 3926 9408 3942 9442
rect 3842 9392 3942 9408
rect 4000 9442 4100 9489
rect 4000 9408 4016 9442
rect 4084 9408 4100 9442
rect 4000 9392 4100 9408
rect 4158 9442 4258 9489
rect 4158 9408 4174 9442
rect 4242 9408 4258 9442
rect 4158 9392 4258 9408
rect 4316 9442 4416 9489
rect 4316 9408 4332 9442
rect 4400 9408 4416 9442
rect 4316 9392 4416 9408
rect 4474 9442 4574 9489
rect 4474 9408 4490 9442
rect 4558 9408 4574 9442
rect 4474 9392 4574 9408
rect 4632 9442 4732 9489
rect 4632 9408 4648 9442
rect 4716 9408 4732 9442
rect 4632 9392 4732 9408
rect 4790 9442 4890 9489
rect 4790 9408 4806 9442
rect 4874 9408 4890 9442
rect 4790 9392 4890 9408
rect 4948 9442 5048 9489
rect 4948 9408 4964 9442
rect 5032 9408 5048 9442
rect 4948 9392 5048 9408
rect 286 8900 386 8916
rect 286 8866 302 8900
rect 370 8866 386 8900
rect 286 8819 386 8866
rect 444 8900 544 8916
rect 444 8866 460 8900
rect 528 8866 544 8900
rect 444 8819 544 8866
rect 602 8900 702 8916
rect 602 8866 618 8900
rect 686 8866 702 8900
rect 602 8819 702 8866
rect 760 8900 860 8916
rect 760 8866 776 8900
rect 844 8866 860 8900
rect 760 8819 860 8866
rect 918 8900 1018 8916
rect 918 8866 934 8900
rect 1002 8866 1018 8900
rect 918 8819 1018 8866
rect 1076 8900 1176 8916
rect 1076 8866 1092 8900
rect 1160 8866 1176 8900
rect 1076 8819 1176 8866
rect 1234 8900 1334 8916
rect 1234 8866 1250 8900
rect 1318 8866 1334 8900
rect 1234 8819 1334 8866
rect 1392 8900 1492 8916
rect 1392 8866 1408 8900
rect 1476 8866 1492 8900
rect 1392 8819 1492 8866
rect 1550 8900 1650 8916
rect 1550 8866 1566 8900
rect 1634 8866 1650 8900
rect 1550 8819 1650 8866
rect 1708 8900 1808 8916
rect 1708 8866 1724 8900
rect 1792 8866 1808 8900
rect 1708 8819 1808 8866
rect 1866 8900 1966 8916
rect 1866 8866 1882 8900
rect 1950 8866 1966 8900
rect 1866 8819 1966 8866
rect 2024 8900 2124 8916
rect 2024 8866 2040 8900
rect 2108 8866 2124 8900
rect 2024 8819 2124 8866
rect 2182 8900 2282 8916
rect 2182 8866 2198 8900
rect 2266 8866 2282 8900
rect 2182 8819 2282 8866
rect 2340 8900 2440 8916
rect 2340 8866 2356 8900
rect 2424 8866 2440 8900
rect 2340 8819 2440 8866
rect 2498 8900 2598 8916
rect 2498 8866 2514 8900
rect 2582 8866 2598 8900
rect 2498 8819 2598 8866
rect 2656 8900 2756 8916
rect 2656 8866 2672 8900
rect 2740 8866 2756 8900
rect 2656 8819 2756 8866
rect 2814 8900 2914 8916
rect 2814 8866 2830 8900
rect 2898 8866 2914 8900
rect 2814 8819 2914 8866
rect 2972 8900 3072 8916
rect 2972 8866 2988 8900
rect 3056 8866 3072 8900
rect 2972 8819 3072 8866
rect 3130 8900 3230 8916
rect 3130 8866 3146 8900
rect 3214 8866 3230 8900
rect 3130 8819 3230 8866
rect 3288 8900 3388 8916
rect 3288 8866 3304 8900
rect 3372 8866 3388 8900
rect 3288 8819 3388 8866
rect 3446 8900 3546 8916
rect 3446 8866 3462 8900
rect 3530 8866 3546 8900
rect 3446 8819 3546 8866
rect 286 7772 386 7819
rect 286 7738 302 7772
rect 370 7738 386 7772
rect 286 7722 386 7738
rect 444 7772 544 7819
rect 444 7738 460 7772
rect 528 7738 544 7772
rect 444 7722 544 7738
rect 602 7772 702 7819
rect 602 7738 618 7772
rect 686 7738 702 7772
rect 602 7722 702 7738
rect 760 7772 860 7819
rect 760 7738 776 7772
rect 844 7738 860 7772
rect 760 7722 860 7738
rect 918 7772 1018 7819
rect 918 7738 934 7772
rect 1002 7738 1018 7772
rect 918 7722 1018 7738
rect 1076 7772 1176 7819
rect 1076 7738 1092 7772
rect 1160 7738 1176 7772
rect 1076 7722 1176 7738
rect 1234 7772 1334 7819
rect 1234 7738 1250 7772
rect 1318 7738 1334 7772
rect 1234 7722 1334 7738
rect 1392 7772 1492 7819
rect 1392 7738 1408 7772
rect 1476 7738 1492 7772
rect 1392 7722 1492 7738
rect 1550 7772 1650 7819
rect 1550 7738 1566 7772
rect 1634 7738 1650 7772
rect 1550 7722 1650 7738
rect 1708 7772 1808 7819
rect 1708 7738 1724 7772
rect 1792 7738 1808 7772
rect 1708 7722 1808 7738
rect 1866 7772 1966 7819
rect 1866 7738 1882 7772
rect 1950 7738 1966 7772
rect 1866 7722 1966 7738
rect 2024 7772 2124 7819
rect 2024 7738 2040 7772
rect 2108 7738 2124 7772
rect 2024 7722 2124 7738
rect 2182 7772 2282 7819
rect 2182 7738 2198 7772
rect 2266 7738 2282 7772
rect 2182 7722 2282 7738
rect 2340 7772 2440 7819
rect 2340 7738 2356 7772
rect 2424 7738 2440 7772
rect 2340 7722 2440 7738
rect 2498 7772 2598 7819
rect 2498 7738 2514 7772
rect 2582 7738 2598 7772
rect 2498 7722 2598 7738
rect 2656 7772 2756 7819
rect 2656 7738 2672 7772
rect 2740 7738 2756 7772
rect 2656 7722 2756 7738
rect 2814 7772 2914 7819
rect 2814 7738 2830 7772
rect 2898 7738 2914 7772
rect 2814 7722 2914 7738
rect 2972 7772 3072 7819
rect 2972 7738 2988 7772
rect 3056 7738 3072 7772
rect 2972 7722 3072 7738
rect 3130 7772 3230 7819
rect 3130 7738 3146 7772
rect 3214 7738 3230 7772
rect 3130 7722 3230 7738
rect 3288 7772 3388 7819
rect 3288 7738 3304 7772
rect 3372 7738 3388 7772
rect 3288 7722 3388 7738
rect 3446 7772 3546 7819
rect 3446 7738 3462 7772
rect 3530 7738 3546 7772
rect 3446 7722 3546 7738
rect 286 7360 386 7376
rect 286 7326 302 7360
rect 370 7326 386 7360
rect 286 7279 386 7326
rect 444 7360 544 7376
rect 444 7326 460 7360
rect 528 7326 544 7360
rect 444 7279 544 7326
rect 602 7360 702 7376
rect 602 7326 618 7360
rect 686 7326 702 7360
rect 602 7279 702 7326
rect 760 7360 860 7376
rect 760 7326 776 7360
rect 844 7326 860 7360
rect 760 7279 860 7326
rect 918 7360 1018 7376
rect 918 7326 934 7360
rect 1002 7326 1018 7360
rect 918 7279 1018 7326
rect 1076 7360 1176 7376
rect 1076 7326 1092 7360
rect 1160 7326 1176 7360
rect 1076 7279 1176 7326
rect 1234 7360 1334 7376
rect 1234 7326 1250 7360
rect 1318 7326 1334 7360
rect 1234 7279 1334 7326
rect 1392 7360 1492 7376
rect 1392 7326 1408 7360
rect 1476 7326 1492 7360
rect 1392 7279 1492 7326
rect 1550 7360 1650 7376
rect 1550 7326 1566 7360
rect 1634 7326 1650 7360
rect 1550 7279 1650 7326
rect 1708 7360 1808 7376
rect 1708 7326 1724 7360
rect 1792 7326 1808 7360
rect 1708 7279 1808 7326
rect 1866 7360 1966 7376
rect 1866 7326 1882 7360
rect 1950 7326 1966 7360
rect 1866 7279 1966 7326
rect 2024 7360 2124 7376
rect 2024 7326 2040 7360
rect 2108 7326 2124 7360
rect 2024 7279 2124 7326
rect 2182 7360 2282 7376
rect 2182 7326 2198 7360
rect 2266 7326 2282 7360
rect 2182 7279 2282 7326
rect 2340 7360 2440 7376
rect 2340 7326 2356 7360
rect 2424 7326 2440 7360
rect 2340 7279 2440 7326
rect 2498 7360 2598 7376
rect 2498 7326 2514 7360
rect 2582 7326 2598 7360
rect 2498 7279 2598 7326
rect 2656 7360 2756 7376
rect 2656 7326 2672 7360
rect 2740 7326 2756 7360
rect 2656 7279 2756 7326
rect 2814 7360 2914 7376
rect 2814 7326 2830 7360
rect 2898 7326 2914 7360
rect 2814 7279 2914 7326
rect 2972 7360 3072 7376
rect 2972 7326 2988 7360
rect 3056 7326 3072 7360
rect 2972 7279 3072 7326
rect 3130 7360 3230 7376
rect 3130 7326 3146 7360
rect 3214 7326 3230 7360
rect 3130 7279 3230 7326
rect 3288 7360 3388 7376
rect 3288 7326 3304 7360
rect 3372 7326 3388 7360
rect 3288 7279 3388 7326
rect 3446 7360 3546 7376
rect 3446 7326 3462 7360
rect 3530 7326 3546 7360
rect 3446 7279 3546 7326
rect 286 6232 386 6279
rect 286 6198 302 6232
rect 370 6198 386 6232
rect 286 6182 386 6198
rect 444 6232 544 6279
rect 444 6198 460 6232
rect 528 6198 544 6232
rect 444 6182 544 6198
rect 602 6232 702 6279
rect 602 6198 618 6232
rect 686 6198 702 6232
rect 602 6182 702 6198
rect 760 6232 860 6279
rect 760 6198 776 6232
rect 844 6198 860 6232
rect 760 6182 860 6198
rect 918 6232 1018 6279
rect 918 6198 934 6232
rect 1002 6198 1018 6232
rect 918 6182 1018 6198
rect 1076 6232 1176 6279
rect 1076 6198 1092 6232
rect 1160 6198 1176 6232
rect 1076 6182 1176 6198
rect 1234 6232 1334 6279
rect 1234 6198 1250 6232
rect 1318 6198 1334 6232
rect 1234 6182 1334 6198
rect 1392 6232 1492 6279
rect 1392 6198 1408 6232
rect 1476 6198 1492 6232
rect 1392 6182 1492 6198
rect 1550 6232 1650 6279
rect 1550 6198 1566 6232
rect 1634 6198 1650 6232
rect 1550 6182 1650 6198
rect 1708 6232 1808 6279
rect 1708 6198 1724 6232
rect 1792 6198 1808 6232
rect 1708 6182 1808 6198
rect 1866 6232 1966 6279
rect 1866 6198 1882 6232
rect 1950 6198 1966 6232
rect 1866 6182 1966 6198
rect 2024 6232 2124 6279
rect 2024 6198 2040 6232
rect 2108 6198 2124 6232
rect 2024 6182 2124 6198
rect 2182 6232 2282 6279
rect 2182 6198 2198 6232
rect 2266 6198 2282 6232
rect 2182 6182 2282 6198
rect 2340 6232 2440 6279
rect 2340 6198 2356 6232
rect 2424 6198 2440 6232
rect 2340 6182 2440 6198
rect 2498 6232 2598 6279
rect 2498 6198 2514 6232
rect 2582 6198 2598 6232
rect 2498 6182 2598 6198
rect 2656 6232 2756 6279
rect 2656 6198 2672 6232
rect 2740 6198 2756 6232
rect 2656 6182 2756 6198
rect 2814 6232 2914 6279
rect 2814 6198 2830 6232
rect 2898 6198 2914 6232
rect 2814 6182 2914 6198
rect 2972 6232 3072 6279
rect 2972 6198 2988 6232
rect 3056 6198 3072 6232
rect 2972 6182 3072 6198
rect 3130 6232 3230 6279
rect 3130 6198 3146 6232
rect 3214 6198 3230 6232
rect 3130 6182 3230 6198
rect 3288 6232 3388 6279
rect 3288 6198 3304 6232
rect 3372 6198 3388 6232
rect 3288 6182 3388 6198
rect 3446 6232 3546 6279
rect 3446 6198 3462 6232
rect 3530 6198 3546 6232
rect 3446 6182 3546 6198
rect 1387 5783 1487 5799
rect 1387 5749 1403 5783
rect 1471 5749 1487 5783
rect 1387 5711 1487 5749
rect 1545 5783 1645 5799
rect 1545 5749 1561 5783
rect 1629 5749 1645 5783
rect 1545 5711 1645 5749
rect 1703 5783 1803 5799
rect 1703 5749 1719 5783
rect 1787 5749 1803 5783
rect 1703 5711 1803 5749
rect 1861 5783 1961 5799
rect 1861 5749 1877 5783
rect 1945 5749 1961 5783
rect 1861 5711 1961 5749
rect 2019 5783 2119 5799
rect 2019 5749 2035 5783
rect 2103 5749 2119 5783
rect 2019 5711 2119 5749
rect 2177 5783 2277 5799
rect 2177 5749 2193 5783
rect 2261 5749 2277 5783
rect 2177 5711 2277 5749
rect 2335 5783 2435 5799
rect 2335 5749 2351 5783
rect 2419 5749 2435 5783
rect 2335 5711 2435 5749
rect 1387 4673 1487 4711
rect 1387 4639 1403 4673
rect 1471 4639 1487 4673
rect 1387 4623 1487 4639
rect 1545 4673 1645 4711
rect 1545 4639 1561 4673
rect 1629 4639 1645 4673
rect 1545 4623 1645 4639
rect 1703 4673 1803 4711
rect 1703 4639 1719 4673
rect 1787 4639 1803 4673
rect 1703 4623 1803 4639
rect 1861 4673 1961 4711
rect 1861 4639 1877 4673
rect 1945 4639 1961 4673
rect 1861 4623 1961 4639
rect 2019 4673 2119 4711
rect 2019 4639 2035 4673
rect 2103 4639 2119 4673
rect 2019 4623 2119 4639
rect 2177 4673 2277 4711
rect 2177 4639 2193 4673
rect 2261 4639 2277 4673
rect 2177 4623 2277 4639
rect 2335 4673 2435 4711
rect 2335 4639 2351 4673
rect 2419 4639 2435 4673
rect 2335 4623 2435 4639
rect 1387 4263 1487 4279
rect 1387 4229 1403 4263
rect 1471 4229 1487 4263
rect 1387 4191 1487 4229
rect 1545 4263 1645 4279
rect 1545 4229 1561 4263
rect 1629 4229 1645 4263
rect 1545 4191 1645 4229
rect 1703 4263 1803 4279
rect 1703 4229 1719 4263
rect 1787 4229 1803 4263
rect 1703 4191 1803 4229
rect 1861 4263 1961 4279
rect 1861 4229 1877 4263
rect 1945 4229 1961 4263
rect 1861 4191 1961 4229
rect 2019 4263 2119 4279
rect 2019 4229 2035 4263
rect 2103 4229 2119 4263
rect 2019 4191 2119 4229
rect 2177 4263 2277 4279
rect 2177 4229 2193 4263
rect 2261 4229 2277 4263
rect 2177 4191 2277 4229
rect 2335 4263 2435 4279
rect 2335 4229 2351 4263
rect 2419 4229 2435 4263
rect 2335 4191 2435 4229
rect 1387 3153 1487 3191
rect 1387 3119 1403 3153
rect 1471 3119 1487 3153
rect 1387 3103 1487 3119
rect 1545 3153 1645 3191
rect 1545 3119 1561 3153
rect 1629 3119 1645 3153
rect 1545 3103 1645 3119
rect 1703 3153 1803 3191
rect 1703 3119 1719 3153
rect 1787 3119 1803 3153
rect 1703 3103 1803 3119
rect 1861 3153 1961 3191
rect 1861 3119 1877 3153
rect 1945 3119 1961 3153
rect 1861 3103 1961 3119
rect 2019 3153 2119 3191
rect 2019 3119 2035 3153
rect 2103 3119 2119 3153
rect 2019 3103 2119 3119
rect 2177 3153 2277 3191
rect 2177 3119 2193 3153
rect 2261 3119 2277 3153
rect 2177 3103 2277 3119
rect 2335 3153 2435 3191
rect 2335 3119 2351 3153
rect 2419 3119 2435 3153
rect 2335 3103 2435 3119
rect 396 2742 596 2758
rect 396 2708 412 2742
rect 580 2708 596 2742
rect 396 2670 596 2708
rect 654 2742 854 2758
rect 654 2708 670 2742
rect 838 2708 854 2742
rect 654 2670 854 2708
rect 912 2742 1112 2758
rect 912 2708 928 2742
rect 1096 2708 1112 2742
rect 912 2670 1112 2708
rect 1170 2742 1370 2758
rect 1170 2708 1186 2742
rect 1354 2708 1370 2742
rect 1170 2670 1370 2708
rect 1428 2742 1628 2758
rect 1428 2708 1444 2742
rect 1612 2708 1628 2742
rect 1428 2670 1628 2708
rect 1686 2742 1886 2758
rect 1686 2708 1702 2742
rect 1870 2708 1886 2742
rect 1686 2670 1886 2708
rect 1944 2742 2144 2758
rect 1944 2708 1960 2742
rect 2128 2708 2144 2742
rect 1944 2670 2144 2708
rect 2202 2742 2402 2758
rect 2202 2708 2218 2742
rect 2386 2708 2402 2742
rect 2202 2670 2402 2708
rect 2460 2742 2660 2758
rect 2460 2708 2476 2742
rect 2644 2708 2660 2742
rect 2460 2670 2660 2708
rect 2718 2742 2918 2758
rect 2718 2708 2734 2742
rect 2902 2708 2918 2742
rect 2718 2670 2918 2708
rect 2976 2742 3176 2758
rect 2976 2708 2992 2742
rect 3160 2708 3176 2742
rect 2976 2670 3176 2708
rect 3234 2742 3434 2758
rect 3234 2708 3250 2742
rect 3418 2708 3434 2742
rect 3234 2670 3434 2708
rect 396 1632 596 1670
rect 396 1598 412 1632
rect 580 1598 596 1632
rect 396 1582 596 1598
rect 654 1632 854 1670
rect 654 1598 670 1632
rect 838 1598 854 1632
rect 654 1582 854 1598
rect 912 1632 1112 1670
rect 912 1598 928 1632
rect 1096 1598 1112 1632
rect 912 1582 1112 1598
rect 1170 1632 1370 1670
rect 1170 1598 1186 1632
rect 1354 1598 1370 1632
rect 1170 1582 1370 1598
rect 1428 1632 1628 1670
rect 1428 1598 1444 1632
rect 1612 1598 1628 1632
rect 1428 1582 1628 1598
rect 1686 1632 1886 1670
rect 1686 1598 1702 1632
rect 1870 1598 1886 1632
rect 1686 1582 1886 1598
rect 1944 1632 2144 1670
rect 1944 1598 1960 1632
rect 2128 1598 2144 1632
rect 1944 1582 2144 1598
rect 2202 1632 2402 1670
rect 2202 1598 2218 1632
rect 2386 1598 2402 1632
rect 2202 1582 2402 1598
rect 2460 1632 2660 1670
rect 2460 1598 2476 1632
rect 2644 1598 2660 1632
rect 2460 1582 2660 1598
rect 2718 1632 2918 1670
rect 2718 1598 2734 1632
rect 2902 1598 2918 1632
rect 2718 1582 2918 1598
rect 2976 1632 3176 1670
rect 2976 1598 2992 1632
rect 3160 1598 3176 1632
rect 2976 1582 3176 1598
rect 3234 1632 3434 1670
rect 3234 1598 3250 1632
rect 3418 1598 3434 1632
rect 3234 1582 3434 1598
rect 136 1222 336 1238
rect 136 1188 152 1222
rect 320 1188 336 1222
rect 136 1150 336 1188
rect 394 1222 594 1238
rect 394 1188 410 1222
rect 578 1188 594 1222
rect 394 1150 594 1188
rect 652 1222 852 1238
rect 652 1188 668 1222
rect 836 1188 852 1222
rect 652 1150 852 1188
rect 910 1222 1110 1238
rect 910 1188 926 1222
rect 1094 1188 1110 1222
rect 910 1150 1110 1188
rect 1168 1222 1368 1238
rect 1168 1188 1184 1222
rect 1352 1188 1368 1222
rect 1168 1150 1368 1188
rect 1426 1222 1626 1238
rect 1426 1188 1442 1222
rect 1610 1188 1626 1222
rect 1426 1150 1626 1188
rect 1684 1222 1884 1238
rect 1684 1188 1700 1222
rect 1868 1188 1884 1222
rect 1684 1150 1884 1188
rect 1942 1222 2142 1238
rect 1942 1188 1958 1222
rect 2126 1188 2142 1222
rect 1942 1150 2142 1188
rect 2200 1222 2400 1238
rect 2200 1188 2216 1222
rect 2384 1188 2400 1222
rect 2200 1150 2400 1188
rect 2458 1222 2658 1238
rect 2458 1188 2474 1222
rect 2642 1188 2658 1222
rect 2458 1150 2658 1188
rect 2716 1222 2916 1238
rect 2716 1188 2732 1222
rect 2900 1188 2916 1222
rect 2716 1150 2916 1188
rect 2974 1222 3174 1238
rect 2974 1188 2990 1222
rect 3158 1188 3174 1222
rect 2974 1150 3174 1188
rect 3232 1222 3432 1238
rect 3232 1188 3248 1222
rect 3416 1188 3432 1222
rect 3232 1150 3432 1188
rect 3490 1222 3690 1238
rect 3490 1188 3506 1222
rect 3674 1188 3690 1222
rect 3490 1150 3690 1188
rect 136 112 336 150
rect 136 78 152 112
rect 320 78 336 112
rect 136 62 336 78
rect 394 112 594 150
rect 394 78 410 112
rect 578 78 594 112
rect 394 62 594 78
rect 652 112 852 150
rect 652 78 668 112
rect 836 78 852 112
rect 652 62 852 78
rect 910 112 1110 150
rect 910 78 926 112
rect 1094 78 1110 112
rect 910 62 1110 78
rect 1168 112 1368 150
rect 1168 78 1184 112
rect 1352 78 1368 112
rect 1168 62 1368 78
rect 1426 112 1626 150
rect 1426 78 1442 112
rect 1610 78 1626 112
rect 1426 62 1626 78
rect 1684 112 1884 150
rect 1684 78 1700 112
rect 1868 78 1884 112
rect 1684 62 1884 78
rect 1942 112 2142 150
rect 1942 78 1958 112
rect 2126 78 2142 112
rect 1942 62 2142 78
rect 2200 112 2400 150
rect 2200 78 2216 112
rect 2384 78 2400 112
rect 2200 62 2400 78
rect 2458 112 2658 150
rect 2458 78 2474 112
rect 2642 78 2658 112
rect 2458 62 2658 78
rect 2716 112 2916 150
rect 2716 78 2732 112
rect 2900 78 2916 112
rect 2716 62 2916 78
rect 2974 112 3174 150
rect 2974 78 2990 112
rect 3158 78 3174 112
rect 2974 62 3174 78
rect 3232 112 3432 150
rect 3232 78 3248 112
rect 3416 78 3432 112
rect 3232 62 3432 78
rect 3490 112 3690 150
rect 3490 78 3506 112
rect 3674 78 3690 112
rect 3490 62 3690 78
<< polycont >>
rect -1198 10536 -1130 10570
rect -1040 10536 -972 10570
rect -882 10536 -814 10570
rect -724 10536 -656 10570
rect -566 10536 -498 10570
rect -408 10536 -340 10570
rect -250 10536 -182 10570
rect -92 10536 -24 10570
rect 66 10536 134 10570
rect 224 10536 292 10570
rect 382 10536 450 10570
rect 540 10536 608 10570
rect 698 10536 766 10570
rect 856 10536 924 10570
rect 1014 10536 1082 10570
rect 1172 10536 1240 10570
rect 1330 10536 1398 10570
rect 1488 10536 1556 10570
rect 1646 10536 1714 10570
rect 1804 10536 1872 10570
rect 1962 10536 2030 10570
rect 2120 10536 2188 10570
rect 2278 10536 2346 10570
rect 2436 10536 2504 10570
rect 2594 10536 2662 10570
rect 2752 10536 2820 10570
rect 2910 10536 2978 10570
rect 3068 10536 3136 10570
rect 3226 10536 3294 10570
rect 3384 10536 3452 10570
rect 3542 10536 3610 10570
rect 3700 10536 3768 10570
rect 3858 10536 3926 10570
rect 4016 10536 4084 10570
rect 4174 10536 4242 10570
rect 4332 10536 4400 10570
rect 4490 10536 4558 10570
rect 4648 10536 4716 10570
rect 4806 10536 4874 10570
rect 4964 10536 5032 10570
rect -1198 9408 -1130 9442
rect -1040 9408 -972 9442
rect -882 9408 -814 9442
rect -724 9408 -656 9442
rect -566 9408 -498 9442
rect -408 9408 -340 9442
rect -250 9408 -182 9442
rect -92 9408 -24 9442
rect 66 9408 134 9442
rect 224 9408 292 9442
rect 382 9408 450 9442
rect 540 9408 608 9442
rect 698 9408 766 9442
rect 856 9408 924 9442
rect 1014 9408 1082 9442
rect 1172 9408 1240 9442
rect 1330 9408 1398 9442
rect 1488 9408 1556 9442
rect 1646 9408 1714 9442
rect 1804 9408 1872 9442
rect 1962 9408 2030 9442
rect 2120 9408 2188 9442
rect 2278 9408 2346 9442
rect 2436 9408 2504 9442
rect 2594 9408 2662 9442
rect 2752 9408 2820 9442
rect 2910 9408 2978 9442
rect 3068 9408 3136 9442
rect 3226 9408 3294 9442
rect 3384 9408 3452 9442
rect 3542 9408 3610 9442
rect 3700 9408 3768 9442
rect 3858 9408 3926 9442
rect 4016 9408 4084 9442
rect 4174 9408 4242 9442
rect 4332 9408 4400 9442
rect 4490 9408 4558 9442
rect 4648 9408 4716 9442
rect 4806 9408 4874 9442
rect 4964 9408 5032 9442
rect 302 8866 370 8900
rect 460 8866 528 8900
rect 618 8866 686 8900
rect 776 8866 844 8900
rect 934 8866 1002 8900
rect 1092 8866 1160 8900
rect 1250 8866 1318 8900
rect 1408 8866 1476 8900
rect 1566 8866 1634 8900
rect 1724 8866 1792 8900
rect 1882 8866 1950 8900
rect 2040 8866 2108 8900
rect 2198 8866 2266 8900
rect 2356 8866 2424 8900
rect 2514 8866 2582 8900
rect 2672 8866 2740 8900
rect 2830 8866 2898 8900
rect 2988 8866 3056 8900
rect 3146 8866 3214 8900
rect 3304 8866 3372 8900
rect 3462 8866 3530 8900
rect 302 7738 370 7772
rect 460 7738 528 7772
rect 618 7738 686 7772
rect 776 7738 844 7772
rect 934 7738 1002 7772
rect 1092 7738 1160 7772
rect 1250 7738 1318 7772
rect 1408 7738 1476 7772
rect 1566 7738 1634 7772
rect 1724 7738 1792 7772
rect 1882 7738 1950 7772
rect 2040 7738 2108 7772
rect 2198 7738 2266 7772
rect 2356 7738 2424 7772
rect 2514 7738 2582 7772
rect 2672 7738 2740 7772
rect 2830 7738 2898 7772
rect 2988 7738 3056 7772
rect 3146 7738 3214 7772
rect 3304 7738 3372 7772
rect 3462 7738 3530 7772
rect 302 7326 370 7360
rect 460 7326 528 7360
rect 618 7326 686 7360
rect 776 7326 844 7360
rect 934 7326 1002 7360
rect 1092 7326 1160 7360
rect 1250 7326 1318 7360
rect 1408 7326 1476 7360
rect 1566 7326 1634 7360
rect 1724 7326 1792 7360
rect 1882 7326 1950 7360
rect 2040 7326 2108 7360
rect 2198 7326 2266 7360
rect 2356 7326 2424 7360
rect 2514 7326 2582 7360
rect 2672 7326 2740 7360
rect 2830 7326 2898 7360
rect 2988 7326 3056 7360
rect 3146 7326 3214 7360
rect 3304 7326 3372 7360
rect 3462 7326 3530 7360
rect 302 6198 370 6232
rect 460 6198 528 6232
rect 618 6198 686 6232
rect 776 6198 844 6232
rect 934 6198 1002 6232
rect 1092 6198 1160 6232
rect 1250 6198 1318 6232
rect 1408 6198 1476 6232
rect 1566 6198 1634 6232
rect 1724 6198 1792 6232
rect 1882 6198 1950 6232
rect 2040 6198 2108 6232
rect 2198 6198 2266 6232
rect 2356 6198 2424 6232
rect 2514 6198 2582 6232
rect 2672 6198 2740 6232
rect 2830 6198 2898 6232
rect 2988 6198 3056 6232
rect 3146 6198 3214 6232
rect 3304 6198 3372 6232
rect 3462 6198 3530 6232
rect 1403 5749 1471 5783
rect 1561 5749 1629 5783
rect 1719 5749 1787 5783
rect 1877 5749 1945 5783
rect 2035 5749 2103 5783
rect 2193 5749 2261 5783
rect 2351 5749 2419 5783
rect 1403 4639 1471 4673
rect 1561 4639 1629 4673
rect 1719 4639 1787 4673
rect 1877 4639 1945 4673
rect 2035 4639 2103 4673
rect 2193 4639 2261 4673
rect 2351 4639 2419 4673
rect 1403 4229 1471 4263
rect 1561 4229 1629 4263
rect 1719 4229 1787 4263
rect 1877 4229 1945 4263
rect 2035 4229 2103 4263
rect 2193 4229 2261 4263
rect 2351 4229 2419 4263
rect 1403 3119 1471 3153
rect 1561 3119 1629 3153
rect 1719 3119 1787 3153
rect 1877 3119 1945 3153
rect 2035 3119 2103 3153
rect 2193 3119 2261 3153
rect 2351 3119 2419 3153
rect 412 2708 580 2742
rect 670 2708 838 2742
rect 928 2708 1096 2742
rect 1186 2708 1354 2742
rect 1444 2708 1612 2742
rect 1702 2708 1870 2742
rect 1960 2708 2128 2742
rect 2218 2708 2386 2742
rect 2476 2708 2644 2742
rect 2734 2708 2902 2742
rect 2992 2708 3160 2742
rect 3250 2708 3418 2742
rect 412 1598 580 1632
rect 670 1598 838 1632
rect 928 1598 1096 1632
rect 1186 1598 1354 1632
rect 1444 1598 1612 1632
rect 1702 1598 1870 1632
rect 1960 1598 2128 1632
rect 2218 1598 2386 1632
rect 2476 1598 2644 1632
rect 2734 1598 2902 1632
rect 2992 1598 3160 1632
rect 3250 1598 3418 1632
rect 152 1188 320 1222
rect 410 1188 578 1222
rect 668 1188 836 1222
rect 926 1188 1094 1222
rect 1184 1188 1352 1222
rect 1442 1188 1610 1222
rect 1700 1188 1868 1222
rect 1958 1188 2126 1222
rect 2216 1188 2384 1222
rect 2474 1188 2642 1222
rect 2732 1188 2900 1222
rect 2990 1188 3158 1222
rect 3248 1188 3416 1222
rect 3506 1188 3674 1222
rect 152 78 320 112
rect 410 78 578 112
rect 668 78 836 112
rect 926 78 1094 112
rect 1184 78 1352 112
rect 1442 78 1610 112
rect 1700 78 1868 112
rect 1958 78 2126 112
rect 2216 78 2384 112
rect 2474 78 2642 112
rect 2732 78 2900 112
rect 2990 78 3158 112
rect 3248 78 3416 112
rect 3506 78 3674 112
<< xpolycontact >>
rect -5047 10273 -4615 11419
rect -2615 10273 -2183 11419
rect -5047 8813 -4615 9959
rect -2615 8813 -2183 9959
rect 6683 10273 7115 11419
rect 9115 10273 9547 11419
rect 6683 8813 7115 9959
rect 9115 8813 9547 9959
<< xpolyres >>
rect -4615 10273 -2615 11419
rect -4615 8813 -2615 9959
rect 7115 10273 9115 11419
rect 7115 8813 9115 9959
<< locali >>
rect -5177 11515 -5081 11549
rect -2149 11515 -2053 11549
rect -5177 11453 -5143 11515
rect -2087 11453 -2053 11515
rect -5177 10177 -5143 10239
rect 6553 11515 6649 11549
rect 9581 11515 9677 11549
rect 6553 11453 6587 11515
rect -2087 10177 -2053 10239
rect -5177 10143 -5081 10177
rect -2149 10143 -2053 10177
rect -1374 10638 -1278 10672
rect 5112 10638 5208 10672
rect -1374 10576 -1340 10638
rect -3832 10089 -3718 10143
rect -5177 10055 -5081 10089
rect -2149 10055 -2053 10089
rect -5177 9993 -5143 10055
rect -2087 9993 -2053 10055
rect -5177 8717 -5143 8779
rect 5174 10576 5208 10638
rect -1214 10536 -1198 10570
rect -1130 10536 -1114 10570
rect -1056 10536 -1040 10570
rect -972 10536 -956 10570
rect -898 10536 -882 10570
rect -814 10536 -798 10570
rect -740 10536 -724 10570
rect -656 10536 -640 10570
rect -582 10536 -566 10570
rect -498 10536 -482 10570
rect -424 10536 -408 10570
rect -340 10536 -324 10570
rect -266 10536 -250 10570
rect -182 10536 -166 10570
rect -108 10536 -92 10570
rect -24 10536 -8 10570
rect 50 10536 66 10570
rect 134 10536 150 10570
rect 208 10536 224 10570
rect 292 10536 308 10570
rect 366 10536 382 10570
rect 450 10536 466 10570
rect 524 10536 540 10570
rect 608 10536 624 10570
rect 682 10536 698 10570
rect 766 10536 782 10570
rect 840 10536 856 10570
rect 924 10536 940 10570
rect 998 10536 1014 10570
rect 1082 10536 1098 10570
rect 1156 10536 1172 10570
rect 1240 10536 1256 10570
rect 1314 10536 1330 10570
rect 1398 10536 1414 10570
rect 1472 10536 1488 10570
rect 1556 10536 1572 10570
rect 1630 10536 1646 10570
rect 1714 10536 1730 10570
rect 1788 10536 1804 10570
rect 1872 10536 1888 10570
rect 1946 10536 1962 10570
rect 2030 10536 2046 10570
rect 2104 10536 2120 10570
rect 2188 10536 2204 10570
rect 2262 10536 2278 10570
rect 2346 10536 2362 10570
rect 2420 10536 2436 10570
rect 2504 10536 2520 10570
rect 2578 10536 2594 10570
rect 2662 10536 2678 10570
rect 2736 10536 2752 10570
rect 2820 10536 2836 10570
rect 2894 10536 2910 10570
rect 2978 10536 2994 10570
rect 3052 10536 3068 10570
rect 3136 10536 3152 10570
rect 3210 10536 3226 10570
rect 3294 10536 3310 10570
rect 3368 10536 3384 10570
rect 3452 10536 3468 10570
rect 3526 10536 3542 10570
rect 3610 10536 3626 10570
rect 3684 10536 3700 10570
rect 3768 10536 3784 10570
rect 3842 10536 3858 10570
rect 3926 10536 3942 10570
rect 4000 10536 4016 10570
rect 4084 10536 4100 10570
rect 4158 10536 4174 10570
rect 4242 10536 4258 10570
rect 4316 10536 4332 10570
rect 4400 10536 4416 10570
rect 4474 10536 4490 10570
rect 4558 10536 4574 10570
rect 4632 10536 4648 10570
rect 4716 10536 4732 10570
rect 4790 10536 4806 10570
rect 4874 10536 4890 10570
rect 4948 10536 4964 10570
rect 5032 10536 5048 10570
rect -1260 10477 -1226 10493
rect -1260 9485 -1226 9501
rect -1102 10477 -1068 10493
rect -1102 9485 -1068 9501
rect -944 10477 -910 10493
rect -944 9485 -910 9501
rect -786 10477 -752 10493
rect -786 9485 -752 9501
rect -628 10477 -594 10493
rect -628 9485 -594 9501
rect -470 10477 -436 10493
rect -470 9485 -436 9501
rect -312 10477 -278 10493
rect -312 9485 -278 9501
rect -154 10477 -120 10493
rect -154 9485 -120 9501
rect 4 10477 38 10493
rect 4 9485 38 9501
rect 162 10477 196 10493
rect 162 9485 196 9501
rect 320 10477 354 10493
rect 320 9485 354 9501
rect 478 10477 512 10493
rect 478 9485 512 9501
rect 636 10477 670 10493
rect 636 9485 670 9501
rect 794 10477 828 10493
rect 794 9485 828 9501
rect 952 10477 986 10493
rect 952 9485 986 9501
rect 1110 10477 1144 10493
rect 1110 9485 1144 9501
rect 1268 10477 1302 10493
rect 1268 9485 1302 9501
rect 1426 10477 1460 10493
rect 1426 9485 1460 9501
rect 1584 10477 1618 10493
rect 1584 9485 1618 9501
rect 1742 10477 1776 10493
rect 1742 9485 1776 9501
rect 1900 10477 1934 10493
rect 1900 9485 1934 9501
rect 2058 10477 2092 10493
rect 2058 9485 2092 9501
rect 2216 10477 2250 10493
rect 2216 9485 2250 9501
rect 2374 10477 2408 10493
rect 2374 9485 2408 9501
rect 2532 10477 2566 10493
rect 2532 9485 2566 9501
rect 2690 10477 2724 10493
rect 2690 9485 2724 9501
rect 2848 10477 2882 10493
rect 2848 9485 2882 9501
rect 3006 10477 3040 10493
rect 3006 9485 3040 9501
rect 3164 10477 3198 10493
rect 3164 9485 3198 9501
rect 3322 10477 3356 10493
rect 3322 9485 3356 9501
rect 3480 10477 3514 10493
rect 3480 9485 3514 9501
rect 3638 10477 3672 10493
rect 3638 9485 3672 9501
rect 3796 10477 3830 10493
rect 3796 9485 3830 9501
rect 3954 10477 3988 10493
rect 3954 9485 3988 9501
rect 4112 10477 4146 10493
rect 4112 9485 4146 9501
rect 4270 10477 4304 10493
rect 4270 9485 4304 9501
rect 4428 10477 4462 10493
rect 4428 9485 4462 9501
rect 4586 10477 4620 10493
rect 4586 9485 4620 9501
rect 4744 10477 4778 10493
rect 4744 9485 4778 9501
rect 4902 10477 4936 10493
rect 4902 9485 4936 9501
rect 5060 10477 5094 10493
rect 5060 9485 5094 9501
rect -1214 9408 -1198 9442
rect -1130 9408 -1114 9442
rect -1056 9408 -1040 9442
rect -972 9408 -956 9442
rect -898 9408 -882 9442
rect -814 9408 -798 9442
rect -740 9408 -724 9442
rect -656 9408 -640 9442
rect -582 9408 -566 9442
rect -498 9408 -482 9442
rect -424 9408 -408 9442
rect -340 9408 -324 9442
rect -266 9408 -250 9442
rect -182 9408 -166 9442
rect -108 9408 -92 9442
rect -24 9408 -8 9442
rect 50 9408 66 9442
rect 134 9408 150 9442
rect 208 9408 224 9442
rect 292 9408 308 9442
rect 366 9408 382 9442
rect 450 9408 466 9442
rect 524 9408 540 9442
rect 608 9408 624 9442
rect 682 9408 698 9442
rect 766 9408 782 9442
rect 840 9408 856 9442
rect 924 9408 940 9442
rect 998 9408 1014 9442
rect 1082 9408 1098 9442
rect 1156 9408 1172 9442
rect 1240 9408 1256 9442
rect 1314 9408 1330 9442
rect 1398 9408 1414 9442
rect 1472 9408 1488 9442
rect 1556 9408 1572 9442
rect 1630 9408 1646 9442
rect 1714 9408 1730 9442
rect 1788 9408 1804 9442
rect 1872 9408 1888 9442
rect 1946 9408 1962 9442
rect 2030 9408 2046 9442
rect 2104 9408 2120 9442
rect 2188 9408 2204 9442
rect 2262 9408 2278 9442
rect 2346 9408 2362 9442
rect 2420 9408 2436 9442
rect 2504 9408 2520 9442
rect 2578 9408 2594 9442
rect 2662 9408 2678 9442
rect 2736 9408 2752 9442
rect 2820 9408 2836 9442
rect 2894 9408 2910 9442
rect 2978 9408 2994 9442
rect 3052 9408 3068 9442
rect 3136 9408 3152 9442
rect 3210 9408 3226 9442
rect 3294 9408 3310 9442
rect 3368 9408 3384 9442
rect 3452 9408 3468 9442
rect 3526 9408 3542 9442
rect 3610 9408 3626 9442
rect 3684 9408 3700 9442
rect 3768 9408 3784 9442
rect 3842 9408 3858 9442
rect 3926 9408 3942 9442
rect 4000 9408 4016 9442
rect 4084 9408 4100 9442
rect 4158 9408 4174 9442
rect 4242 9408 4258 9442
rect 4316 9408 4332 9442
rect 4400 9408 4416 9442
rect 4474 9408 4490 9442
rect 4558 9408 4574 9442
rect 4632 9408 4648 9442
rect 4716 9408 4732 9442
rect 4790 9408 4806 9442
rect 4874 9408 4890 9442
rect 4948 9408 4964 9442
rect 5032 9408 5048 9442
rect -1374 9340 -1340 9402
rect 9643 11453 9677 11515
rect 6553 10177 6587 10239
rect 9643 10177 9677 10239
rect 6553 10143 6649 10177
rect 9581 10143 9677 10177
rect 7832 10089 8034 10143
rect 5174 9340 5208 9402
rect -1374 9306 -1278 9340
rect 5112 9306 5208 9340
rect 6553 10055 6649 10089
rect 9581 10055 9677 10089
rect 6553 9993 6587 10055
rect -2087 8717 -2053 8779
rect -5177 8683 -5081 8717
rect -2149 8683 -2053 8717
rect 126 8968 222 9002
rect 3610 8968 3706 9002
rect 126 8906 160 8968
rect -4610 8220 -4480 8236
rect -4610 8044 -4480 8060
rect -2940 8230 -2810 8246
rect -2940 8054 -2810 8070
rect 3672 8906 3706 8968
rect 286 8866 302 8900
rect 370 8866 386 8900
rect 444 8866 460 8900
rect 528 8866 544 8900
rect 602 8866 618 8900
rect 686 8866 702 8900
rect 760 8866 776 8900
rect 844 8866 860 8900
rect 918 8866 934 8900
rect 1002 8866 1018 8900
rect 1076 8866 1092 8900
rect 1160 8866 1176 8900
rect 1234 8866 1250 8900
rect 1318 8866 1334 8900
rect 1392 8866 1408 8900
rect 1476 8866 1492 8900
rect 1550 8866 1566 8900
rect 1634 8866 1650 8900
rect 1708 8866 1724 8900
rect 1792 8866 1808 8900
rect 1866 8866 1882 8900
rect 1950 8866 1966 8900
rect 2024 8866 2040 8900
rect 2108 8866 2124 8900
rect 2182 8866 2198 8900
rect 2266 8866 2282 8900
rect 2340 8866 2356 8900
rect 2424 8866 2440 8900
rect 2498 8866 2514 8900
rect 2582 8866 2598 8900
rect 2656 8866 2672 8900
rect 2740 8866 2756 8900
rect 2814 8866 2830 8900
rect 2898 8866 2914 8900
rect 2972 8866 2988 8900
rect 3056 8866 3072 8900
rect 3130 8866 3146 8900
rect 3214 8866 3230 8900
rect 3288 8866 3304 8900
rect 3372 8866 3388 8900
rect 3446 8866 3462 8900
rect 3530 8866 3546 8900
rect 240 8807 274 8823
rect 240 7815 274 7831
rect 398 8807 432 8823
rect 398 7815 432 7831
rect 556 8807 590 8823
rect 556 7815 590 7831
rect 714 8807 748 8823
rect 714 7815 748 7831
rect 872 8807 906 8823
rect 872 7815 906 7831
rect 1030 8807 1064 8823
rect 1030 7815 1064 7831
rect 1188 8807 1222 8823
rect 1188 7815 1222 7831
rect 1346 8807 1380 8823
rect 1346 7815 1380 7831
rect 1504 8807 1538 8823
rect 1504 7815 1538 7831
rect 1662 8807 1696 8823
rect 1662 7815 1696 7831
rect 1820 8807 1854 8823
rect 1820 7815 1854 7831
rect 1978 8807 2012 8823
rect 1978 7815 2012 7831
rect 2136 8807 2170 8823
rect 2136 7815 2170 7831
rect 2294 8807 2328 8823
rect 2294 7815 2328 7831
rect 2452 8807 2486 8823
rect 2452 7815 2486 7831
rect 2610 8807 2644 8823
rect 2610 7815 2644 7831
rect 2768 8807 2802 8823
rect 2768 7815 2802 7831
rect 2926 8807 2960 8823
rect 2926 7815 2960 7831
rect 3084 8807 3118 8823
rect 3084 7815 3118 7831
rect 3242 8807 3276 8823
rect 3242 7815 3276 7831
rect 3400 8807 3434 8823
rect 3400 7815 3434 7831
rect 3558 8807 3592 8823
rect 3558 7815 3592 7831
rect 286 7738 302 7772
rect 370 7738 386 7772
rect 444 7738 460 7772
rect 528 7738 544 7772
rect 602 7738 618 7772
rect 686 7738 702 7772
rect 760 7738 776 7772
rect 844 7738 860 7772
rect 918 7738 934 7772
rect 1002 7738 1018 7772
rect 1076 7738 1092 7772
rect 1160 7738 1176 7772
rect 1234 7738 1250 7772
rect 1318 7738 1334 7772
rect 1392 7738 1408 7772
rect 1476 7738 1492 7772
rect 1550 7738 1566 7772
rect 1634 7738 1650 7772
rect 1708 7738 1724 7772
rect 1792 7738 1808 7772
rect 1866 7738 1882 7772
rect 1950 7738 1966 7772
rect 2024 7738 2040 7772
rect 2108 7738 2124 7772
rect 2182 7738 2198 7772
rect 2266 7738 2282 7772
rect 2340 7738 2356 7772
rect 2424 7738 2440 7772
rect 2498 7738 2514 7772
rect 2582 7738 2598 7772
rect 2656 7738 2672 7772
rect 2740 7738 2756 7772
rect 2814 7738 2830 7772
rect 2898 7738 2914 7772
rect 2972 7738 2988 7772
rect 3056 7738 3072 7772
rect 3130 7738 3146 7772
rect 3214 7738 3230 7772
rect 3288 7738 3304 7772
rect 3372 7738 3388 7772
rect 3446 7738 3462 7772
rect 3530 7738 3546 7772
rect 126 7670 160 7732
rect 9643 9993 9677 10055
rect 6553 8717 6587 8779
rect 9643 8717 9677 8779
rect 6553 8683 6649 8717
rect 9581 8683 9677 8717
rect 7010 8360 7120 8376
rect 7010 8214 7120 8230
rect 8890 8350 9000 8366
rect 8890 8204 9000 8220
rect 3672 7670 3706 7732
rect 126 7636 222 7670
rect 3610 7636 3706 7670
rect 126 7428 222 7462
rect 3610 7428 3706 7462
rect 126 7366 160 7428
rect 3672 7366 3706 7428
rect 286 7326 302 7360
rect 370 7326 386 7360
rect 444 7326 460 7360
rect 528 7326 544 7360
rect 602 7326 618 7360
rect 686 7326 702 7360
rect 760 7326 776 7360
rect 844 7326 860 7360
rect 918 7326 934 7360
rect 1002 7326 1018 7360
rect 1076 7326 1092 7360
rect 1160 7326 1176 7360
rect 1234 7326 1250 7360
rect 1318 7326 1334 7360
rect 1392 7326 1408 7360
rect 1476 7326 1492 7360
rect 1550 7326 1566 7360
rect 1634 7326 1650 7360
rect 1708 7326 1724 7360
rect 1792 7326 1808 7360
rect 1866 7326 1882 7360
rect 1950 7326 1966 7360
rect 2024 7326 2040 7360
rect 2108 7326 2124 7360
rect 2182 7326 2198 7360
rect 2266 7326 2282 7360
rect 2340 7326 2356 7360
rect 2424 7326 2440 7360
rect 2498 7326 2514 7360
rect 2582 7326 2598 7360
rect 2656 7326 2672 7360
rect 2740 7326 2756 7360
rect 2814 7326 2830 7360
rect 2898 7326 2914 7360
rect 2972 7326 2988 7360
rect 3056 7326 3072 7360
rect 3130 7326 3146 7360
rect 3214 7326 3230 7360
rect 3288 7326 3304 7360
rect 3372 7326 3388 7360
rect 3446 7326 3462 7360
rect 3530 7326 3546 7360
rect 240 7267 274 7283
rect 240 6275 274 6291
rect 398 7267 432 7283
rect 398 6275 432 6291
rect 556 7267 590 7283
rect 556 6275 590 6291
rect 714 7267 748 7283
rect 714 6275 748 6291
rect 872 7267 906 7283
rect 872 6275 906 6291
rect 1030 7267 1064 7283
rect 1030 6275 1064 6291
rect 1188 7267 1222 7283
rect 1188 6275 1222 6291
rect 1346 7267 1380 7283
rect 1346 6275 1380 6291
rect 1504 7267 1538 7283
rect 1504 6275 1538 6291
rect 1662 7267 1696 7283
rect 1662 6275 1696 6291
rect 1820 7267 1854 7283
rect 1820 6275 1854 6291
rect 1978 7267 2012 7283
rect 1978 6275 2012 6291
rect 2136 7267 2170 7283
rect 2136 6275 2170 6291
rect 2294 7267 2328 7283
rect 2294 6275 2328 6291
rect 2452 7267 2486 7283
rect 2452 6275 2486 6291
rect 2610 7267 2644 7283
rect 2610 6275 2644 6291
rect 2768 7267 2802 7283
rect 2768 6275 2802 6291
rect 2926 7267 2960 7283
rect 2926 6275 2960 6291
rect 3084 7267 3118 7283
rect 3084 6275 3118 6291
rect 3242 7267 3276 7283
rect 3242 6275 3276 6291
rect 3400 7267 3434 7283
rect 3400 6275 3434 6291
rect 3558 7267 3592 7283
rect 3558 6275 3592 6291
rect 286 6198 302 6232
rect 370 6198 386 6232
rect 444 6198 460 6232
rect 528 6198 544 6232
rect 602 6198 618 6232
rect 686 6198 702 6232
rect 760 6198 776 6232
rect 844 6198 860 6232
rect 918 6198 934 6232
rect 1002 6198 1018 6232
rect 1076 6198 1092 6232
rect 1160 6198 1176 6232
rect 1234 6198 1250 6232
rect 1318 6198 1334 6232
rect 1392 6198 1408 6232
rect 1476 6198 1492 6232
rect 1550 6198 1566 6232
rect 1634 6198 1650 6232
rect 1708 6198 1724 6232
rect 1792 6198 1808 6232
rect 1866 6198 1882 6232
rect 1950 6198 1966 6232
rect 2024 6198 2040 6232
rect 2108 6198 2124 6232
rect 2182 6198 2198 6232
rect 2266 6198 2282 6232
rect 2340 6198 2356 6232
rect 2424 6198 2440 6232
rect 2498 6198 2514 6232
rect 2582 6198 2598 6232
rect 2656 6198 2672 6232
rect 2740 6198 2756 6232
rect 2814 6198 2830 6232
rect 2898 6198 2914 6232
rect 2972 6198 2988 6232
rect 3056 6198 3072 6232
rect 3130 6198 3146 6232
rect 3214 6198 3230 6232
rect 3288 6198 3304 6232
rect 3372 6198 3388 6232
rect 3446 6198 3462 6232
rect 3530 6198 3546 6232
rect 126 6130 160 6192
rect 3672 6130 3706 6192
rect 126 6096 222 6130
rect 3610 6096 3706 6130
rect 1227 5851 1323 5885
rect 2499 5851 2595 5885
rect 1227 5789 1261 5851
rect 2561 5789 2595 5851
rect 1387 5749 1403 5783
rect 1471 5749 1487 5783
rect 1545 5749 1561 5783
rect 1629 5749 1645 5783
rect 1703 5749 1719 5783
rect 1787 5749 1803 5783
rect 1861 5749 1877 5783
rect 1945 5749 1961 5783
rect 2019 5749 2035 5783
rect 2103 5749 2119 5783
rect 2177 5749 2193 5783
rect 2261 5749 2277 5783
rect 2335 5749 2351 5783
rect 2419 5749 2435 5783
rect 1341 5699 1375 5715
rect 1341 4707 1375 4723
rect 1499 5699 1533 5715
rect 1499 4707 1533 4723
rect 1657 5699 1691 5715
rect 1657 4707 1691 4723
rect 1815 5699 1849 5715
rect 1815 4707 1849 4723
rect 1973 5699 2007 5715
rect 1973 4707 2007 4723
rect 2131 5699 2165 5715
rect 2131 4707 2165 4723
rect 2289 5699 2323 5715
rect 2289 4707 2323 4723
rect 2447 5699 2481 5715
rect 2447 4707 2481 4723
rect 1387 4639 1403 4673
rect 1471 4639 1487 4673
rect 1545 4639 1561 4673
rect 1629 4639 1645 4673
rect 1703 4639 1719 4673
rect 1787 4639 1803 4673
rect 1861 4639 1877 4673
rect 1945 4639 1961 4673
rect 2019 4639 2035 4673
rect 2103 4639 2119 4673
rect 2177 4639 2193 4673
rect 2261 4639 2277 4673
rect 2335 4639 2351 4673
rect 2419 4639 2435 4673
rect 1227 4571 1261 4633
rect 2561 4571 2595 4633
rect 1227 4537 1323 4571
rect 2499 4537 2595 4571
rect 1227 4331 1323 4365
rect 2499 4331 2595 4365
rect 1227 4269 1261 4331
rect 2561 4269 2595 4331
rect 1387 4229 1403 4263
rect 1471 4229 1487 4263
rect 1545 4229 1561 4263
rect 1629 4229 1645 4263
rect 1703 4229 1719 4263
rect 1787 4229 1803 4263
rect 1861 4229 1877 4263
rect 1945 4229 1961 4263
rect 2019 4229 2035 4263
rect 2103 4229 2119 4263
rect 2177 4229 2193 4263
rect 2261 4229 2277 4263
rect 2335 4229 2351 4263
rect 2419 4229 2435 4263
rect 1341 4179 1375 4195
rect 1341 3187 1375 3203
rect 1499 4179 1533 4195
rect 1499 3187 1533 3203
rect 1657 4179 1691 4195
rect 1657 3187 1691 3203
rect 1815 4179 1849 4195
rect 1815 3187 1849 3203
rect 1973 4179 2007 4195
rect 1973 3187 2007 3203
rect 2131 4179 2165 4195
rect 2131 3187 2165 3203
rect 2289 4179 2323 4195
rect 2289 3187 2323 3203
rect 2447 4179 2481 4195
rect 2447 3187 2481 3203
rect 1387 3119 1403 3153
rect 1471 3119 1487 3153
rect 1545 3119 1561 3153
rect 1629 3119 1645 3153
rect 1703 3119 1719 3153
rect 1787 3119 1803 3153
rect 1861 3119 1877 3153
rect 1945 3119 1961 3153
rect 2019 3119 2035 3153
rect 2103 3119 2119 3153
rect 2177 3119 2193 3153
rect 2261 3119 2277 3153
rect 2335 3119 2351 3153
rect 2419 3119 2435 3153
rect 1227 3051 1261 3113
rect 2561 3051 2595 3113
rect 1227 3017 1323 3051
rect 2499 3017 2595 3051
rect 236 2810 332 2844
rect 3498 2810 3594 2844
rect 236 2748 270 2810
rect 3560 2748 3594 2810
rect 396 2708 412 2742
rect 580 2708 596 2742
rect 654 2708 670 2742
rect 838 2708 854 2742
rect 912 2708 928 2742
rect 1096 2708 1112 2742
rect 1170 2708 1186 2742
rect 1354 2708 1370 2742
rect 1428 2708 1444 2742
rect 1612 2708 1628 2742
rect 1686 2708 1702 2742
rect 1870 2708 1886 2742
rect 1944 2708 1960 2742
rect 2128 2708 2144 2742
rect 2202 2708 2218 2742
rect 2386 2708 2402 2742
rect 2460 2708 2476 2742
rect 2644 2708 2660 2742
rect 2718 2708 2734 2742
rect 2902 2708 2918 2742
rect 2976 2708 2992 2742
rect 3160 2708 3176 2742
rect 3234 2708 3250 2742
rect 3418 2708 3434 2742
rect 350 2658 384 2674
rect 350 1666 384 1682
rect 608 2658 642 2674
rect 608 1666 642 1682
rect 866 2658 900 2674
rect 866 1666 900 1682
rect 1124 2658 1158 2674
rect 1124 1666 1158 1682
rect 1382 2658 1416 2674
rect 1382 1666 1416 1682
rect 1640 2658 1674 2674
rect 1640 1666 1674 1682
rect 1898 2658 1932 2674
rect 1898 1666 1932 1682
rect 2156 2658 2190 2674
rect 2156 1666 2190 1682
rect 2414 2658 2448 2674
rect 2414 1666 2448 1682
rect 2672 2658 2706 2674
rect 2672 1666 2706 1682
rect 2930 2658 2964 2674
rect 2930 1666 2964 1682
rect 3188 2658 3222 2674
rect 3188 1666 3222 1682
rect 3446 2658 3480 2674
rect 3446 1666 3480 1682
rect 396 1598 412 1632
rect 580 1598 596 1632
rect 654 1598 670 1632
rect 838 1598 854 1632
rect 912 1598 928 1632
rect 1096 1598 1112 1632
rect 1170 1598 1186 1632
rect 1354 1598 1370 1632
rect 1428 1598 1444 1632
rect 1612 1598 1628 1632
rect 1686 1598 1702 1632
rect 1870 1598 1886 1632
rect 1944 1598 1960 1632
rect 2128 1598 2144 1632
rect 2202 1598 2218 1632
rect 2386 1598 2402 1632
rect 2460 1598 2476 1632
rect 2644 1598 2660 1632
rect 2718 1598 2734 1632
rect 2902 1598 2918 1632
rect 2976 1598 2992 1632
rect 3160 1598 3176 1632
rect 3234 1598 3250 1632
rect 3418 1598 3434 1632
rect 236 1530 270 1592
rect 3560 1530 3594 1592
rect 236 1496 332 1530
rect 3498 1496 3594 1530
rect -24 1290 72 1324
rect 3754 1290 3850 1324
rect -24 1228 10 1290
rect 3816 1228 3850 1290
rect 136 1188 152 1222
rect 320 1188 336 1222
rect 394 1188 410 1222
rect 578 1188 594 1222
rect 652 1188 668 1222
rect 836 1188 852 1222
rect 910 1188 926 1222
rect 1094 1188 1110 1222
rect 1168 1188 1184 1222
rect 1352 1188 1368 1222
rect 1426 1188 1442 1222
rect 1610 1188 1626 1222
rect 1684 1188 1700 1222
rect 1868 1188 1884 1222
rect 1942 1188 1958 1222
rect 2126 1188 2142 1222
rect 2200 1188 2216 1222
rect 2384 1188 2400 1222
rect 2458 1188 2474 1222
rect 2642 1188 2658 1222
rect 2716 1188 2732 1222
rect 2900 1188 2916 1222
rect 2974 1188 2990 1222
rect 3158 1188 3174 1222
rect 3232 1188 3248 1222
rect 3416 1188 3432 1222
rect 3490 1188 3506 1222
rect 3674 1188 3690 1222
rect 90 1138 124 1154
rect 90 146 124 162
rect 348 1138 382 1154
rect 348 146 382 162
rect 606 1138 640 1154
rect 606 146 640 162
rect 864 1138 898 1154
rect 864 146 898 162
rect 1122 1138 1156 1154
rect 1122 146 1156 162
rect 1380 1138 1414 1154
rect 1380 146 1414 162
rect 1638 1138 1672 1154
rect 1638 146 1672 162
rect 1896 1138 1930 1154
rect 1896 146 1930 162
rect 2154 1138 2188 1154
rect 2154 146 2188 162
rect 2412 1138 2446 1154
rect 2412 146 2446 162
rect 2670 1138 2704 1154
rect 2670 146 2704 162
rect 2928 1138 2962 1154
rect 2928 146 2962 162
rect 3186 1138 3220 1154
rect 3186 146 3220 162
rect 3444 1138 3478 1154
rect 3444 146 3478 162
rect 3702 1138 3736 1154
rect 3702 146 3736 162
rect 136 78 152 112
rect 320 78 336 112
rect 394 78 410 112
rect 578 78 594 112
rect 652 78 668 112
rect 836 78 852 112
rect 910 78 926 112
rect 1094 78 1110 112
rect 1168 78 1184 112
rect 1352 78 1368 112
rect 1426 78 1442 112
rect 1610 78 1626 112
rect 1684 78 1700 112
rect 1868 78 1884 112
rect 1942 78 1958 112
rect 2126 78 2142 112
rect 2200 78 2216 112
rect 2384 78 2400 112
rect 2458 78 2474 112
rect 2642 78 2658 112
rect 2716 78 2732 112
rect 2900 78 2916 112
rect 2974 78 2990 112
rect 3158 78 3174 112
rect 3232 78 3248 112
rect 3416 78 3432 112
rect 3490 78 3506 112
rect 3674 78 3690 112
rect -24 10 10 72
rect 3816 10 3850 72
rect -24 -24 72 10
rect 3754 -24 3850 10
<< viali >>
rect -5029 10289 -4632 11403
rect -2598 10289 -2201 11403
rect 289 10638 3545 10672
rect -5029 8829 -4632 9943
rect -2598 8829 -2201 9943
rect -1198 10536 -1130 10570
rect -1040 10536 -972 10570
rect -882 10536 -814 10570
rect -724 10536 -656 10570
rect -566 10536 -498 10570
rect -408 10536 -340 10570
rect -250 10536 -182 10570
rect -92 10536 -24 10570
rect 66 10536 134 10570
rect 224 10536 292 10570
rect 382 10536 450 10570
rect 540 10536 608 10570
rect 698 10536 766 10570
rect 856 10536 924 10570
rect 1014 10536 1082 10570
rect 1172 10536 1240 10570
rect 1330 10536 1398 10570
rect 1488 10536 1556 10570
rect 1646 10536 1714 10570
rect 1804 10536 1872 10570
rect 1962 10536 2030 10570
rect 2120 10536 2188 10570
rect 2278 10536 2346 10570
rect 2436 10536 2504 10570
rect 2594 10536 2662 10570
rect 2752 10536 2820 10570
rect 2910 10536 2978 10570
rect 3068 10536 3136 10570
rect 3226 10536 3294 10570
rect 3384 10536 3452 10570
rect 3542 10536 3610 10570
rect 3700 10536 3768 10570
rect 3858 10536 3926 10570
rect 4016 10536 4084 10570
rect 4174 10536 4242 10570
rect 4332 10536 4400 10570
rect 4490 10536 4558 10570
rect 4648 10536 4716 10570
rect 4806 10536 4874 10570
rect 4964 10536 5032 10570
rect -1260 9501 -1226 10477
rect -1102 9501 -1068 10477
rect -944 9501 -910 10477
rect -786 9501 -752 10477
rect -628 9501 -594 10477
rect -470 9501 -436 10477
rect -312 9501 -278 10477
rect -154 9501 -120 10477
rect 4 9501 38 10477
rect 162 9501 196 10477
rect 320 9501 354 10477
rect 478 9501 512 10477
rect 636 9501 670 10477
rect 794 9501 828 10477
rect 952 9501 986 10477
rect 1110 9501 1144 10477
rect 1268 9501 1302 10477
rect 1426 9501 1460 10477
rect 1584 9501 1618 10477
rect 1742 9501 1776 10477
rect 1900 9501 1934 10477
rect 2058 9501 2092 10477
rect 2216 9501 2250 10477
rect 2374 9501 2408 10477
rect 2532 9501 2566 10477
rect 2690 9501 2724 10477
rect 2848 9501 2882 10477
rect 3006 9501 3040 10477
rect 3164 9501 3198 10477
rect 3322 9501 3356 10477
rect 3480 9501 3514 10477
rect 3638 9501 3672 10477
rect 3796 9501 3830 10477
rect 3954 9501 3988 10477
rect 4112 9501 4146 10477
rect 4270 9501 4304 10477
rect 4428 9501 4462 10477
rect 4586 9501 4620 10477
rect 4744 9501 4778 10477
rect 4902 9501 4936 10477
rect 5060 9501 5094 10477
rect -1198 9408 -1130 9442
rect -1040 9408 -972 9442
rect -882 9408 -814 9442
rect -724 9408 -656 9442
rect -566 9408 -498 9442
rect -408 9408 -340 9442
rect -250 9408 -182 9442
rect -92 9408 -24 9442
rect 66 9408 134 9442
rect 224 9408 292 9442
rect 382 9408 450 9442
rect 540 9408 608 9442
rect 698 9408 766 9442
rect 856 9408 924 9442
rect 1014 9408 1082 9442
rect 1172 9408 1240 9442
rect 1330 9408 1398 9442
rect 1488 9408 1556 9442
rect 1646 9408 1714 9442
rect 1804 9408 1872 9442
rect 1962 9408 2030 9442
rect 2120 9408 2188 9442
rect 2278 9408 2346 9442
rect 2436 9408 2504 9442
rect 2594 9408 2662 9442
rect 2752 9408 2820 9442
rect 2910 9408 2978 9442
rect 3068 9408 3136 9442
rect 3226 9408 3294 9442
rect 3384 9408 3452 9442
rect 3542 9408 3610 9442
rect 3700 9408 3768 9442
rect 3858 9408 3926 9442
rect 4016 9408 4084 9442
rect 4174 9408 4242 9442
rect 4332 9408 4400 9442
rect 4490 9408 4558 9442
rect 4648 9408 4716 9442
rect 4806 9408 4874 9442
rect 4964 9408 5032 9442
rect 6701 10289 7098 11403
rect 9132 10289 9529 11403
rect 289 9306 3545 9340
rect -3912 8717 -3682 8722
rect -3912 8683 -3682 8717
rect 1038 8968 2794 9002
rect -3912 8636 -3682 8683
rect -4610 8060 -4480 8220
rect -2940 8070 -2810 8230
rect 302 8866 370 8900
rect 460 8866 528 8900
rect 618 8866 686 8900
rect 776 8866 844 8900
rect 934 8866 1002 8900
rect 1092 8866 1160 8900
rect 1250 8866 1318 8900
rect 1408 8866 1476 8900
rect 1566 8866 1634 8900
rect 1724 8866 1792 8900
rect 1882 8866 1950 8900
rect 2040 8866 2108 8900
rect 2198 8866 2266 8900
rect 2356 8866 2424 8900
rect 2514 8866 2582 8900
rect 2672 8866 2740 8900
rect 2830 8866 2898 8900
rect 2988 8866 3056 8900
rect 3146 8866 3214 8900
rect 3304 8866 3372 8900
rect 3462 8866 3530 8900
rect 240 7831 274 8807
rect 398 7831 432 8807
rect 556 7831 590 8807
rect 714 7831 748 8807
rect 872 7831 906 8807
rect 1030 7831 1064 8807
rect 1188 7831 1222 8807
rect 1346 7831 1380 8807
rect 1504 7831 1538 8807
rect 1662 7831 1696 8807
rect 1820 7831 1854 8807
rect 1978 7831 2012 8807
rect 2136 7831 2170 8807
rect 2294 7831 2328 8807
rect 2452 7831 2486 8807
rect 2610 7831 2644 8807
rect 2768 7831 2802 8807
rect 2926 7831 2960 8807
rect 3084 7831 3118 8807
rect 3242 7831 3276 8807
rect 3400 7831 3434 8807
rect 3558 7831 3592 8807
rect 302 7738 370 7772
rect 460 7738 528 7772
rect 618 7738 686 7772
rect 776 7738 844 7772
rect 934 7738 1002 7772
rect 1092 7738 1160 7772
rect 1250 7738 1318 7772
rect 1408 7738 1476 7772
rect 1566 7738 1634 7772
rect 1724 7738 1792 7772
rect 1882 7738 1950 7772
rect 2040 7738 2108 7772
rect 2198 7738 2266 7772
rect 2356 7738 2424 7772
rect 2514 7738 2582 7772
rect 2672 7738 2740 7772
rect 2830 7738 2898 7772
rect 2988 7738 3056 7772
rect 3146 7738 3214 7772
rect 3304 7738 3372 7772
rect 3462 7738 3530 7772
rect 6701 8829 7098 9943
rect 9132 8829 9529 9943
rect 7656 8683 7874 8706
rect 7656 8614 7874 8683
rect 7010 8230 7120 8360
rect 8890 8220 9000 8350
rect 900 7636 1470 7670
rect 2370 7636 2940 7670
rect 900 7462 1470 7636
rect 2370 7462 2940 7636
rect 900 7430 1470 7462
rect 2370 7430 2940 7462
rect 302 7326 370 7360
rect 460 7326 528 7360
rect 618 7326 686 7360
rect 776 7326 844 7360
rect 934 7326 1002 7360
rect 1092 7326 1160 7360
rect 1250 7326 1318 7360
rect 1408 7326 1476 7360
rect 1566 7326 1634 7360
rect 1724 7326 1792 7360
rect 1882 7326 1950 7360
rect 2040 7326 2108 7360
rect 2198 7326 2266 7360
rect 2356 7326 2424 7360
rect 2514 7326 2582 7360
rect 2672 7326 2740 7360
rect 2830 7326 2898 7360
rect 2988 7326 3056 7360
rect 3146 7326 3214 7360
rect 3304 7326 3372 7360
rect 3462 7326 3530 7360
rect 240 6291 274 7267
rect 398 6291 432 7267
rect 556 6291 590 7267
rect 714 6291 748 7267
rect 872 6291 906 7267
rect 1030 6291 1064 7267
rect 1188 6291 1222 7267
rect 1346 6291 1380 7267
rect 1504 6291 1538 7267
rect 1662 6291 1696 7267
rect 1820 6291 1854 7267
rect 1978 6291 2012 7267
rect 2136 6291 2170 7267
rect 2294 6291 2328 7267
rect 2452 6291 2486 7267
rect 2610 6291 2644 7267
rect 2768 6291 2802 7267
rect 2926 6291 2960 7267
rect 3084 6291 3118 7267
rect 3242 6291 3276 7267
rect 3400 6291 3434 7267
rect 3558 6291 3592 7267
rect 302 6198 370 6232
rect 460 6198 528 6232
rect 618 6198 686 6232
rect 776 6198 844 6232
rect 934 6198 1002 6232
rect 1092 6198 1160 6232
rect 1250 6198 1318 6232
rect 1408 6198 1476 6232
rect 1566 6198 1634 6232
rect 1724 6198 1792 6232
rect 1882 6198 1950 6232
rect 2040 6198 2108 6232
rect 2198 6198 2266 6232
rect 2356 6198 2424 6232
rect 2514 6198 2582 6232
rect 2672 6198 2740 6232
rect 2830 6198 2898 6232
rect 2988 6198 3056 6232
rect 3146 6198 3214 6232
rect 3304 6198 3372 6232
rect 3462 6198 3530 6232
rect 1586 5851 2236 5885
rect 1403 5749 1471 5783
rect 1561 5749 1629 5783
rect 1719 5749 1787 5783
rect 1877 5749 1945 5783
rect 2035 5749 2103 5783
rect 2193 5749 2261 5783
rect 2351 5749 2419 5783
rect 1341 4723 1375 5699
rect 1499 4723 1533 5699
rect 1657 4723 1691 5699
rect 1815 4723 1849 5699
rect 1973 4723 2007 5699
rect 2131 4723 2165 5699
rect 2289 4723 2323 5699
rect 2447 4723 2481 5699
rect 1403 4639 1471 4673
rect 1561 4639 1629 4673
rect 1719 4639 1787 4673
rect 1877 4639 1945 4673
rect 2035 4639 2103 4673
rect 2193 4639 2261 4673
rect 2351 4639 2419 4673
rect 1586 4537 2236 4571
rect 1586 4331 2236 4365
rect 1403 4229 1471 4263
rect 1561 4229 1629 4263
rect 1719 4229 1787 4263
rect 1877 4229 1945 4263
rect 2035 4229 2103 4263
rect 2193 4229 2261 4263
rect 2351 4229 2419 4263
rect 1341 3203 1375 4179
rect 1499 3203 1533 4179
rect 1657 3203 1691 4179
rect 1815 3203 1849 4179
rect 1973 3203 2007 4179
rect 2131 3203 2165 4179
rect 2289 3203 2323 4179
rect 2447 3203 2481 4179
rect 1403 3119 1471 3153
rect 1561 3119 1629 3153
rect 1719 3119 1787 3153
rect 1877 3119 1945 3153
rect 2035 3119 2103 3153
rect 2193 3119 2261 3153
rect 2351 3119 2419 3153
rect 1586 3017 2236 3051
rect 1093 2810 2737 2844
rect 412 2708 580 2742
rect 670 2708 838 2742
rect 928 2708 1096 2742
rect 1186 2708 1354 2742
rect 1444 2708 1612 2742
rect 1702 2708 1870 2742
rect 1960 2708 2128 2742
rect 2218 2708 2386 2742
rect 2476 2708 2644 2742
rect 2734 2708 2902 2742
rect 2992 2708 3160 2742
rect 3250 2708 3418 2742
rect 350 1682 384 2658
rect 608 1682 642 2658
rect 866 1682 900 2658
rect 1124 1682 1158 2658
rect 1382 1682 1416 2658
rect 1640 1682 1674 2658
rect 1898 1682 1932 2658
rect 2156 1682 2190 2658
rect 2414 1682 2448 2658
rect 2672 1682 2706 2658
rect 2930 1682 2964 2658
rect 3188 1682 3222 2658
rect 3446 1682 3480 2658
rect 412 1598 580 1632
rect 670 1598 838 1632
rect 928 1598 1096 1632
rect 1186 1598 1354 1632
rect 1444 1598 1612 1632
rect 1702 1598 1870 1632
rect 1960 1598 2128 1632
rect 2218 1598 2386 1632
rect 2476 1598 2644 1632
rect 2734 1598 2902 1632
rect 2992 1598 3160 1632
rect 3250 1598 3418 1632
rect 1093 1496 2737 1530
rect 962 1290 2864 1324
rect 152 1188 320 1222
rect 410 1188 578 1222
rect 668 1188 836 1222
rect 926 1188 1094 1222
rect 1184 1188 1352 1222
rect 1442 1188 1610 1222
rect 1700 1188 1868 1222
rect 1958 1188 2126 1222
rect 2216 1188 2384 1222
rect 2474 1188 2642 1222
rect 2732 1188 2900 1222
rect 2990 1188 3158 1222
rect 3248 1188 3416 1222
rect 3506 1188 3674 1222
rect 90 162 124 1138
rect 348 162 382 1138
rect 606 162 640 1138
rect 864 162 898 1138
rect 1122 162 1156 1138
rect 1380 162 1414 1138
rect 1638 162 1672 1138
rect 1896 162 1930 1138
rect 2154 162 2188 1138
rect 2412 162 2446 1138
rect 2670 162 2704 1138
rect 2928 162 2962 1138
rect 3186 162 3220 1138
rect 3444 162 3478 1138
rect 3702 162 3736 1138
rect 152 78 320 112
rect 410 78 578 112
rect 668 78 836 112
rect 926 78 1094 112
rect 1184 78 1352 112
rect 1442 78 1610 112
rect 1700 78 1868 112
rect 1958 78 2126 112
rect 2216 78 2384 112
rect 2474 78 2642 112
rect 2732 78 2900 112
rect 2990 78 3158 112
rect 3248 78 3416 112
rect 3506 78 3674 112
rect 962 -24 2864 10
<< metal1 >>
rect -5540 11890 -5100 11930
rect -5540 11820 -5390 11890
rect -5320 11820 -5100 11890
rect -5540 11770 -5100 11820
rect -5540 11700 -5390 11770
rect -5320 11700 -5100 11770
rect -5540 11650 -5100 11700
rect -5540 11580 -5390 11650
rect -5320 11580 -5100 11650
rect -5540 11530 -5100 11580
rect -5540 11460 -5390 11530
rect -5320 11460 -5100 11530
rect -5540 11310 -5100 11460
rect 9000 11890 9440 11930
rect 9000 11820 9200 11890
rect 9270 11820 9440 11890
rect 9000 11770 9440 11820
rect 9000 11700 9200 11770
rect 9270 11700 9440 11770
rect 9000 11650 9440 11700
rect 9000 11580 9200 11650
rect 9270 11580 9440 11650
rect 9000 11530 9440 11580
rect 9000 11460 9200 11530
rect 9270 11460 9440 11530
rect 9000 11415 9440 11460
rect -5035 11403 -4626 11415
rect -5035 11310 -5029 11403
rect -5540 10289 -5029 11310
rect -4632 10289 -4626 11403
rect -2604 11403 -2195 11415
rect -2604 11310 -2598 11403
rect -5540 10277 -4626 10289
rect -2730 10289 -2598 11310
rect -2201 10289 -2195 11403
rect 6695 11403 7104 11415
rect 6695 11310 6701 11403
rect 1240 10930 2620 10980
rect 1240 10678 1270 10930
rect 277 10672 1270 10678
rect 1540 10672 2320 10930
rect 2590 10678 2620 10930
rect 2590 10672 3557 10678
rect 277 10638 289 10672
rect 3545 10638 3557 10672
rect 277 10632 3557 10638
rect -2730 10277 -2195 10289
rect -1410 10570 5250 10580
rect -1410 10536 -1198 10570
rect -1130 10536 -1040 10570
rect -972 10536 -882 10570
rect -814 10536 -724 10570
rect -656 10536 -566 10570
rect -498 10536 -408 10570
rect -340 10536 -250 10570
rect -182 10536 -92 10570
rect -24 10536 66 10570
rect 134 10536 224 10570
rect 292 10536 382 10570
rect 450 10536 540 10570
rect 608 10536 698 10570
rect 766 10536 856 10570
rect 924 10536 1014 10570
rect 1082 10536 1172 10570
rect 1240 10536 1330 10570
rect 1398 10536 1488 10570
rect 1556 10536 1646 10570
rect 1714 10536 1804 10570
rect 1872 10536 1962 10570
rect 2030 10536 2120 10570
rect 2188 10536 2278 10570
rect 2346 10536 2436 10570
rect 2504 10536 2594 10570
rect 2662 10536 2752 10570
rect 2820 10536 2910 10570
rect 2978 10536 3068 10570
rect 3136 10536 3226 10570
rect 3294 10536 3384 10570
rect 3452 10536 3542 10570
rect 3610 10536 3700 10570
rect 3768 10536 3858 10570
rect 3926 10536 4016 10570
rect 4084 10536 4174 10570
rect 4242 10536 4332 10570
rect 4400 10536 4490 10570
rect 4558 10536 4648 10570
rect 4716 10536 4806 10570
rect 4874 10536 4964 10570
rect 5032 10536 5250 10570
rect -1410 10530 5250 10536
rect -5540 9955 -4730 10277
rect -2730 10150 -2290 10277
rect -1410 10150 -1330 10530
rect -1266 10477 -1220 10489
rect -1266 10450 -1260 10477
rect -1226 10450 -1220 10477
rect -1108 10477 -1062 10489
rect -1290 10380 -1280 10450
rect -1210 10380 -1200 10450
rect -1266 10210 -1260 10380
rect -1226 10210 -1220 10380
rect -5540 9943 -4626 9955
rect -5540 8829 -5029 9943
rect -4632 8829 -4626 9943
rect -5540 8817 -4626 8829
rect -2730 9943 -1330 10150
rect -1290 10140 -1280 10210
rect -1210 10140 -1200 10210
rect -2730 8829 -2598 9943
rect -2201 9860 -1330 9943
rect -2201 8829 -2195 9860
rect -1410 9450 -1330 9860
rect -1266 9501 -1260 10140
rect -1226 9501 -1220 10140
rect -1108 9840 -1102 10477
rect -1068 9840 -1062 10477
rect -950 10477 -904 10489
rect -950 10450 -944 10477
rect -910 10450 -904 10477
rect -792 10477 -746 10489
rect -970 10380 -960 10450
rect -890 10380 -880 10450
rect -950 10210 -944 10380
rect -910 10210 -904 10380
rect -970 10140 -960 10210
rect -890 10140 -880 10210
rect -1130 9770 -1120 9840
rect -1050 9770 -1040 9840
rect -1108 9600 -1102 9770
rect -1068 9600 -1062 9770
rect -1130 9530 -1120 9600
rect -1050 9530 -1040 9600
rect -1266 9489 -1220 9501
rect -1108 9501 -1102 9530
rect -1068 9501 -1062 9530
rect -1108 9489 -1062 9501
rect -950 9501 -944 10140
rect -910 9501 -904 10140
rect -792 9840 -786 10477
rect -752 9840 -746 10477
rect -634 10477 -588 10489
rect -634 10450 -628 10477
rect -594 10450 -588 10477
rect -476 10477 -430 10489
rect -660 10380 -650 10450
rect -580 10380 -570 10450
rect -634 10210 -628 10380
rect -594 10210 -588 10380
rect -660 10140 -650 10210
rect -580 10140 -570 10210
rect -820 9770 -810 9840
rect -740 9770 -730 9840
rect -792 9600 -786 9770
rect -752 9600 -746 9770
rect -820 9530 -810 9600
rect -740 9530 -730 9600
rect -950 9489 -904 9501
rect -792 9501 -786 9530
rect -752 9501 -746 9530
rect -792 9489 -746 9501
rect -634 9501 -628 10140
rect -594 9501 -588 10140
rect -476 9840 -470 10477
rect -436 9840 -430 10477
rect -318 10477 -272 10489
rect -318 10450 -312 10477
rect -278 10450 -272 10477
rect -160 10477 -114 10489
rect -340 10380 -330 10450
rect -260 10380 -250 10450
rect -318 10210 -312 10380
rect -278 10210 -272 10380
rect -340 10140 -330 10210
rect -260 10140 -250 10210
rect -500 9770 -490 9840
rect -420 9770 -410 9840
rect -476 9600 -470 9770
rect -436 9600 -430 9770
rect -500 9530 -490 9600
rect -420 9530 -410 9600
rect -634 9489 -588 9501
rect -476 9501 -470 9530
rect -436 9501 -430 9530
rect -476 9489 -430 9501
rect -318 9501 -312 10140
rect -278 9501 -272 10140
rect -160 9840 -154 10477
rect -120 9840 -114 10477
rect -2 10477 44 10489
rect -2 10450 4 10477
rect 38 10450 44 10477
rect 156 10477 202 10489
rect -30 10380 -20 10450
rect 50 10380 60 10450
rect -2 10210 4 10380
rect 38 10210 44 10380
rect -30 10140 -20 10210
rect 50 10140 60 10210
rect -180 9770 -170 9840
rect -100 9770 -90 9840
rect -160 9600 -154 9770
rect -120 9600 -114 9770
rect -180 9530 -170 9600
rect -100 9530 -90 9600
rect -318 9489 -272 9501
rect -160 9501 -154 9530
rect -120 9501 -114 9530
rect -160 9489 -114 9501
rect -2 9501 4 10140
rect 38 9501 44 10140
rect 156 9840 162 10477
rect 196 9840 202 10477
rect 314 10477 360 10489
rect 314 10450 320 10477
rect 354 10450 360 10477
rect 472 10477 518 10489
rect 290 10380 300 10450
rect 370 10380 380 10450
rect 314 10210 320 10380
rect 354 10210 360 10380
rect 290 10140 300 10210
rect 370 10140 380 10210
rect 130 9770 140 9840
rect 210 9770 220 9840
rect 156 9600 162 9770
rect 196 9600 202 9770
rect 130 9530 140 9600
rect 210 9530 220 9600
rect -2 9489 44 9501
rect 156 9501 162 9530
rect 196 9501 202 9530
rect 156 9489 202 9501
rect 314 9501 320 10140
rect 354 9501 360 10140
rect 472 9840 478 10477
rect 512 9840 518 10477
rect 630 10477 676 10489
rect 630 10450 636 10477
rect 670 10450 676 10477
rect 788 10477 834 10489
rect 610 10380 620 10450
rect 690 10380 700 10450
rect 630 10210 636 10380
rect 670 10210 676 10380
rect 610 10140 620 10210
rect 690 10140 700 10210
rect 450 9770 460 9840
rect 530 9770 540 9840
rect 472 9600 478 9770
rect 512 9600 518 9770
rect 450 9530 460 9600
rect 530 9530 540 9600
rect 314 9489 360 9501
rect 472 9501 478 9530
rect 512 9501 518 9530
rect 472 9489 518 9501
rect 630 9501 636 10140
rect 670 9501 676 10140
rect 788 9840 794 10477
rect 828 9840 834 10477
rect 946 10477 992 10489
rect 946 10450 952 10477
rect 986 10450 992 10477
rect 1104 10477 1150 10489
rect 920 10380 930 10450
rect 1000 10380 1010 10450
rect 946 10210 952 10380
rect 986 10210 992 10380
rect 920 10140 930 10210
rect 1000 10140 1010 10210
rect 760 9770 770 9840
rect 840 9770 850 9840
rect 788 9600 794 9770
rect 828 9600 834 9770
rect 760 9530 770 9600
rect 840 9530 850 9600
rect 630 9489 676 9501
rect 788 9501 794 9530
rect 828 9501 834 9530
rect 788 9489 834 9501
rect 946 9501 952 10140
rect 986 9501 992 10140
rect 1104 9840 1110 10477
rect 1144 9840 1150 10477
rect 1262 10477 1308 10489
rect 1262 10450 1268 10477
rect 1302 10450 1308 10477
rect 1420 10477 1466 10489
rect 1240 10380 1250 10450
rect 1320 10380 1330 10450
rect 1262 10210 1268 10380
rect 1302 10210 1308 10380
rect 1240 10140 1250 10210
rect 1320 10140 1330 10210
rect 1080 9770 1090 9840
rect 1160 9770 1170 9840
rect 1104 9600 1110 9770
rect 1144 9600 1150 9770
rect 1080 9530 1090 9600
rect 1160 9530 1170 9600
rect 946 9489 992 9501
rect 1104 9501 1110 9530
rect 1144 9501 1150 9530
rect 1104 9489 1150 9501
rect 1262 9501 1268 10140
rect 1302 9501 1308 10140
rect 1420 9840 1426 10477
rect 1460 9840 1466 10477
rect 1578 10477 1624 10489
rect 1578 10450 1584 10477
rect 1618 10450 1624 10477
rect 1736 10477 1782 10489
rect 1560 10380 1570 10450
rect 1640 10380 1650 10450
rect 1578 10210 1584 10380
rect 1618 10210 1624 10380
rect 1560 10140 1570 10210
rect 1640 10140 1650 10210
rect 1400 9770 1410 9840
rect 1480 9770 1490 9840
rect 1420 9600 1426 9770
rect 1460 9600 1466 9770
rect 1400 9530 1410 9600
rect 1480 9530 1490 9600
rect 1262 9489 1308 9501
rect 1420 9501 1426 9530
rect 1460 9501 1466 9530
rect 1420 9489 1466 9501
rect 1578 9501 1584 10140
rect 1618 9501 1624 10140
rect 1736 9840 1742 10477
rect 1776 9840 1782 10477
rect 1894 10477 1940 10489
rect 1894 10450 1900 10477
rect 1934 10450 1940 10477
rect 2052 10477 2098 10489
rect 1870 10380 1880 10450
rect 1950 10380 1960 10450
rect 1894 10210 1900 10380
rect 1934 10210 1940 10380
rect 1870 10140 1880 10210
rect 1950 10140 1960 10210
rect 1710 9770 1720 9840
rect 1790 9770 1800 9840
rect 1736 9600 1742 9770
rect 1776 9600 1782 9770
rect 1710 9530 1720 9600
rect 1790 9530 1800 9600
rect 1578 9489 1624 9501
rect 1736 9501 1742 9530
rect 1776 9501 1782 9530
rect 1736 9489 1782 9501
rect 1894 9501 1900 10140
rect 1934 9501 1940 10140
rect 2052 9840 2058 10477
rect 2092 9840 2098 10477
rect 2210 10477 2256 10489
rect 2210 10450 2216 10477
rect 2250 10450 2256 10477
rect 2368 10477 2414 10489
rect 2190 10380 2200 10450
rect 2270 10380 2280 10450
rect 2210 10210 2216 10380
rect 2250 10210 2256 10380
rect 2190 10140 2200 10210
rect 2270 10140 2280 10210
rect 2030 9770 2040 9840
rect 2110 9770 2120 9840
rect 2052 9600 2058 9770
rect 2092 9600 2098 9770
rect 2030 9530 2040 9600
rect 2110 9530 2120 9600
rect 1894 9489 1940 9501
rect 2052 9501 2058 9530
rect 2092 9501 2098 9530
rect 2052 9489 2098 9501
rect 2210 9501 2216 10140
rect 2250 9501 2256 10140
rect 2368 9840 2374 10477
rect 2408 9840 2414 10477
rect 2526 10477 2572 10489
rect 2526 10450 2532 10477
rect 2566 10450 2572 10477
rect 2684 10477 2730 10489
rect 2500 10380 2510 10450
rect 2580 10380 2590 10450
rect 2526 10210 2532 10380
rect 2566 10210 2572 10380
rect 2500 10140 2510 10210
rect 2580 10140 2590 10210
rect 2350 9770 2360 9840
rect 2430 9770 2440 9840
rect 2368 9600 2374 9770
rect 2408 9600 2414 9770
rect 2350 9530 2360 9600
rect 2430 9530 2440 9600
rect 2210 9489 2256 9501
rect 2368 9501 2374 9530
rect 2408 9501 2414 9530
rect 2368 9489 2414 9501
rect 2526 9501 2532 10140
rect 2566 9501 2572 10140
rect 2684 9840 2690 10477
rect 2724 9840 2730 10477
rect 2842 10477 2888 10489
rect 2842 10450 2848 10477
rect 2882 10450 2888 10477
rect 3000 10477 3046 10489
rect 2820 10380 2830 10450
rect 2900 10380 2910 10450
rect 2842 10210 2848 10380
rect 2882 10210 2888 10380
rect 2820 10140 2830 10210
rect 2900 10140 2910 10210
rect 2660 9770 2670 9840
rect 2740 9770 2750 9840
rect 2684 9600 2690 9770
rect 2724 9600 2730 9770
rect 2660 9530 2670 9600
rect 2740 9530 2750 9600
rect 2526 9489 2572 9501
rect 2684 9501 2690 9530
rect 2724 9501 2730 9530
rect 2684 9489 2730 9501
rect 2842 9501 2848 10140
rect 2882 9501 2888 10140
rect 3000 9840 3006 10477
rect 3040 9840 3046 10477
rect 3158 10477 3204 10489
rect 3158 10450 3164 10477
rect 3198 10450 3204 10477
rect 3316 10477 3362 10489
rect 3140 10380 3150 10450
rect 3220 10380 3230 10450
rect 3158 10210 3164 10380
rect 3198 10210 3204 10380
rect 3140 10140 3150 10210
rect 3220 10140 3230 10210
rect 2980 9770 2990 9840
rect 3060 9770 3070 9840
rect 3000 9600 3006 9770
rect 3040 9600 3046 9770
rect 2980 9530 2990 9600
rect 3060 9530 3070 9600
rect 2842 9489 2888 9501
rect 3000 9501 3006 9530
rect 3040 9501 3046 9530
rect 3000 9489 3046 9501
rect 3158 9501 3164 10140
rect 3198 9501 3204 10140
rect 3316 9840 3322 10477
rect 3356 9840 3362 10477
rect 3474 10477 3520 10489
rect 3474 10450 3480 10477
rect 3514 10450 3520 10477
rect 3632 10477 3678 10489
rect 3450 10380 3460 10450
rect 3530 10380 3540 10450
rect 3474 10210 3480 10380
rect 3514 10210 3520 10380
rect 3450 10140 3460 10210
rect 3530 10140 3540 10210
rect 3290 9770 3300 9840
rect 3370 9770 3380 9840
rect 3316 9600 3322 9770
rect 3356 9600 3362 9770
rect 3290 9530 3300 9600
rect 3370 9530 3380 9600
rect 3158 9489 3204 9501
rect 3316 9501 3322 9530
rect 3356 9501 3362 9530
rect 3316 9489 3362 9501
rect 3474 9501 3480 10140
rect 3514 9501 3520 10140
rect 3632 9840 3638 10477
rect 3672 9840 3678 10477
rect 3790 10477 3836 10489
rect 3790 10450 3796 10477
rect 3830 10450 3836 10477
rect 3948 10477 3994 10489
rect 3770 10380 3780 10450
rect 3850 10380 3860 10450
rect 3790 10210 3796 10380
rect 3830 10210 3836 10380
rect 3770 10140 3780 10210
rect 3850 10140 3860 10210
rect 3610 9770 3620 9840
rect 3690 9770 3700 9840
rect 3632 9600 3638 9770
rect 3672 9600 3678 9770
rect 3610 9530 3620 9600
rect 3690 9530 3700 9600
rect 3474 9489 3520 9501
rect 3632 9501 3638 9530
rect 3672 9501 3678 9530
rect 3632 9489 3678 9501
rect 3790 9501 3796 10140
rect 3830 9501 3836 10140
rect 3948 9840 3954 10477
rect 3988 9840 3994 10477
rect 4106 10477 4152 10489
rect 4106 10450 4112 10477
rect 4146 10450 4152 10477
rect 4264 10477 4310 10489
rect 4080 10380 4090 10450
rect 4160 10380 4170 10450
rect 4106 10210 4112 10380
rect 4146 10210 4152 10380
rect 4080 10140 4090 10210
rect 4160 10140 4170 10210
rect 3930 9770 3940 9840
rect 4010 9770 4020 9840
rect 3948 9600 3954 9770
rect 3988 9600 3994 9770
rect 3930 9530 3940 9600
rect 4010 9530 4020 9600
rect 3790 9489 3836 9501
rect 3948 9501 3954 9530
rect 3988 9501 3994 9530
rect 3948 9489 3994 9501
rect 4106 9501 4112 10140
rect 4146 9501 4152 10140
rect 4264 9840 4270 10477
rect 4304 9840 4310 10477
rect 4422 10477 4468 10489
rect 4422 10450 4428 10477
rect 4462 10450 4468 10477
rect 4580 10477 4626 10489
rect 4400 10380 4410 10450
rect 4480 10380 4490 10450
rect 4422 10210 4428 10380
rect 4462 10210 4468 10380
rect 4400 10140 4410 10210
rect 4480 10140 4490 10210
rect 4240 9770 4250 9840
rect 4320 9770 4330 9840
rect 4264 9600 4270 9770
rect 4304 9600 4310 9770
rect 4240 9530 4250 9600
rect 4320 9530 4330 9600
rect 4106 9489 4152 9501
rect 4264 9501 4270 9530
rect 4304 9501 4310 9530
rect 4264 9489 4310 9501
rect 4422 9501 4428 10140
rect 4462 9501 4468 10140
rect 4580 9840 4586 10477
rect 4620 9840 4626 10477
rect 4738 10477 4784 10489
rect 4738 10450 4744 10477
rect 4778 10450 4784 10477
rect 4896 10477 4942 10489
rect 4720 10380 4730 10450
rect 4800 10380 4810 10450
rect 4738 10210 4744 10380
rect 4778 10210 4784 10380
rect 4720 10140 4730 10210
rect 4800 10140 4810 10210
rect 4560 9770 4570 9840
rect 4640 9770 4650 9840
rect 4580 9600 4586 9770
rect 4620 9600 4626 9770
rect 4560 9530 4570 9600
rect 4640 9530 4650 9600
rect 4422 9489 4468 9501
rect 4580 9501 4586 9530
rect 4620 9501 4626 9530
rect 4580 9489 4626 9501
rect 4738 9501 4744 10140
rect 4778 9501 4784 10140
rect 4896 9840 4902 10477
rect 4936 9840 4942 10477
rect 5054 10477 5100 10489
rect 5054 10450 5060 10477
rect 5094 10450 5100 10477
rect 5030 10380 5040 10450
rect 5110 10380 5120 10450
rect 5054 10210 5060 10380
rect 5094 10210 5100 10380
rect 5030 10140 5040 10210
rect 5110 10140 5120 10210
rect 5170 10150 5250 10530
rect 6570 10289 6701 11310
rect 7098 10289 7104 11403
rect 6570 10277 7104 10289
rect 9000 11403 9535 11415
rect 9000 10289 9132 11403
rect 9529 10289 9535 11403
rect 9000 10277 9535 10289
rect 6570 10150 7010 10277
rect 4880 9770 4890 9840
rect 4960 9770 4970 9840
rect 4896 9600 4902 9770
rect 4936 9600 4942 9770
rect 4880 9530 4890 9600
rect 4960 9530 4970 9600
rect 4738 9489 4784 9501
rect 4896 9501 4902 9530
rect 4936 9501 4942 9530
rect 4896 9489 4942 9501
rect 5054 9501 5060 10140
rect 5094 9501 5100 10140
rect 5054 9489 5100 9501
rect 5170 9955 7010 10150
rect 9000 9955 9440 10277
rect 5170 9943 7104 9955
rect 5170 9860 6701 9943
rect 5170 9450 5250 9860
rect -1410 9442 5250 9450
rect -1410 9408 -1198 9442
rect -1130 9408 -1040 9442
rect -972 9408 -882 9442
rect -814 9408 -724 9442
rect -656 9408 -566 9442
rect -498 9408 -408 9442
rect -340 9408 -250 9442
rect -182 9430 -92 9442
rect -182 9408 -160 9430
rect -24 9408 66 9442
rect 134 9408 224 9442
rect 292 9408 382 9442
rect 450 9408 540 9442
rect 608 9408 698 9442
rect 766 9408 856 9442
rect 924 9408 1014 9442
rect 1082 9408 1172 9442
rect 1240 9408 1330 9442
rect 1398 9408 1488 9442
rect 1556 9408 1646 9442
rect 1714 9408 1804 9442
rect 1872 9408 1962 9442
rect 2030 9408 2120 9442
rect 2188 9408 2278 9442
rect 2346 9408 2436 9442
rect 2504 9408 2594 9442
rect 2662 9408 2752 9442
rect 2820 9408 2910 9442
rect 2978 9408 3068 9442
rect 3136 9408 3226 9442
rect 3294 9408 3384 9442
rect 3452 9408 3542 9442
rect 3610 9408 3700 9442
rect 3768 9408 3858 9442
rect 3926 9430 4016 9442
rect 3980 9408 4016 9430
rect 4084 9408 4174 9442
rect 4242 9408 4332 9442
rect 4400 9408 4490 9442
rect 4558 9408 4648 9442
rect 4716 9408 4806 9442
rect 4874 9408 4964 9442
rect 5032 9408 5250 9442
rect -1410 9400 -160 9408
rect -200 9350 -160 9400
rect -80 9400 3900 9408
rect -80 9350 -40 9400
rect 3860 9350 3900 9400
rect 3980 9400 5250 9408
rect 3980 9350 4020 9400
rect -200 9340 -40 9350
rect 1020 9346 2810 9350
rect 277 9340 3557 9346
rect 3860 9340 4020 9350
rect 277 9306 289 9340
rect 3545 9306 3557 9340
rect 277 9300 3557 9306
rect 1020 9290 2810 9300
rect 1020 9020 1270 9290
rect 1540 9020 2320 9290
rect 2590 9020 2810 9290
rect 1020 9002 2810 9020
rect 1020 8968 1038 9002
rect 2794 8968 2810 9002
rect 1020 8960 2810 8968
rect -2730 8817 -2195 8829
rect 90 8900 3740 8910
rect 90 8866 302 8900
rect 370 8866 460 8900
rect 528 8866 618 8900
rect 686 8866 776 8900
rect 844 8866 934 8900
rect 1002 8866 1092 8900
rect 1160 8866 1250 8900
rect 1318 8866 1408 8900
rect 1476 8866 1566 8900
rect 1634 8866 1724 8900
rect 1792 8866 1882 8900
rect 1950 8866 2040 8900
rect 2108 8866 2198 8900
rect 2266 8866 2356 8900
rect 2424 8866 2514 8900
rect 2582 8866 2672 8900
rect 2740 8866 2830 8900
rect 2898 8866 2988 8900
rect 3056 8866 3146 8900
rect 3214 8866 3304 8900
rect 3372 8866 3462 8900
rect 3530 8866 3740 8900
rect 90 8860 3740 8866
rect -5540 8700 -4730 8817
rect -3924 8722 -3670 8728
rect -4074 8636 -3912 8722
rect -3682 8636 -3482 8722
rect -2730 8700 -2290 8817
rect -4074 8360 -3482 8636
rect -4950 8230 -2500 8360
rect -4950 8220 -2940 8230
rect -4950 8060 -4610 8220
rect -4480 8070 -2940 8220
rect -2810 8070 -2500 8230
rect -4480 8060 -2500 8070
rect -4950 7920 -2500 8060
rect -4060 1290 -3540 7920
rect 90 7780 170 8860
rect 234 8807 280 8819
rect 234 8780 240 8807
rect 274 8780 280 8807
rect 392 8807 438 8819
rect 210 8710 220 8780
rect 290 8710 300 8780
rect 234 8570 240 8710
rect 274 8570 280 8710
rect 210 8500 220 8570
rect 290 8500 300 8570
rect 234 7831 240 8500
rect 274 7831 280 8500
rect 392 8140 398 8807
rect 432 8140 438 8807
rect 550 8807 596 8819
rect 550 8780 556 8807
rect 590 8780 596 8807
rect 708 8807 754 8819
rect 530 8710 540 8780
rect 610 8710 620 8780
rect 550 8570 556 8710
rect 590 8570 596 8710
rect 530 8500 540 8570
rect 610 8500 620 8570
rect 370 8070 380 8140
rect 450 8070 460 8140
rect 392 7930 398 8070
rect 432 7930 438 8070
rect 370 7860 380 7930
rect 450 7860 460 7930
rect 234 7819 280 7831
rect 392 7831 398 7860
rect 432 7831 438 7860
rect 392 7819 438 7831
rect 550 7831 556 8500
rect 590 7831 596 8500
rect 708 8140 714 8807
rect 748 8140 754 8807
rect 866 8807 912 8819
rect 866 8780 872 8807
rect 906 8780 912 8807
rect 1024 8807 1070 8819
rect 840 8710 850 8780
rect 920 8710 930 8780
rect 866 8570 872 8710
rect 906 8570 912 8710
rect 840 8500 850 8570
rect 920 8500 930 8570
rect 690 8070 700 8140
rect 770 8070 780 8140
rect 708 7930 714 8070
rect 748 7930 754 8070
rect 690 7860 700 7930
rect 770 7860 780 7930
rect 550 7819 596 7831
rect 708 7831 714 7860
rect 748 7831 754 7860
rect 708 7819 754 7831
rect 866 7831 872 8500
rect 906 7831 912 8500
rect 1024 8140 1030 8807
rect 1064 8140 1070 8807
rect 1182 8807 1228 8819
rect 1182 8780 1188 8807
rect 1222 8780 1228 8807
rect 1340 8807 1386 8819
rect 1160 8710 1170 8780
rect 1240 8710 1250 8780
rect 1182 8570 1188 8710
rect 1222 8570 1228 8710
rect 1160 8500 1170 8570
rect 1240 8500 1250 8570
rect 1000 8070 1010 8140
rect 1080 8070 1090 8140
rect 1024 7930 1030 8070
rect 1064 7930 1070 8070
rect 1000 7860 1010 7930
rect 1080 7860 1090 7930
rect 866 7819 912 7831
rect 1024 7831 1030 7860
rect 1064 7831 1070 7860
rect 1024 7819 1070 7831
rect 1182 7831 1188 8500
rect 1222 7831 1228 8500
rect 1340 8140 1346 8807
rect 1380 8140 1386 8807
rect 1498 8807 1544 8819
rect 1498 8780 1504 8807
rect 1538 8780 1544 8807
rect 1656 8807 1702 8819
rect 1480 8710 1490 8780
rect 1560 8710 1570 8780
rect 1498 8570 1504 8710
rect 1538 8570 1544 8710
rect 1480 8500 1490 8570
rect 1560 8500 1570 8570
rect 1320 8070 1330 8140
rect 1400 8070 1410 8140
rect 1340 7930 1346 8070
rect 1380 7930 1386 8070
rect 1320 7860 1330 7930
rect 1400 7860 1410 7930
rect 1182 7819 1228 7831
rect 1340 7831 1346 7860
rect 1380 7831 1386 7860
rect 1340 7819 1386 7831
rect 1498 7831 1504 8500
rect 1538 7831 1544 8500
rect 1656 8140 1662 8807
rect 1696 8140 1702 8807
rect 1814 8807 1860 8819
rect 1814 8780 1820 8807
rect 1854 8780 1860 8807
rect 1972 8807 2018 8819
rect 1790 8710 1800 8780
rect 1870 8710 1880 8780
rect 1814 8570 1820 8710
rect 1854 8570 1860 8710
rect 1790 8500 1800 8570
rect 1870 8500 1880 8570
rect 1640 8070 1650 8140
rect 1720 8070 1730 8140
rect 1656 7930 1662 8070
rect 1696 7930 1702 8070
rect 1640 7860 1650 7930
rect 1720 7860 1730 7930
rect 1498 7819 1544 7831
rect 1656 7831 1662 7860
rect 1696 7831 1702 7860
rect 1656 7819 1702 7831
rect 1814 7831 1820 8500
rect 1854 7831 1860 8500
rect 1972 8140 1978 8807
rect 2012 8140 2018 8807
rect 2130 8807 2176 8819
rect 2130 8780 2136 8807
rect 2170 8780 2176 8807
rect 2288 8807 2334 8819
rect 2110 8710 2120 8780
rect 2190 8710 2200 8780
rect 2130 8570 2136 8710
rect 2170 8570 2176 8710
rect 2110 8500 2120 8570
rect 2190 8500 2200 8570
rect 1950 8070 1960 8140
rect 2030 8070 2040 8140
rect 1972 7930 1978 8070
rect 2012 7930 2018 8070
rect 1950 7860 1960 7930
rect 2030 7860 2040 7930
rect 1814 7819 1860 7831
rect 1972 7831 1978 7860
rect 2012 7831 2018 7860
rect 1972 7819 2018 7831
rect 2130 7831 2136 8500
rect 2170 7831 2176 8500
rect 2288 8140 2294 8807
rect 2328 8140 2334 8807
rect 2446 8807 2492 8819
rect 2446 8780 2452 8807
rect 2486 8780 2492 8807
rect 2604 8807 2650 8819
rect 2430 8710 2440 8780
rect 2510 8710 2520 8780
rect 2446 8570 2452 8710
rect 2486 8570 2492 8710
rect 2430 8500 2440 8570
rect 2510 8500 2520 8570
rect 2270 8070 2280 8140
rect 2350 8070 2360 8140
rect 2288 7930 2294 8070
rect 2328 7930 2334 8070
rect 2270 7860 2280 7930
rect 2350 7860 2360 7930
rect 2130 7819 2176 7831
rect 2288 7831 2294 7860
rect 2328 7831 2334 7860
rect 2288 7819 2334 7831
rect 2446 7831 2452 8500
rect 2486 7831 2492 8500
rect 2604 8140 2610 8807
rect 2644 8140 2650 8807
rect 2762 8807 2808 8819
rect 2762 8780 2768 8807
rect 2802 8780 2808 8807
rect 2920 8807 2966 8819
rect 2740 8710 2750 8780
rect 2820 8710 2830 8780
rect 2762 8570 2768 8710
rect 2802 8570 2808 8710
rect 2740 8500 2750 8570
rect 2820 8500 2830 8570
rect 2580 8070 2590 8140
rect 2660 8070 2670 8140
rect 2604 7930 2610 8070
rect 2644 7930 2650 8070
rect 2580 7860 2590 7930
rect 2660 7860 2670 7930
rect 2446 7819 2492 7831
rect 2604 7831 2610 7860
rect 2644 7831 2650 7860
rect 2604 7819 2650 7831
rect 2762 7831 2768 8500
rect 2802 7831 2808 8500
rect 2920 8140 2926 8807
rect 2960 8140 2966 8807
rect 3078 8807 3124 8819
rect 3078 8780 3084 8807
rect 3118 8780 3124 8807
rect 3236 8807 3282 8819
rect 3060 8710 3070 8780
rect 3140 8710 3150 8780
rect 3078 8570 3084 8710
rect 3118 8570 3124 8710
rect 3060 8500 3070 8570
rect 3140 8500 3150 8570
rect 2900 8070 2910 8140
rect 2980 8070 2990 8140
rect 2920 7930 2926 8070
rect 2960 7930 2966 8070
rect 2900 7860 2910 7930
rect 2980 7860 2990 7930
rect 2762 7819 2808 7831
rect 2920 7831 2926 7860
rect 2960 7831 2966 7860
rect 2920 7819 2966 7831
rect 3078 7831 3084 8500
rect 3118 7831 3124 8500
rect 3236 8140 3242 8807
rect 3276 8140 3282 8807
rect 3394 8807 3440 8819
rect 3394 8780 3400 8807
rect 3434 8780 3440 8807
rect 3552 8807 3598 8819
rect 3370 8710 3380 8780
rect 3450 8710 3460 8780
rect 3394 8570 3400 8710
rect 3434 8570 3440 8710
rect 3370 8500 3380 8570
rect 3450 8500 3460 8570
rect 3220 8070 3230 8140
rect 3300 8070 3310 8140
rect 3236 7930 3242 8070
rect 3276 7930 3282 8070
rect 3220 7860 3230 7930
rect 3300 7860 3310 7930
rect 3078 7819 3124 7831
rect 3236 7831 3242 7860
rect 3276 7831 3282 7860
rect 3236 7819 3282 7831
rect 3394 7831 3400 8500
rect 3434 7831 3440 8500
rect 3552 8140 3558 8807
rect 3592 8140 3598 8807
rect 3530 8070 3540 8140
rect 3610 8070 3620 8140
rect 3552 7930 3558 8070
rect 3592 7930 3598 8070
rect 3530 7860 3540 7930
rect 3610 7860 3620 7930
rect 3394 7819 3440 7831
rect 3552 7831 3558 7860
rect 3592 7831 3598 7860
rect 3552 7819 3598 7831
rect 3660 7780 3740 8860
rect 6570 8829 6701 9860
rect 7098 8829 7104 9943
rect 6570 8817 7104 8829
rect 9000 9943 9535 9955
rect 9000 8829 9132 9943
rect 9529 8829 9535 9943
rect 9000 8817 9535 8829
rect 6570 8700 7010 8817
rect 7594 8706 7996 8714
rect 7594 8614 7656 8706
rect 7874 8614 7996 8706
rect 9000 8700 9440 8817
rect 7594 8410 7996 8614
rect 6580 8360 9480 8410
rect 6580 8230 7010 8360
rect 7120 8350 9480 8360
rect 7120 8230 8890 8350
rect 6580 8220 8890 8230
rect 9000 8220 9480 8350
rect 6580 8150 9480 8220
rect 90 7772 3740 7780
rect 90 7738 302 7772
rect 370 7738 460 7772
rect 528 7738 618 7772
rect 686 7738 776 7772
rect 844 7738 934 7772
rect 1002 7738 1092 7772
rect 1160 7738 1250 7772
rect 1318 7738 1408 7772
rect 1476 7738 1566 7772
rect 1634 7738 1724 7772
rect 1792 7738 1882 7772
rect 1950 7738 2040 7772
rect 2108 7738 2198 7772
rect 2266 7738 2356 7772
rect 2424 7738 2514 7772
rect 2582 7738 2672 7772
rect 2740 7738 2830 7772
rect 2898 7738 2988 7772
rect 3056 7738 3146 7772
rect 3214 7738 3304 7772
rect 3372 7738 3462 7772
rect 3530 7738 3740 7772
rect 90 7730 3740 7738
rect 280 7370 550 7730
rect 1030 7676 1040 7680
rect 888 7670 1040 7676
rect 1300 7676 1310 7680
rect 1300 7670 1482 7676
rect 888 7430 900 7670
rect 1470 7430 1482 7670
rect 888 7424 1040 7430
rect 1030 7420 1040 7424
rect 1300 7424 1482 7430
rect 1300 7420 1310 7424
rect 1780 7370 2050 7730
rect 2530 7676 2540 7680
rect 2358 7670 2540 7676
rect 2800 7676 2810 7680
rect 2800 7670 2952 7676
rect 2358 7430 2370 7670
rect 2940 7430 2952 7670
rect 2358 7424 2540 7430
rect 2530 7420 2540 7424
rect 2800 7424 2952 7430
rect 2800 7420 2810 7424
rect 3280 7370 3550 7730
rect 280 7360 3550 7370
rect 280 7326 302 7360
rect 370 7326 460 7360
rect 528 7326 618 7360
rect 686 7326 776 7360
rect 844 7326 934 7360
rect 1002 7326 1092 7360
rect 1160 7326 1250 7360
rect 1318 7326 1408 7360
rect 1476 7326 1566 7360
rect 1634 7326 1724 7360
rect 1792 7326 1882 7360
rect 1950 7326 2040 7360
rect 2108 7326 2198 7360
rect 2266 7326 2356 7360
rect 2424 7326 2514 7360
rect 2582 7326 2672 7360
rect 2740 7326 2830 7360
rect 2898 7326 2988 7360
rect 3056 7326 3146 7360
rect 3214 7326 3304 7360
rect 3372 7326 3462 7360
rect 3530 7326 3550 7360
rect 280 7320 3550 7326
rect 234 7267 280 7279
rect 234 7230 240 7267
rect 274 7230 280 7267
rect 392 7267 438 7279
rect 210 7160 220 7230
rect 290 7160 300 7230
rect 234 7020 240 7160
rect 274 7020 280 7160
rect 210 6950 220 7020
rect 290 6950 300 7020
rect 234 6291 240 6950
rect 274 6291 280 6950
rect 392 6600 398 7267
rect 432 6600 438 7267
rect 550 7267 596 7279
rect 550 7230 556 7267
rect 590 7230 596 7267
rect 700 7267 760 7320
rect 530 7160 540 7230
rect 610 7160 620 7230
rect 550 7020 556 7160
rect 590 7020 596 7160
rect 530 6950 540 7020
rect 610 6950 620 7020
rect 370 6530 380 6600
rect 450 6530 460 6600
rect 392 6390 398 6530
rect 432 6390 438 6530
rect 370 6320 380 6390
rect 450 6320 460 6390
rect 234 6279 280 6291
rect 392 6291 398 6320
rect 432 6291 438 6320
rect 392 6279 438 6291
rect 550 6291 556 6950
rect 590 6291 596 6950
rect 700 6600 714 7267
rect 748 6600 760 7267
rect 866 7267 912 7279
rect 866 7230 872 7267
rect 906 7230 912 7267
rect 1020 7267 1080 7320
rect 840 7160 850 7230
rect 920 7160 930 7230
rect 866 7020 872 7160
rect 906 7020 912 7160
rect 840 6950 850 7020
rect 920 6950 930 7020
rect 690 6530 700 6600
rect 770 6530 780 6600
rect 700 6390 714 6530
rect 748 6390 760 6530
rect 690 6320 700 6390
rect 770 6320 780 6390
rect 550 6279 596 6291
rect 700 6291 714 6320
rect 748 6291 760 6320
rect 700 6240 760 6291
rect 866 6291 872 6950
rect 906 6291 912 6950
rect 1020 6600 1030 7267
rect 1064 6600 1080 7267
rect 1182 7267 1228 7279
rect 1182 7230 1188 7267
rect 1222 7230 1228 7267
rect 1340 7267 1386 7279
rect 1160 7160 1170 7230
rect 1240 7160 1250 7230
rect 1182 7020 1188 7160
rect 1222 7020 1228 7160
rect 1160 6950 1170 7020
rect 1240 6950 1250 7020
rect 1000 6530 1010 6600
rect 1080 6530 1090 6600
rect 1020 6390 1030 6530
rect 1064 6390 1080 6530
rect 1000 6320 1010 6390
rect 1080 6320 1090 6390
rect 866 6279 912 6291
rect 1020 6291 1030 6320
rect 1064 6291 1080 6320
rect 1020 6240 1080 6291
rect 1182 6291 1188 6950
rect 1222 6291 1228 6950
rect 1340 6600 1346 7267
rect 1380 6600 1386 7267
rect 1498 7267 1544 7279
rect 1498 7230 1504 7267
rect 1538 7230 1544 7267
rect 1656 7267 1702 7279
rect 1480 7160 1490 7230
rect 1560 7160 1570 7230
rect 1498 7020 1504 7160
rect 1538 7020 1544 7160
rect 1480 6950 1490 7020
rect 1560 6950 1570 7020
rect 1320 6530 1330 6600
rect 1400 6530 1410 6600
rect 1340 6390 1346 6530
rect 1380 6390 1386 6530
rect 1320 6320 1330 6390
rect 1400 6320 1410 6390
rect 1182 6279 1228 6291
rect 1340 6291 1346 6320
rect 1380 6291 1386 6320
rect 1340 6279 1386 6291
rect 1498 6291 1504 6950
rect 1538 6291 1544 6950
rect 1656 6600 1662 7267
rect 1696 6600 1702 7267
rect 1814 7267 1860 7279
rect 1814 7230 1820 7267
rect 1854 7230 1860 7267
rect 1972 7267 2018 7279
rect 1790 7160 1800 7230
rect 1870 7160 1880 7230
rect 1814 7020 1820 7160
rect 1854 7020 1860 7160
rect 1790 6950 1800 7020
rect 1870 6950 1880 7020
rect 1630 6530 1640 6600
rect 1710 6530 1720 6600
rect 1656 6390 1662 6530
rect 1696 6390 1702 6530
rect 1630 6320 1640 6390
rect 1710 6320 1720 6390
rect 1498 6279 1544 6291
rect 1656 6291 1662 6320
rect 1696 6291 1702 6320
rect 1656 6279 1702 6291
rect 1814 6291 1820 6950
rect 1854 6291 1860 6950
rect 1972 6600 1978 7267
rect 2012 6600 2018 7267
rect 2130 7267 2176 7279
rect 2130 7230 2136 7267
rect 2170 7230 2176 7267
rect 2288 7267 2334 7279
rect 2110 7160 2120 7230
rect 2190 7160 2200 7230
rect 2130 7020 2136 7160
rect 2170 7020 2176 7160
rect 2110 6950 2120 7020
rect 2190 6950 2200 7020
rect 1950 6530 1960 6600
rect 2030 6530 2040 6600
rect 1972 6390 1978 6530
rect 2012 6390 2018 6530
rect 1950 6320 1960 6390
rect 2030 6320 2040 6390
rect 1814 6279 1860 6291
rect 1972 6291 1978 6320
rect 2012 6291 2018 6320
rect 1972 6279 2018 6291
rect 2130 6291 2136 6950
rect 2170 6291 2176 6950
rect 2288 6600 2294 7267
rect 2328 6600 2334 7267
rect 2446 7267 2492 7279
rect 2446 7230 2452 7267
rect 2486 7230 2492 7267
rect 2604 7267 2650 7279
rect 2420 7160 2430 7230
rect 2500 7160 2510 7230
rect 2446 7020 2452 7160
rect 2486 7020 2492 7160
rect 2420 6950 2430 7020
rect 2500 6950 2510 7020
rect 2270 6530 2280 6600
rect 2350 6530 2360 6600
rect 2288 6390 2294 6530
rect 2328 6390 2334 6530
rect 2270 6320 2280 6390
rect 2350 6320 2360 6390
rect 2130 6279 2176 6291
rect 2288 6291 2294 6320
rect 2328 6291 2334 6320
rect 2288 6279 2334 6291
rect 2446 6291 2452 6950
rect 2486 6291 2492 6950
rect 2604 6600 2610 7267
rect 2644 6600 2650 7267
rect 2762 7267 2808 7279
rect 2762 7230 2768 7267
rect 2802 7230 2808 7267
rect 2910 7267 2970 7320
rect 2740 7160 2750 7230
rect 2820 7160 2830 7230
rect 2762 7020 2768 7160
rect 2802 7020 2808 7160
rect 2740 6950 2750 7020
rect 2820 6950 2830 7020
rect 2580 6530 2590 6600
rect 2660 6530 2670 6600
rect 2604 6390 2610 6530
rect 2644 6390 2650 6530
rect 2580 6320 2590 6390
rect 2660 6320 2670 6390
rect 2446 6279 2492 6291
rect 2604 6291 2610 6320
rect 2644 6291 2650 6320
rect 2604 6279 2650 6291
rect 2762 6291 2768 6950
rect 2802 6291 2808 6950
rect 2910 6600 2926 7267
rect 2960 6600 2970 7267
rect 3078 7267 3124 7279
rect 3078 7230 3084 7267
rect 3118 7230 3124 7267
rect 3230 7267 3290 7320
rect 3060 7160 3070 7230
rect 3140 7160 3150 7230
rect 3078 7020 3084 7160
rect 3118 7020 3124 7160
rect 3060 6950 3070 7020
rect 3140 6950 3150 7020
rect 2900 6530 2910 6600
rect 2980 6530 2990 6600
rect 2910 6390 2926 6530
rect 2960 6390 2970 6530
rect 2900 6320 2910 6390
rect 2980 6320 2990 6390
rect 2762 6279 2808 6291
rect 2910 6291 2926 6320
rect 2960 6291 2970 6320
rect 2910 6240 2970 6291
rect 3078 6291 3084 6950
rect 3118 6291 3124 6950
rect 3230 6600 3242 7267
rect 3276 6600 3290 7267
rect 3394 7267 3440 7279
rect 3394 7230 3400 7267
rect 3434 7230 3440 7267
rect 3552 7267 3598 7279
rect 3370 7160 3380 7230
rect 3450 7160 3460 7230
rect 3394 7020 3400 7160
rect 3434 7020 3440 7160
rect 3370 6950 3380 7020
rect 3450 6950 3460 7020
rect 3210 6530 3220 6600
rect 3290 6530 3300 6600
rect 3230 6390 3242 6530
rect 3276 6390 3290 6530
rect 3210 6320 3220 6390
rect 3290 6320 3300 6390
rect 3078 6279 3124 6291
rect 3230 6291 3242 6320
rect 3276 6291 3290 6320
rect 3230 6240 3290 6291
rect 3394 6291 3400 6950
rect 3434 6291 3440 6950
rect 3552 6600 3558 7267
rect 3592 6600 3598 7267
rect 3530 6530 3540 6600
rect 3610 6530 3620 6600
rect 3552 6390 3558 6530
rect 3592 6390 3598 6530
rect 3530 6320 3540 6390
rect 3610 6320 3620 6390
rect 3394 6279 3440 6291
rect 3552 6291 3558 6320
rect 3592 6291 3598 6320
rect 3552 6279 3598 6291
rect 280 6232 3550 6240
rect 280 6198 302 6232
rect 370 6198 460 6232
rect 528 6198 618 6232
rect 686 6198 776 6232
rect 844 6198 934 6232
rect 1002 6198 1092 6232
rect 1160 6198 1250 6232
rect 1318 6198 1408 6232
rect 1476 6198 1566 6232
rect 1634 6198 1724 6232
rect 1792 6198 1882 6232
rect 1950 6198 2040 6232
rect 2108 6198 2198 6232
rect 2266 6198 2356 6232
rect 2424 6198 2514 6232
rect 2582 6198 2672 6232
rect 2740 6198 2830 6232
rect 2898 6198 2988 6232
rect 3056 6198 3146 6232
rect 3214 6198 3304 6232
rect 3372 6198 3462 6232
rect 3530 6198 3550 6232
rect 280 6190 3550 6198
rect 1574 5885 2248 5891
rect 1574 5851 1586 5885
rect 2236 5851 2248 5885
rect 1574 5845 2248 5851
rect 1130 5783 2690 5790
rect 1130 5749 1403 5783
rect 1471 5749 1561 5783
rect 1629 5749 1719 5783
rect 1787 5749 1877 5783
rect 1945 5749 2035 5783
rect 2103 5749 2193 5783
rect 2261 5749 2351 5783
rect 2419 5749 2690 5783
rect 1130 5740 2690 5749
rect 1130 4680 1210 5740
rect 1335 5699 1381 5711
rect 1335 5670 1341 5699
rect 1375 5670 1381 5699
rect 1493 5699 1539 5711
rect 1310 5600 1320 5670
rect 1390 5600 1400 5670
rect 1335 5380 1341 5600
rect 1375 5380 1381 5600
rect 1310 5310 1320 5380
rect 1390 5310 1400 5380
rect 1335 4723 1341 5310
rect 1375 4723 1381 5310
rect 1493 5110 1499 5699
rect 1533 5110 1539 5699
rect 1651 5699 1697 5711
rect 1651 5670 1657 5699
rect 1691 5670 1697 5699
rect 1809 5699 1855 5711
rect 1630 5600 1640 5670
rect 1710 5600 1720 5670
rect 1651 5380 1657 5600
rect 1691 5380 1697 5600
rect 1630 5310 1640 5380
rect 1710 5310 1720 5380
rect 1470 5040 1480 5110
rect 1550 5040 1560 5110
rect 1493 4820 1499 5040
rect 1533 4820 1539 5040
rect 1470 4750 1480 4820
rect 1550 4750 1560 4820
rect 1335 4711 1381 4723
rect 1493 4723 1499 4750
rect 1533 4723 1539 4750
rect 1493 4711 1539 4723
rect 1651 4723 1657 5310
rect 1691 4723 1697 5310
rect 1809 5110 1815 5699
rect 1849 5110 1855 5699
rect 1967 5699 2013 5711
rect 1967 5670 1973 5699
rect 2007 5670 2013 5699
rect 2125 5699 2171 5711
rect 1940 5600 1950 5670
rect 2020 5600 2030 5670
rect 1967 5380 1973 5600
rect 2007 5380 2013 5600
rect 1940 5310 1950 5380
rect 2020 5310 2030 5380
rect 1780 5040 1790 5110
rect 1860 5040 1870 5110
rect 1809 4820 1815 5040
rect 1849 4820 1855 5040
rect 1780 4750 1790 4820
rect 1860 4750 1870 4820
rect 1651 4711 1697 4723
rect 1809 4723 1815 4750
rect 1849 4723 1855 4750
rect 1809 4711 1855 4723
rect 1967 4723 1973 5310
rect 2007 4723 2013 5310
rect 2125 5110 2131 5699
rect 2165 5110 2171 5699
rect 2283 5699 2329 5711
rect 2283 5670 2289 5699
rect 2323 5670 2329 5699
rect 2441 5699 2487 5711
rect 2260 5600 2270 5670
rect 2340 5600 2350 5670
rect 2283 5380 2289 5600
rect 2323 5380 2329 5600
rect 2260 5310 2270 5380
rect 2340 5310 2350 5380
rect 2100 5040 2110 5110
rect 2180 5040 2190 5110
rect 2125 4820 2131 5040
rect 2165 4820 2171 5040
rect 2100 4750 2110 4820
rect 2180 4750 2190 4820
rect 1967 4711 2013 4723
rect 2125 4723 2131 4750
rect 2165 4723 2171 4750
rect 2125 4711 2171 4723
rect 2283 4723 2289 5310
rect 2323 4723 2329 5310
rect 2441 5110 2447 5699
rect 2481 5110 2487 5699
rect 2420 5040 2430 5110
rect 2500 5040 2510 5110
rect 2441 4820 2447 5040
rect 2481 4820 2487 5040
rect 2420 4750 2430 4820
rect 2500 4750 2510 4820
rect 2283 4711 2329 4723
rect 2441 4723 2447 4750
rect 2481 4723 2487 4750
rect 2441 4711 2487 4723
rect 2610 4680 2690 5740
rect 1130 4673 2690 4680
rect 1130 4639 1403 4673
rect 1471 4639 1561 4673
rect 1629 4639 1719 4673
rect 1787 4639 1877 4673
rect 1945 4639 2035 4673
rect 2103 4639 2193 4673
rect 2261 4639 2351 4673
rect 2419 4639 2690 4673
rect 1130 4630 2690 4639
rect 1770 4577 1780 4580
rect 1574 4571 1780 4577
rect 2040 4577 2050 4580
rect 2040 4571 2248 4577
rect 1574 4537 1586 4571
rect 2236 4537 2248 4571
rect 1574 4531 1780 4537
rect 1770 4371 1780 4531
rect 1574 4365 1780 4371
rect 2040 4531 2248 4537
rect 2040 4371 2050 4531
rect 2040 4365 2248 4371
rect 1574 4331 1586 4365
rect 2236 4331 2248 4365
rect 1574 4325 1780 4331
rect 1770 4320 1780 4325
rect 2040 4325 2248 4331
rect 2040 4320 2050 4325
rect 1130 4263 2690 4270
rect 1130 4229 1403 4263
rect 1471 4229 1561 4263
rect 1629 4229 1719 4263
rect 1787 4229 1877 4263
rect 1945 4229 2035 4263
rect 2103 4229 2193 4263
rect 2261 4229 2351 4263
rect 2419 4229 2690 4263
rect 1130 4220 2690 4229
rect 1130 3160 1210 4220
rect 1335 4179 1381 4191
rect 1335 4150 1341 4179
rect 1375 4150 1381 4179
rect 1493 4179 1539 4191
rect 1310 4080 1320 4150
rect 1390 4080 1400 4150
rect 1335 3860 1341 4080
rect 1375 3860 1381 4080
rect 1310 3790 1320 3860
rect 1390 3790 1400 3860
rect 1335 3203 1341 3790
rect 1375 3203 1381 3790
rect 1493 3590 1499 4179
rect 1533 3590 1539 4179
rect 1651 4179 1697 4191
rect 1651 4150 1657 4179
rect 1691 4150 1697 4179
rect 1809 4179 1855 4191
rect 1630 4080 1640 4150
rect 1710 4080 1720 4150
rect 1651 3860 1657 4080
rect 1691 3860 1697 4080
rect 1630 3790 1640 3860
rect 1710 3790 1720 3860
rect 1470 3520 1480 3590
rect 1550 3520 1560 3590
rect 1493 3300 1499 3520
rect 1533 3300 1539 3520
rect 1470 3230 1480 3300
rect 1550 3230 1560 3300
rect 1335 3191 1381 3203
rect 1493 3203 1499 3230
rect 1533 3203 1539 3230
rect 1493 3191 1539 3203
rect 1651 3203 1657 3790
rect 1691 3203 1697 3790
rect 1809 3590 1815 4179
rect 1849 3590 1855 4179
rect 1967 4179 2013 4191
rect 1967 4150 1973 4179
rect 2007 4150 2013 4179
rect 2125 4179 2171 4191
rect 1940 4080 1950 4150
rect 2020 4080 2030 4150
rect 1967 3860 1973 4080
rect 2007 3860 2013 4080
rect 1940 3790 1950 3860
rect 2020 3790 2030 3860
rect 1780 3520 1790 3590
rect 1860 3520 1870 3590
rect 1809 3300 1815 3520
rect 1849 3300 1855 3520
rect 1780 3230 1790 3300
rect 1860 3230 1870 3300
rect 1651 3191 1697 3203
rect 1809 3203 1815 3230
rect 1849 3203 1855 3230
rect 1809 3191 1855 3203
rect 1967 3203 1973 3790
rect 2007 3203 2013 3790
rect 2125 3590 2131 4179
rect 2165 3590 2171 4179
rect 2283 4179 2329 4191
rect 2283 4150 2289 4179
rect 2323 4150 2329 4179
rect 2441 4179 2487 4191
rect 2260 4080 2270 4150
rect 2340 4080 2350 4150
rect 2283 3860 2289 4080
rect 2323 3860 2329 4080
rect 2260 3790 2270 3860
rect 2340 3790 2350 3860
rect 2100 3520 2110 3590
rect 2180 3520 2190 3590
rect 2125 3300 2131 3520
rect 2165 3300 2171 3520
rect 2100 3230 2110 3300
rect 2180 3230 2190 3300
rect 1967 3191 2013 3203
rect 2125 3203 2131 3230
rect 2165 3203 2171 3230
rect 2125 3191 2171 3203
rect 2283 3203 2289 3790
rect 2323 3203 2329 3790
rect 2441 3590 2447 4179
rect 2481 3590 2487 4179
rect 2420 3520 2430 3590
rect 2500 3520 2510 3590
rect 2441 3300 2447 3520
rect 2481 3300 2487 3520
rect 2420 3230 2430 3300
rect 2500 3230 2510 3300
rect 2283 3191 2329 3203
rect 2441 3203 2447 3230
rect 2481 3203 2487 3230
rect 2441 3191 2487 3203
rect 2610 3160 2690 4220
rect 1130 3153 2690 3160
rect 1130 3119 1403 3153
rect 1471 3119 1561 3153
rect 1629 3119 1719 3153
rect 1787 3119 1877 3153
rect 1945 3119 2035 3153
rect 2103 3119 2193 3153
rect 2261 3119 2351 3153
rect 2419 3119 2690 3153
rect 1130 3110 2690 3119
rect 1770 3057 1780 3060
rect 1574 3051 1780 3057
rect 2040 3057 2050 3060
rect 2040 3051 2248 3057
rect 1574 3017 1586 3051
rect 2236 3017 2248 3051
rect 1574 3011 1780 3017
rect 1770 2850 1780 3011
rect 1081 2844 1780 2850
rect 2040 3011 2248 3017
rect 2040 2850 2050 3011
rect 2040 2844 2749 2850
rect 1081 2810 1093 2844
rect 2737 2810 2749 2844
rect 1081 2804 1780 2810
rect 1770 2800 1780 2804
rect 2040 2804 2749 2810
rect 2040 2800 2050 2804
rect -490 2750 -480 2780
rect -500 2700 -480 2750
rect -490 2670 -480 2700
rect -370 2750 -360 2780
rect -240 2750 -230 2780
rect -370 2700 -230 2750
rect -370 2670 -360 2700
rect -240 2670 -230 2700
rect -120 2750 -110 2780
rect 3910 2750 3920 2780
rect -120 2742 3920 2750
rect -120 2708 412 2742
rect 580 2708 670 2742
rect 838 2708 928 2742
rect 1096 2708 1186 2742
rect 1354 2708 1444 2742
rect 1612 2708 1702 2742
rect 1870 2708 1960 2742
rect 2128 2708 2218 2742
rect 2386 2708 2476 2742
rect 2644 2708 2734 2742
rect 2902 2708 2992 2742
rect 3160 2708 3250 2742
rect 3418 2708 3920 2742
rect -120 2700 3920 2708
rect -120 2670 -110 2700
rect 3910 2670 3920 2700
rect 4030 2750 4040 2780
rect 4160 2750 4170 2780
rect 4030 2700 4170 2750
rect 4030 2670 4040 2700
rect 4160 2670 4170 2700
rect 4280 2750 4290 2780
rect 4280 2700 4300 2750
rect 4280 2670 4290 2700
rect 344 2658 390 2670
rect 344 2630 350 2658
rect 384 2630 390 2658
rect 602 2658 648 2670
rect 320 2560 330 2630
rect 400 2560 410 2630
rect 344 2450 350 2560
rect 384 2450 390 2560
rect 320 2380 330 2450
rect 400 2380 410 2450
rect 344 1682 350 2380
rect 384 1682 390 2380
rect 602 1960 608 2658
rect 642 1960 648 2658
rect 860 2658 906 2670
rect 860 2630 866 2658
rect 900 2630 906 2658
rect 1118 2658 1164 2670
rect 840 2560 850 2630
rect 920 2560 930 2630
rect 860 2450 866 2560
rect 900 2450 906 2560
rect 840 2380 850 2450
rect 920 2380 930 2450
rect 580 1890 590 1960
rect 660 1890 670 1960
rect 602 1780 608 1890
rect 642 1780 648 1890
rect 580 1710 590 1780
rect 660 1710 670 1780
rect 344 1670 390 1682
rect 602 1682 608 1710
rect 642 1682 648 1710
rect 602 1670 648 1682
rect 860 1682 866 2380
rect 900 1682 906 2380
rect 1118 1960 1124 2658
rect 1158 1960 1164 2658
rect 1376 2658 1422 2670
rect 1376 2630 1382 2658
rect 1416 2630 1422 2658
rect 1634 2658 1680 2670
rect 1350 2560 1360 2630
rect 1430 2560 1440 2630
rect 1376 2450 1382 2560
rect 1416 2450 1422 2560
rect 1350 2380 1360 2450
rect 1430 2380 1440 2450
rect 1090 1890 1100 1960
rect 1170 1890 1180 1960
rect 1118 1780 1124 1890
rect 1158 1780 1164 1890
rect 1090 1710 1100 1780
rect 1170 1710 1180 1780
rect 860 1670 906 1682
rect 1118 1682 1124 1710
rect 1158 1682 1164 1710
rect 1118 1670 1164 1682
rect 1376 1682 1382 2380
rect 1416 1682 1422 2380
rect 1634 1960 1640 2658
rect 1674 1960 1680 2658
rect 1892 2658 1938 2670
rect 1892 2630 1898 2658
rect 1932 2630 1938 2658
rect 2150 2658 2196 2670
rect 1870 2560 1880 2630
rect 1950 2560 1960 2630
rect 1892 2450 1898 2560
rect 1932 2450 1938 2560
rect 1870 2380 1880 2450
rect 1950 2380 1960 2450
rect 1610 1890 1620 1960
rect 1690 1890 1700 1960
rect 1634 1780 1640 1890
rect 1674 1780 1680 1890
rect 1610 1710 1620 1780
rect 1690 1710 1700 1780
rect 1376 1670 1422 1682
rect 1634 1682 1640 1710
rect 1674 1682 1680 1710
rect 1634 1670 1680 1682
rect 1892 1682 1898 2380
rect 1932 1682 1938 2380
rect 2150 1960 2156 2658
rect 2190 1960 2196 2658
rect 2408 2658 2454 2670
rect 2408 2630 2414 2658
rect 2448 2630 2454 2658
rect 2666 2658 2712 2670
rect 2380 2560 2390 2630
rect 2460 2560 2470 2630
rect 2408 2450 2414 2560
rect 2448 2450 2454 2560
rect 2380 2380 2390 2450
rect 2460 2380 2470 2450
rect 2130 1890 2140 1960
rect 2210 1890 2220 1960
rect 2150 1780 2156 1890
rect 2190 1780 2196 1890
rect 2130 1710 2140 1780
rect 2210 1710 2220 1780
rect 1892 1670 1938 1682
rect 2150 1682 2156 1710
rect 2190 1682 2196 1710
rect 2150 1670 2196 1682
rect 2408 1682 2414 2380
rect 2448 1682 2454 2380
rect 2666 1960 2672 2658
rect 2706 1960 2712 2658
rect 2924 2658 2970 2670
rect 2924 2630 2930 2658
rect 2964 2630 2970 2658
rect 3182 2658 3228 2670
rect 2900 2560 2910 2630
rect 2980 2560 2990 2630
rect 2924 2450 2930 2560
rect 2964 2450 2970 2560
rect 2900 2380 2910 2450
rect 2980 2380 2990 2450
rect 2640 1890 2650 1960
rect 2720 1890 2730 1960
rect 2666 1780 2672 1890
rect 2706 1780 2712 1890
rect 2640 1710 2650 1780
rect 2720 1710 2730 1780
rect 2408 1670 2454 1682
rect 2666 1682 2672 1710
rect 2706 1682 2712 1710
rect 2666 1670 2712 1682
rect 2924 1682 2930 2380
rect 2964 1682 2970 2380
rect 3182 1960 3188 2658
rect 3222 1960 3228 2658
rect 3440 2658 3486 2670
rect 3440 2630 3446 2658
rect 3480 2630 3486 2658
rect 3420 2560 3430 2630
rect 3500 2560 3510 2630
rect 3440 2450 3446 2560
rect 3480 2450 3486 2560
rect 3420 2380 3430 2450
rect 3500 2380 3510 2450
rect 3160 1890 3170 1960
rect 3240 1890 3250 1960
rect 3182 1780 3188 1890
rect 3222 1780 3228 1890
rect 3160 1710 3170 1780
rect 3240 1710 3250 1780
rect 2924 1670 2970 1682
rect 3182 1682 3188 1710
rect 3222 1682 3228 1710
rect 3182 1670 3228 1682
rect 3440 1682 3446 2380
rect 3480 1682 3486 2380
rect 3440 1670 3486 1682
rect -490 1640 -480 1670
rect -500 1590 -480 1640
rect -490 1560 -480 1590
rect -370 1640 -360 1670
rect -240 1640 -230 1670
rect -370 1590 -230 1640
rect -370 1560 -360 1590
rect -240 1560 -230 1590
rect -120 1640 -110 1670
rect 3910 1640 3920 1670
rect -120 1632 3920 1640
rect -120 1598 412 1632
rect 580 1598 670 1632
rect 838 1598 928 1632
rect 1096 1598 1186 1632
rect 1354 1598 1444 1632
rect 1612 1598 1702 1632
rect 1870 1598 1960 1632
rect 2128 1598 2218 1632
rect 2386 1598 2476 1632
rect 2644 1598 2734 1632
rect 2902 1598 2992 1632
rect 3160 1598 3250 1632
rect 3418 1598 3920 1632
rect -120 1590 3920 1598
rect -120 1560 -110 1590
rect 3910 1560 3920 1590
rect 4030 1640 4040 1670
rect 4160 1640 4170 1670
rect 4030 1590 4170 1640
rect 4030 1560 4040 1590
rect 4160 1560 4170 1590
rect 4280 1640 4290 1670
rect 4280 1590 4300 1640
rect 4280 1560 4290 1590
rect 1780 1536 1790 1540
rect 1081 1530 1790 1536
rect 2040 1536 2050 1540
rect 2040 1530 2749 1536
rect 1081 1496 1093 1530
rect 2737 1496 2749 1530
rect 1081 1490 1790 1496
rect 1780 1330 1790 1490
rect 950 1324 1790 1330
rect 2040 1490 2749 1496
rect 2040 1330 2050 1490
rect 2040 1324 2876 1330
rect 950 1290 962 1324
rect 2864 1290 2876 1324
rect -4060 1280 -1570 1290
rect 950 1284 2876 1290
rect 1780 1280 2050 1284
rect -4060 1270 -750 1280
rect -4060 850 -1350 1270
rect -760 850 -750 1270
rect -490 1230 -480 1260
rect -500 1180 -480 1230
rect -490 1150 -480 1180
rect -370 1230 -360 1260
rect -240 1230 -230 1260
rect -370 1180 -230 1230
rect -370 1150 -360 1180
rect -240 1150 -230 1180
rect -120 1230 -110 1260
rect 3910 1230 3920 1260
rect -120 1222 3920 1230
rect -120 1188 152 1222
rect 320 1188 410 1222
rect 578 1188 668 1222
rect 836 1188 926 1222
rect 1094 1188 1184 1222
rect 1352 1188 1442 1222
rect 1610 1188 1700 1222
rect 1868 1188 1958 1222
rect 2126 1188 2216 1222
rect 2384 1188 2474 1222
rect 2642 1188 2732 1222
rect 2900 1188 2990 1222
rect 3158 1188 3248 1222
rect 3416 1188 3506 1222
rect 3674 1188 3920 1222
rect -120 1180 3920 1188
rect -120 1150 -110 1180
rect 3910 1150 3920 1180
rect 4030 1230 4040 1260
rect 4160 1230 4170 1260
rect 4030 1180 4170 1230
rect 4030 1150 4040 1180
rect 4160 1150 4170 1180
rect 4280 1230 4290 1260
rect 4280 1180 4300 1230
rect 7330 1200 8240 8150
rect 4280 1150 4290 1180
rect 84 1138 130 1150
rect 84 1110 90 1138
rect 124 1110 130 1138
rect 342 1138 388 1150
rect 60 1040 70 1110
rect 140 1040 150 1110
rect 84 930 90 1040
rect 124 930 130 1040
rect 60 860 70 930
rect 140 860 150 930
rect -4060 840 -750 850
rect 84 162 90 860
rect 124 162 130 860
rect 342 440 348 1138
rect 382 440 388 1138
rect 600 1138 646 1150
rect 600 1110 606 1138
rect 640 1110 646 1138
rect 858 1138 904 1150
rect 580 1040 590 1110
rect 660 1040 670 1110
rect 600 930 606 1040
rect 640 930 646 1040
rect 580 860 590 930
rect 660 860 670 930
rect 320 370 330 440
rect 400 370 410 440
rect 342 260 348 370
rect 382 260 388 370
rect 320 190 330 260
rect 400 190 410 260
rect 84 150 130 162
rect 342 162 348 190
rect 382 162 388 190
rect 342 150 388 162
rect 600 162 606 860
rect 640 162 646 860
rect 858 440 864 1138
rect 898 440 904 1138
rect 1116 1138 1162 1150
rect 1116 1110 1122 1138
rect 1156 1110 1162 1138
rect 1374 1138 1420 1150
rect 1090 1040 1100 1110
rect 1170 1040 1180 1110
rect 1116 930 1122 1040
rect 1156 930 1162 1040
rect 1090 860 1100 930
rect 1170 860 1180 930
rect 830 370 840 440
rect 910 370 920 440
rect 858 260 864 370
rect 898 260 904 370
rect 830 190 840 260
rect 910 190 920 260
rect 600 150 646 162
rect 858 162 864 190
rect 898 162 904 190
rect 858 150 904 162
rect 1116 162 1122 860
rect 1156 162 1162 860
rect 1374 440 1380 1138
rect 1414 440 1420 1138
rect 1632 1138 1678 1150
rect 1632 1110 1638 1138
rect 1672 1110 1678 1138
rect 1890 1138 1936 1150
rect 1610 1040 1620 1110
rect 1690 1040 1700 1110
rect 1632 930 1638 1040
rect 1672 930 1678 1040
rect 1610 860 1620 930
rect 1690 860 1700 930
rect 1350 370 1360 440
rect 1430 370 1440 440
rect 1374 260 1380 370
rect 1414 260 1420 370
rect 1350 190 1360 260
rect 1430 190 1440 260
rect 1116 150 1162 162
rect 1374 162 1380 190
rect 1414 162 1420 190
rect 1374 150 1420 162
rect 1632 162 1638 860
rect 1672 162 1678 860
rect 1890 440 1896 1138
rect 1930 440 1936 1138
rect 2148 1138 2194 1150
rect 2148 1110 2154 1138
rect 2188 1110 2194 1138
rect 2406 1138 2452 1150
rect 2120 1040 2130 1110
rect 2200 1040 2210 1110
rect 2148 930 2154 1040
rect 2188 930 2194 1040
rect 2120 860 2130 930
rect 2200 860 2210 930
rect 1870 370 1880 440
rect 1950 370 1960 440
rect 1890 260 1896 370
rect 1930 260 1936 370
rect 1870 190 1880 260
rect 1950 190 1960 260
rect 1632 150 1678 162
rect 1890 162 1896 190
rect 1930 162 1936 190
rect 1890 150 1936 162
rect 2148 162 2154 860
rect 2188 162 2194 860
rect 2406 440 2412 1138
rect 2446 440 2452 1138
rect 2664 1138 2710 1150
rect 2664 1110 2670 1138
rect 2704 1110 2710 1138
rect 2922 1138 2968 1150
rect 2640 1040 2650 1110
rect 2720 1040 2730 1110
rect 2664 930 2670 1040
rect 2704 930 2710 1040
rect 2640 860 2650 930
rect 2720 860 2730 930
rect 2380 370 2390 440
rect 2460 370 2470 440
rect 2406 260 2412 370
rect 2446 260 2452 370
rect 2380 190 2390 260
rect 2460 190 2470 260
rect 2148 150 2194 162
rect 2406 162 2412 190
rect 2446 162 2452 190
rect 2406 150 2452 162
rect 2664 162 2670 860
rect 2704 162 2710 860
rect 2922 440 2928 1138
rect 2962 440 2968 1138
rect 3180 1138 3226 1150
rect 3180 1110 3186 1138
rect 3220 1110 3226 1138
rect 3438 1138 3484 1150
rect 3160 1040 3170 1110
rect 3240 1040 3250 1110
rect 3180 930 3186 1040
rect 3220 930 3226 1040
rect 3160 860 3170 930
rect 3240 860 3250 930
rect 2900 370 2910 440
rect 2980 370 2990 440
rect 2922 260 2928 370
rect 2962 260 2968 370
rect 2900 190 2910 260
rect 2980 190 2990 260
rect 2664 150 2710 162
rect 2922 162 2928 190
rect 2962 162 2968 190
rect 2922 150 2968 162
rect 3180 162 3186 860
rect 3220 162 3226 860
rect 3438 440 3444 1138
rect 3478 440 3484 1138
rect 3696 1138 3742 1150
rect 3696 1110 3702 1138
rect 3736 1110 3742 1138
rect 3670 1040 3680 1110
rect 3750 1040 3760 1110
rect 3696 930 3702 1040
rect 3736 930 3742 1040
rect 4600 940 4610 1200
rect 5100 950 8240 1200
rect 5100 940 7510 950
rect 3670 860 3680 930
rect 3750 860 3760 930
rect 3410 370 3420 440
rect 3490 370 3500 440
rect 3438 260 3444 370
rect 3478 260 3484 370
rect 3410 190 3420 260
rect 3490 190 3500 260
rect 3180 150 3226 162
rect 3438 162 3444 190
rect 3478 162 3484 190
rect 3438 150 3484 162
rect 3696 162 3702 860
rect 3736 162 3742 860
rect 3696 150 3742 162
rect -490 120 -480 150
rect -500 70 -480 120
rect -490 40 -480 70
rect -370 120 -360 150
rect -240 120 -230 150
rect -370 70 -230 120
rect -370 40 -360 70
rect -240 40 -230 70
rect -120 120 -110 150
rect 3910 120 3920 150
rect -120 112 3920 120
rect -120 78 152 112
rect 320 78 410 112
rect 578 78 668 112
rect 836 78 926 112
rect 1094 78 1184 112
rect 1352 78 1442 112
rect 1610 78 1700 112
rect 1868 78 1958 112
rect 2126 78 2216 112
rect 2384 78 2474 112
rect 2642 78 2732 112
rect 2900 78 2990 112
rect 3158 78 3248 112
rect 3416 78 3506 112
rect 3674 78 3920 112
rect -120 70 3920 78
rect -120 40 -110 70
rect 3910 40 3920 70
rect 4030 120 4040 150
rect 4160 120 4170 150
rect 4030 70 4170 120
rect 4030 40 4040 70
rect 4160 40 4170 70
rect 4280 120 4290 150
rect 4280 70 4300 120
rect 4280 40 4290 70
rect 950 10 2876 16
rect 950 -24 962 10
rect 2864 -24 2876 10
rect 950 -30 1790 -24
rect 1780 -240 1790 -30
rect 2040 -30 2876 -24
rect 2040 -240 2050 -30
<< via1 >>
rect -5390 11820 -5320 11890
rect -5390 11700 -5320 11770
rect -5390 11580 -5320 11650
rect -5390 11460 -5320 11530
rect 9200 11820 9270 11890
rect 9200 11700 9270 11770
rect 9200 11580 9270 11650
rect 9200 11460 9270 11530
rect 1270 10672 1540 10930
rect 2320 10672 2590 10930
rect 1270 10660 1540 10672
rect 2320 10660 2590 10672
rect -1280 10380 -1260 10450
rect -1260 10380 -1226 10450
rect -1226 10380 -1210 10450
rect -1280 10140 -1260 10210
rect -1260 10140 -1226 10210
rect -1226 10140 -1210 10210
rect -960 10380 -944 10450
rect -944 10380 -910 10450
rect -910 10380 -890 10450
rect -960 10140 -944 10210
rect -944 10140 -910 10210
rect -910 10140 -890 10210
rect -1120 9770 -1102 9840
rect -1102 9770 -1068 9840
rect -1068 9770 -1050 9840
rect -1120 9530 -1102 9600
rect -1102 9530 -1068 9600
rect -1068 9530 -1050 9600
rect -650 10380 -628 10450
rect -628 10380 -594 10450
rect -594 10380 -580 10450
rect -650 10140 -628 10210
rect -628 10140 -594 10210
rect -594 10140 -580 10210
rect -810 9770 -786 9840
rect -786 9770 -752 9840
rect -752 9770 -740 9840
rect -810 9530 -786 9600
rect -786 9530 -752 9600
rect -752 9530 -740 9600
rect -330 10380 -312 10450
rect -312 10380 -278 10450
rect -278 10380 -260 10450
rect -330 10140 -312 10210
rect -312 10140 -278 10210
rect -278 10140 -260 10210
rect -490 9770 -470 9840
rect -470 9770 -436 9840
rect -436 9770 -420 9840
rect -490 9530 -470 9600
rect -470 9530 -436 9600
rect -436 9530 -420 9600
rect -20 10380 4 10450
rect 4 10380 38 10450
rect 38 10380 50 10450
rect -20 10140 4 10210
rect 4 10140 38 10210
rect 38 10140 50 10210
rect -170 9770 -154 9840
rect -154 9770 -120 9840
rect -120 9770 -100 9840
rect -170 9530 -154 9600
rect -154 9530 -120 9600
rect -120 9530 -100 9600
rect 300 10380 320 10450
rect 320 10380 354 10450
rect 354 10380 370 10450
rect 300 10140 320 10210
rect 320 10140 354 10210
rect 354 10140 370 10210
rect 140 9770 162 9840
rect 162 9770 196 9840
rect 196 9770 210 9840
rect 140 9530 162 9600
rect 162 9530 196 9600
rect 196 9530 210 9600
rect 620 10380 636 10450
rect 636 10380 670 10450
rect 670 10380 690 10450
rect 620 10140 636 10210
rect 636 10140 670 10210
rect 670 10140 690 10210
rect 460 9770 478 9840
rect 478 9770 512 9840
rect 512 9770 530 9840
rect 460 9530 478 9600
rect 478 9530 512 9600
rect 512 9530 530 9600
rect 930 10380 952 10450
rect 952 10380 986 10450
rect 986 10380 1000 10450
rect 930 10140 952 10210
rect 952 10140 986 10210
rect 986 10140 1000 10210
rect 770 9770 794 9840
rect 794 9770 828 9840
rect 828 9770 840 9840
rect 770 9530 794 9600
rect 794 9530 828 9600
rect 828 9530 840 9600
rect 1250 10380 1268 10450
rect 1268 10380 1302 10450
rect 1302 10380 1320 10450
rect 1250 10140 1268 10210
rect 1268 10140 1302 10210
rect 1302 10140 1320 10210
rect 1090 9770 1110 9840
rect 1110 9770 1144 9840
rect 1144 9770 1160 9840
rect 1090 9530 1110 9600
rect 1110 9530 1144 9600
rect 1144 9530 1160 9600
rect 1570 10380 1584 10450
rect 1584 10380 1618 10450
rect 1618 10380 1640 10450
rect 1570 10140 1584 10210
rect 1584 10140 1618 10210
rect 1618 10140 1640 10210
rect 1410 9770 1426 9840
rect 1426 9770 1460 9840
rect 1460 9770 1480 9840
rect 1410 9530 1426 9600
rect 1426 9530 1460 9600
rect 1460 9530 1480 9600
rect 1880 10380 1900 10450
rect 1900 10380 1934 10450
rect 1934 10380 1950 10450
rect 1880 10140 1900 10210
rect 1900 10140 1934 10210
rect 1934 10140 1950 10210
rect 1720 9770 1742 9840
rect 1742 9770 1776 9840
rect 1776 9770 1790 9840
rect 1720 9530 1742 9600
rect 1742 9530 1776 9600
rect 1776 9530 1790 9600
rect 2200 10380 2216 10450
rect 2216 10380 2250 10450
rect 2250 10380 2270 10450
rect 2200 10140 2216 10210
rect 2216 10140 2250 10210
rect 2250 10140 2270 10210
rect 2040 9770 2058 9840
rect 2058 9770 2092 9840
rect 2092 9770 2110 9840
rect 2040 9530 2058 9600
rect 2058 9530 2092 9600
rect 2092 9530 2110 9600
rect 2510 10380 2532 10450
rect 2532 10380 2566 10450
rect 2566 10380 2580 10450
rect 2510 10140 2532 10210
rect 2532 10140 2566 10210
rect 2566 10140 2580 10210
rect 2360 9770 2374 9840
rect 2374 9770 2408 9840
rect 2408 9770 2430 9840
rect 2360 9530 2374 9600
rect 2374 9530 2408 9600
rect 2408 9530 2430 9600
rect 2830 10380 2848 10450
rect 2848 10380 2882 10450
rect 2882 10380 2900 10450
rect 2830 10140 2848 10210
rect 2848 10140 2882 10210
rect 2882 10140 2900 10210
rect 2670 9770 2690 9840
rect 2690 9770 2724 9840
rect 2724 9770 2740 9840
rect 2670 9530 2690 9600
rect 2690 9530 2724 9600
rect 2724 9530 2740 9600
rect 3150 10380 3164 10450
rect 3164 10380 3198 10450
rect 3198 10380 3220 10450
rect 3150 10140 3164 10210
rect 3164 10140 3198 10210
rect 3198 10140 3220 10210
rect 2990 9770 3006 9840
rect 3006 9770 3040 9840
rect 3040 9770 3060 9840
rect 2990 9530 3006 9600
rect 3006 9530 3040 9600
rect 3040 9530 3060 9600
rect 3460 10380 3480 10450
rect 3480 10380 3514 10450
rect 3514 10380 3530 10450
rect 3460 10140 3480 10210
rect 3480 10140 3514 10210
rect 3514 10140 3530 10210
rect 3300 9770 3322 9840
rect 3322 9770 3356 9840
rect 3356 9770 3370 9840
rect 3300 9530 3322 9600
rect 3322 9530 3356 9600
rect 3356 9530 3370 9600
rect 3780 10380 3796 10450
rect 3796 10380 3830 10450
rect 3830 10380 3850 10450
rect 3780 10140 3796 10210
rect 3796 10140 3830 10210
rect 3830 10140 3850 10210
rect 3620 9770 3638 9840
rect 3638 9770 3672 9840
rect 3672 9770 3690 9840
rect 3620 9530 3638 9600
rect 3638 9530 3672 9600
rect 3672 9530 3690 9600
rect 4090 10380 4112 10450
rect 4112 10380 4146 10450
rect 4146 10380 4160 10450
rect 4090 10140 4112 10210
rect 4112 10140 4146 10210
rect 4146 10140 4160 10210
rect 3940 9770 3954 9840
rect 3954 9770 3988 9840
rect 3988 9770 4010 9840
rect 3940 9530 3954 9600
rect 3954 9530 3988 9600
rect 3988 9530 4010 9600
rect 4410 10380 4428 10450
rect 4428 10380 4462 10450
rect 4462 10380 4480 10450
rect 4410 10140 4428 10210
rect 4428 10140 4462 10210
rect 4462 10140 4480 10210
rect 4250 9770 4270 9840
rect 4270 9770 4304 9840
rect 4304 9770 4320 9840
rect 4250 9530 4270 9600
rect 4270 9530 4304 9600
rect 4304 9530 4320 9600
rect 4730 10380 4744 10450
rect 4744 10380 4778 10450
rect 4778 10380 4800 10450
rect 4730 10140 4744 10210
rect 4744 10140 4778 10210
rect 4778 10140 4800 10210
rect 4570 9770 4586 9840
rect 4586 9770 4620 9840
rect 4620 9770 4640 9840
rect 4570 9530 4586 9600
rect 4586 9530 4620 9600
rect 4620 9530 4640 9600
rect 5040 10380 5060 10450
rect 5060 10380 5094 10450
rect 5094 10380 5110 10450
rect 5040 10140 5060 10210
rect 5060 10140 5094 10210
rect 5094 10140 5110 10210
rect 4890 9770 4902 9840
rect 4902 9770 4936 9840
rect 4936 9770 4960 9840
rect 4890 9530 4902 9600
rect 4902 9530 4936 9600
rect 4936 9530 4960 9600
rect -160 9408 -92 9430
rect -92 9408 -80 9430
rect 3900 9408 3926 9430
rect 3926 9408 3980 9430
rect -160 9350 -80 9408
rect 3900 9350 3980 9408
rect 1270 9020 1540 9290
rect 2320 9020 2590 9290
rect 220 8710 240 8780
rect 240 8710 274 8780
rect 274 8710 290 8780
rect 220 8500 240 8570
rect 240 8500 274 8570
rect 274 8500 290 8570
rect 540 8710 556 8780
rect 556 8710 590 8780
rect 590 8710 610 8780
rect 540 8500 556 8570
rect 556 8500 590 8570
rect 590 8500 610 8570
rect 380 8070 398 8140
rect 398 8070 432 8140
rect 432 8070 450 8140
rect 380 7860 398 7930
rect 398 7860 432 7930
rect 432 7860 450 7930
rect 850 8710 872 8780
rect 872 8710 906 8780
rect 906 8710 920 8780
rect 850 8500 872 8570
rect 872 8500 906 8570
rect 906 8500 920 8570
rect 700 8070 714 8140
rect 714 8070 748 8140
rect 748 8070 770 8140
rect 700 7860 714 7930
rect 714 7860 748 7930
rect 748 7860 770 7930
rect 1170 8710 1188 8780
rect 1188 8710 1222 8780
rect 1222 8710 1240 8780
rect 1170 8500 1188 8570
rect 1188 8500 1222 8570
rect 1222 8500 1240 8570
rect 1010 8070 1030 8140
rect 1030 8070 1064 8140
rect 1064 8070 1080 8140
rect 1010 7860 1030 7930
rect 1030 7860 1064 7930
rect 1064 7860 1080 7930
rect 1490 8710 1504 8780
rect 1504 8710 1538 8780
rect 1538 8710 1560 8780
rect 1490 8500 1504 8570
rect 1504 8500 1538 8570
rect 1538 8500 1560 8570
rect 1330 8070 1346 8140
rect 1346 8070 1380 8140
rect 1380 8070 1400 8140
rect 1330 7860 1346 7930
rect 1346 7860 1380 7930
rect 1380 7860 1400 7930
rect 1800 8710 1820 8780
rect 1820 8710 1854 8780
rect 1854 8710 1870 8780
rect 1800 8500 1820 8570
rect 1820 8500 1854 8570
rect 1854 8500 1870 8570
rect 1650 8070 1662 8140
rect 1662 8070 1696 8140
rect 1696 8070 1720 8140
rect 1650 7860 1662 7930
rect 1662 7860 1696 7930
rect 1696 7860 1720 7930
rect 2120 8710 2136 8780
rect 2136 8710 2170 8780
rect 2170 8710 2190 8780
rect 2120 8500 2136 8570
rect 2136 8500 2170 8570
rect 2170 8500 2190 8570
rect 1960 8070 1978 8140
rect 1978 8070 2012 8140
rect 2012 8070 2030 8140
rect 1960 7860 1978 7930
rect 1978 7860 2012 7930
rect 2012 7860 2030 7930
rect 2440 8710 2452 8780
rect 2452 8710 2486 8780
rect 2486 8710 2510 8780
rect 2440 8500 2452 8570
rect 2452 8500 2486 8570
rect 2486 8500 2510 8570
rect 2280 8070 2294 8140
rect 2294 8070 2328 8140
rect 2328 8070 2350 8140
rect 2280 7860 2294 7930
rect 2294 7860 2328 7930
rect 2328 7860 2350 7930
rect 2750 8710 2768 8780
rect 2768 8710 2802 8780
rect 2802 8710 2820 8780
rect 2750 8500 2768 8570
rect 2768 8500 2802 8570
rect 2802 8500 2820 8570
rect 2590 8070 2610 8140
rect 2610 8070 2644 8140
rect 2644 8070 2660 8140
rect 2590 7860 2610 7930
rect 2610 7860 2644 7930
rect 2644 7860 2660 7930
rect 3070 8710 3084 8780
rect 3084 8710 3118 8780
rect 3118 8710 3140 8780
rect 3070 8500 3084 8570
rect 3084 8500 3118 8570
rect 3118 8500 3140 8570
rect 2910 8070 2926 8140
rect 2926 8070 2960 8140
rect 2960 8070 2980 8140
rect 2910 7860 2926 7930
rect 2926 7860 2960 7930
rect 2960 7860 2980 7930
rect 3380 8710 3400 8780
rect 3400 8710 3434 8780
rect 3434 8710 3450 8780
rect 3380 8500 3400 8570
rect 3400 8500 3434 8570
rect 3434 8500 3450 8570
rect 3230 8070 3242 8140
rect 3242 8070 3276 8140
rect 3276 8070 3300 8140
rect 3230 7860 3242 7930
rect 3242 7860 3276 7930
rect 3276 7860 3300 7930
rect 3540 8070 3558 8140
rect 3558 8070 3592 8140
rect 3592 8070 3610 8140
rect 3540 7860 3558 7930
rect 3558 7860 3592 7930
rect 3592 7860 3610 7930
rect 1040 7670 1300 7680
rect 1040 7430 1300 7670
rect 1040 7420 1300 7430
rect 2540 7670 2800 7680
rect 2540 7430 2800 7670
rect 2540 7420 2800 7430
rect 220 7160 240 7230
rect 240 7160 274 7230
rect 274 7160 290 7230
rect 220 6950 240 7020
rect 240 6950 274 7020
rect 274 6950 290 7020
rect 540 7160 556 7230
rect 556 7160 590 7230
rect 590 7160 610 7230
rect 540 6950 556 7020
rect 556 6950 590 7020
rect 590 6950 610 7020
rect 380 6530 398 6600
rect 398 6530 432 6600
rect 432 6530 450 6600
rect 380 6320 398 6390
rect 398 6320 432 6390
rect 432 6320 450 6390
rect 850 7160 872 7230
rect 872 7160 906 7230
rect 906 7160 920 7230
rect 850 6950 872 7020
rect 872 6950 906 7020
rect 906 6950 920 7020
rect 700 6530 714 6600
rect 714 6530 748 6600
rect 748 6530 770 6600
rect 700 6320 714 6390
rect 714 6320 748 6390
rect 748 6320 770 6390
rect 1170 7160 1188 7230
rect 1188 7160 1222 7230
rect 1222 7160 1240 7230
rect 1170 6950 1188 7020
rect 1188 6950 1222 7020
rect 1222 6950 1240 7020
rect 1010 6530 1030 6600
rect 1030 6530 1064 6600
rect 1064 6530 1080 6600
rect 1010 6320 1030 6390
rect 1030 6320 1064 6390
rect 1064 6320 1080 6390
rect 1490 7160 1504 7230
rect 1504 7160 1538 7230
rect 1538 7160 1560 7230
rect 1490 6950 1504 7020
rect 1504 6950 1538 7020
rect 1538 6950 1560 7020
rect 1330 6530 1346 6600
rect 1346 6530 1380 6600
rect 1380 6530 1400 6600
rect 1330 6320 1346 6390
rect 1346 6320 1380 6390
rect 1380 6320 1400 6390
rect 1800 7160 1820 7230
rect 1820 7160 1854 7230
rect 1854 7160 1870 7230
rect 1800 6950 1820 7020
rect 1820 6950 1854 7020
rect 1854 6950 1870 7020
rect 1640 6530 1662 6600
rect 1662 6530 1696 6600
rect 1696 6530 1710 6600
rect 1640 6320 1662 6390
rect 1662 6320 1696 6390
rect 1696 6320 1710 6390
rect 2120 7160 2136 7230
rect 2136 7160 2170 7230
rect 2170 7160 2190 7230
rect 2120 6950 2136 7020
rect 2136 6950 2170 7020
rect 2170 6950 2190 7020
rect 1960 6530 1978 6600
rect 1978 6530 2012 6600
rect 2012 6530 2030 6600
rect 1960 6320 1978 6390
rect 1978 6320 2012 6390
rect 2012 6320 2030 6390
rect 2430 7160 2452 7230
rect 2452 7160 2486 7230
rect 2486 7160 2500 7230
rect 2430 6950 2452 7020
rect 2452 6950 2486 7020
rect 2486 6950 2500 7020
rect 2280 6530 2294 6600
rect 2294 6530 2328 6600
rect 2328 6530 2350 6600
rect 2280 6320 2294 6390
rect 2294 6320 2328 6390
rect 2328 6320 2350 6390
rect 2750 7160 2768 7230
rect 2768 7160 2802 7230
rect 2802 7160 2820 7230
rect 2750 6950 2768 7020
rect 2768 6950 2802 7020
rect 2802 6950 2820 7020
rect 2590 6530 2610 6600
rect 2610 6530 2644 6600
rect 2644 6530 2660 6600
rect 2590 6320 2610 6390
rect 2610 6320 2644 6390
rect 2644 6320 2660 6390
rect 3070 7160 3084 7230
rect 3084 7160 3118 7230
rect 3118 7160 3140 7230
rect 3070 6950 3084 7020
rect 3084 6950 3118 7020
rect 3118 6950 3140 7020
rect 2910 6530 2926 6600
rect 2926 6530 2960 6600
rect 2960 6530 2980 6600
rect 2910 6320 2926 6390
rect 2926 6320 2960 6390
rect 2960 6320 2980 6390
rect 3380 7160 3400 7230
rect 3400 7160 3434 7230
rect 3434 7160 3450 7230
rect 3380 6950 3400 7020
rect 3400 6950 3434 7020
rect 3434 6950 3450 7020
rect 3220 6530 3242 6600
rect 3242 6530 3276 6600
rect 3276 6530 3290 6600
rect 3220 6320 3242 6390
rect 3242 6320 3276 6390
rect 3276 6320 3290 6390
rect 3540 6530 3558 6600
rect 3558 6530 3592 6600
rect 3592 6530 3610 6600
rect 3540 6320 3558 6390
rect 3558 6320 3592 6390
rect 3592 6320 3610 6390
rect 1320 5600 1341 5670
rect 1341 5600 1375 5670
rect 1375 5600 1390 5670
rect 1320 5310 1341 5380
rect 1341 5310 1375 5380
rect 1375 5310 1390 5380
rect 1640 5600 1657 5670
rect 1657 5600 1691 5670
rect 1691 5600 1710 5670
rect 1640 5310 1657 5380
rect 1657 5310 1691 5380
rect 1691 5310 1710 5380
rect 1480 5040 1499 5110
rect 1499 5040 1533 5110
rect 1533 5040 1550 5110
rect 1480 4750 1499 4820
rect 1499 4750 1533 4820
rect 1533 4750 1550 4820
rect 1950 5600 1973 5670
rect 1973 5600 2007 5670
rect 2007 5600 2020 5670
rect 1950 5310 1973 5380
rect 1973 5310 2007 5380
rect 2007 5310 2020 5380
rect 1790 5040 1815 5110
rect 1815 5040 1849 5110
rect 1849 5040 1860 5110
rect 1790 4750 1815 4820
rect 1815 4750 1849 4820
rect 1849 4750 1860 4820
rect 2270 5600 2289 5670
rect 2289 5600 2323 5670
rect 2323 5600 2340 5670
rect 2270 5310 2289 5380
rect 2289 5310 2323 5380
rect 2323 5310 2340 5380
rect 2110 5040 2131 5110
rect 2131 5040 2165 5110
rect 2165 5040 2180 5110
rect 2110 4750 2131 4820
rect 2131 4750 2165 4820
rect 2165 4750 2180 4820
rect 2430 5040 2447 5110
rect 2447 5040 2481 5110
rect 2481 5040 2500 5110
rect 2430 4750 2447 4820
rect 2447 4750 2481 4820
rect 2481 4750 2500 4820
rect 1780 4571 2040 4580
rect 1780 4537 2040 4571
rect 1780 4365 2040 4537
rect 1780 4331 2040 4365
rect 1780 4320 2040 4331
rect 1320 4080 1341 4150
rect 1341 4080 1375 4150
rect 1375 4080 1390 4150
rect 1320 3790 1341 3860
rect 1341 3790 1375 3860
rect 1375 3790 1390 3860
rect 1640 4080 1657 4150
rect 1657 4080 1691 4150
rect 1691 4080 1710 4150
rect 1640 3790 1657 3860
rect 1657 3790 1691 3860
rect 1691 3790 1710 3860
rect 1480 3520 1499 3590
rect 1499 3520 1533 3590
rect 1533 3520 1550 3590
rect 1480 3230 1499 3300
rect 1499 3230 1533 3300
rect 1533 3230 1550 3300
rect 1950 4080 1973 4150
rect 1973 4080 2007 4150
rect 2007 4080 2020 4150
rect 1950 3790 1973 3860
rect 1973 3790 2007 3860
rect 2007 3790 2020 3860
rect 1790 3520 1815 3590
rect 1815 3520 1849 3590
rect 1849 3520 1860 3590
rect 1790 3230 1815 3300
rect 1815 3230 1849 3300
rect 1849 3230 1860 3300
rect 2270 4080 2289 4150
rect 2289 4080 2323 4150
rect 2323 4080 2340 4150
rect 2270 3790 2289 3860
rect 2289 3790 2323 3860
rect 2323 3790 2340 3860
rect 2110 3520 2131 3590
rect 2131 3520 2165 3590
rect 2165 3520 2180 3590
rect 2110 3230 2131 3300
rect 2131 3230 2165 3300
rect 2165 3230 2180 3300
rect 2430 3520 2447 3590
rect 2447 3520 2481 3590
rect 2481 3520 2500 3590
rect 2430 3230 2447 3300
rect 2447 3230 2481 3300
rect 2481 3230 2500 3300
rect 1780 3051 2040 3060
rect 1780 3017 2040 3051
rect 1780 2844 2040 3017
rect 1780 2810 2040 2844
rect 1780 2800 2040 2810
rect -480 2670 -370 2780
rect -230 2670 -120 2780
rect 3920 2670 4030 2780
rect 4170 2670 4280 2780
rect 330 2560 350 2630
rect 350 2560 384 2630
rect 384 2560 400 2630
rect 330 2380 350 2450
rect 350 2380 384 2450
rect 384 2380 400 2450
rect 850 2560 866 2630
rect 866 2560 900 2630
rect 900 2560 920 2630
rect 850 2380 866 2450
rect 866 2380 900 2450
rect 900 2380 920 2450
rect 590 1890 608 1960
rect 608 1890 642 1960
rect 642 1890 660 1960
rect 590 1710 608 1780
rect 608 1710 642 1780
rect 642 1710 660 1780
rect 1360 2560 1382 2630
rect 1382 2560 1416 2630
rect 1416 2560 1430 2630
rect 1360 2380 1382 2450
rect 1382 2380 1416 2450
rect 1416 2380 1430 2450
rect 1100 1890 1124 1960
rect 1124 1890 1158 1960
rect 1158 1890 1170 1960
rect 1100 1710 1124 1780
rect 1124 1710 1158 1780
rect 1158 1710 1170 1780
rect 1880 2560 1898 2630
rect 1898 2560 1932 2630
rect 1932 2560 1950 2630
rect 1880 2380 1898 2450
rect 1898 2380 1932 2450
rect 1932 2380 1950 2450
rect 1620 1890 1640 1960
rect 1640 1890 1674 1960
rect 1674 1890 1690 1960
rect 1620 1710 1640 1780
rect 1640 1710 1674 1780
rect 1674 1710 1690 1780
rect 2390 2560 2414 2630
rect 2414 2560 2448 2630
rect 2448 2560 2460 2630
rect 2390 2380 2414 2450
rect 2414 2380 2448 2450
rect 2448 2380 2460 2450
rect 2140 1890 2156 1960
rect 2156 1890 2190 1960
rect 2190 1890 2210 1960
rect 2140 1710 2156 1780
rect 2156 1710 2190 1780
rect 2190 1710 2210 1780
rect 2910 2560 2930 2630
rect 2930 2560 2964 2630
rect 2964 2560 2980 2630
rect 2910 2380 2930 2450
rect 2930 2380 2964 2450
rect 2964 2380 2980 2450
rect 2650 1890 2672 1960
rect 2672 1890 2706 1960
rect 2706 1890 2720 1960
rect 2650 1710 2672 1780
rect 2672 1710 2706 1780
rect 2706 1710 2720 1780
rect 3430 2560 3446 2630
rect 3446 2560 3480 2630
rect 3480 2560 3500 2630
rect 3430 2380 3446 2450
rect 3446 2380 3480 2450
rect 3480 2380 3500 2450
rect 3170 1890 3188 1960
rect 3188 1890 3222 1960
rect 3222 1890 3240 1960
rect 3170 1710 3188 1780
rect 3188 1710 3222 1780
rect 3222 1710 3240 1780
rect -480 1560 -370 1670
rect -230 1560 -120 1670
rect 3920 1560 4030 1670
rect 4170 1560 4280 1670
rect 1790 1530 2040 1540
rect 1790 1496 2040 1530
rect 1790 1324 2040 1496
rect 1790 1290 2040 1324
rect -1350 850 -760 1270
rect -480 1150 -370 1260
rect -230 1150 -120 1260
rect 3920 1150 4030 1260
rect 4170 1150 4280 1260
rect 70 1040 90 1110
rect 90 1040 124 1110
rect 124 1040 140 1110
rect 70 860 90 930
rect 90 860 124 930
rect 124 860 140 930
rect 590 1040 606 1110
rect 606 1040 640 1110
rect 640 1040 660 1110
rect 590 860 606 930
rect 606 860 640 930
rect 640 860 660 930
rect 330 370 348 440
rect 348 370 382 440
rect 382 370 400 440
rect 330 190 348 260
rect 348 190 382 260
rect 382 190 400 260
rect 1100 1040 1122 1110
rect 1122 1040 1156 1110
rect 1156 1040 1170 1110
rect 1100 860 1122 930
rect 1122 860 1156 930
rect 1156 860 1170 930
rect 840 370 864 440
rect 864 370 898 440
rect 898 370 910 440
rect 840 190 864 260
rect 864 190 898 260
rect 898 190 910 260
rect 1620 1040 1638 1110
rect 1638 1040 1672 1110
rect 1672 1040 1690 1110
rect 1620 860 1638 930
rect 1638 860 1672 930
rect 1672 860 1690 930
rect 1360 370 1380 440
rect 1380 370 1414 440
rect 1414 370 1430 440
rect 1360 190 1380 260
rect 1380 190 1414 260
rect 1414 190 1430 260
rect 2130 1040 2154 1110
rect 2154 1040 2188 1110
rect 2188 1040 2200 1110
rect 2130 860 2154 930
rect 2154 860 2188 930
rect 2188 860 2200 930
rect 1880 370 1896 440
rect 1896 370 1930 440
rect 1930 370 1950 440
rect 1880 190 1896 260
rect 1896 190 1930 260
rect 1930 190 1950 260
rect 2650 1040 2670 1110
rect 2670 1040 2704 1110
rect 2704 1040 2720 1110
rect 2650 860 2670 930
rect 2670 860 2704 930
rect 2704 860 2720 930
rect 2390 370 2412 440
rect 2412 370 2446 440
rect 2446 370 2460 440
rect 2390 190 2412 260
rect 2412 190 2446 260
rect 2446 190 2460 260
rect 3170 1040 3186 1110
rect 3186 1040 3220 1110
rect 3220 1040 3240 1110
rect 3170 860 3186 930
rect 3186 860 3220 930
rect 3220 860 3240 930
rect 2910 370 2928 440
rect 2928 370 2962 440
rect 2962 370 2980 440
rect 2910 190 2928 260
rect 2928 190 2962 260
rect 2962 190 2980 260
rect 3680 1040 3702 1110
rect 3702 1040 3736 1110
rect 3736 1040 3750 1110
rect 4610 940 5100 1200
rect 3680 860 3702 930
rect 3702 860 3736 930
rect 3736 860 3750 930
rect 3420 370 3444 440
rect 3444 370 3478 440
rect 3478 370 3490 440
rect 3420 190 3444 260
rect 3444 190 3478 260
rect 3478 190 3490 260
rect -480 40 -370 150
rect -230 40 -120 150
rect 3920 40 4030 150
rect 4170 40 4280 150
rect 1790 -24 2040 10
rect 1790 -240 2040 -24
<< metal2 >>
rect -6510 16440 -6420 16450
rect -6510 16320 -6420 16330
rect -5390 11890 -5320 11900
rect -5390 11810 -5320 11820
rect 9200 11890 9270 11900
rect 9200 11810 9270 11820
rect -5390 11770 -5320 11780
rect -5390 11690 -5320 11700
rect 9200 11770 9270 11780
rect 9200 11690 9270 11700
rect -5390 11650 -5320 11660
rect -5390 11570 -5320 11580
rect 9200 11650 9270 11660
rect 9200 11570 9270 11580
rect -5390 11530 -5320 11540
rect -5390 11450 -5320 11460
rect 9200 11530 9270 11540
rect 9200 11450 9270 11460
rect 1270 10930 1540 10940
rect 1270 10650 1540 10660
rect 2320 10930 2590 10940
rect 2320 10650 2590 10660
rect -1280 10450 -1210 10460
rect -1280 10370 -1210 10380
rect -960 10450 -890 10460
rect -960 10370 -890 10380
rect -650 10450 -580 10460
rect -650 10370 -580 10380
rect -330 10450 -260 10460
rect -330 10370 -260 10380
rect -20 10450 50 10460
rect -20 10370 50 10380
rect 300 10450 370 10460
rect 300 10370 370 10380
rect 620 10450 690 10460
rect 620 10370 690 10380
rect 930 10450 1000 10460
rect 930 10370 1000 10380
rect 1250 10450 1320 10460
rect 1250 10370 1320 10380
rect 1570 10450 1640 10460
rect 1570 10370 1640 10380
rect 1880 10450 1950 10460
rect 1880 10370 1950 10380
rect 2200 10450 2270 10460
rect 2200 10370 2270 10380
rect 2510 10450 2580 10460
rect 2510 10370 2580 10380
rect 2830 10450 2900 10460
rect 2830 10370 2900 10380
rect 3150 10450 3220 10460
rect 3150 10370 3220 10380
rect 3460 10450 3530 10460
rect 3460 10370 3530 10380
rect 3780 10450 3850 10460
rect 3780 10370 3850 10380
rect 4090 10450 4160 10460
rect 4090 10370 4160 10380
rect 4410 10450 4480 10460
rect 4410 10370 4480 10380
rect 4730 10450 4800 10460
rect 4730 10370 4800 10380
rect 5040 10450 5110 10460
rect 5040 10370 5110 10380
rect -1280 10210 -1210 10220
rect -1280 10130 -1210 10140
rect -960 10210 -890 10220
rect -960 10130 -890 10140
rect -650 10210 -580 10220
rect -650 10130 -580 10140
rect -330 10210 -260 10220
rect -330 10130 -260 10140
rect -20 10210 50 10220
rect -20 10130 50 10140
rect 300 10210 370 10220
rect 300 10130 370 10140
rect 620 10210 690 10220
rect 620 10130 690 10140
rect 930 10210 1000 10220
rect 930 10130 1000 10140
rect 1250 10210 1320 10220
rect 1250 10130 1320 10140
rect 1570 10210 1640 10220
rect 1570 10130 1640 10140
rect 1880 10210 1950 10220
rect 1880 10130 1950 10140
rect 2200 10210 2270 10220
rect 2200 10130 2270 10140
rect 2510 10210 2580 10220
rect 2510 10130 2580 10140
rect 2830 10210 2900 10220
rect 2830 10130 2900 10140
rect 3150 10210 3220 10220
rect 3150 10130 3220 10140
rect 3460 10210 3530 10220
rect 3460 10130 3530 10140
rect 3780 10210 3850 10220
rect 3780 10130 3850 10140
rect 4090 10210 4160 10220
rect 4090 10130 4160 10140
rect 4410 10210 4480 10220
rect 4410 10130 4480 10140
rect 4730 10210 4800 10220
rect 4730 10130 4800 10140
rect 5040 10210 5110 10220
rect 5040 10130 5110 10140
rect -1150 9840 -1020 9850
rect -1150 9770 -1120 9840
rect -1050 9770 -1020 9840
rect -1150 9600 -1020 9770
rect -810 9840 -740 9850
rect -810 9760 -740 9770
rect -490 9840 -420 9850
rect -490 9760 -420 9770
rect -170 9840 -100 9850
rect -170 9760 -100 9770
rect 140 9840 210 9850
rect 140 9760 210 9770
rect 460 9840 530 9850
rect 460 9760 530 9770
rect 770 9840 840 9850
rect 770 9760 840 9770
rect 1090 9840 1160 9850
rect 1090 9760 1160 9770
rect 1410 9840 1480 9850
rect 1410 9760 1480 9770
rect 1720 9840 1790 9850
rect 1720 9760 1790 9770
rect 2040 9840 2110 9850
rect 2040 9760 2110 9770
rect 2360 9840 2430 9850
rect 2360 9760 2430 9770
rect 2670 9840 2740 9850
rect 2670 9760 2740 9770
rect 2990 9840 3060 9850
rect 2990 9760 3060 9770
rect 3300 9840 3370 9850
rect 3300 9760 3370 9770
rect 3620 9840 3690 9850
rect 3620 9760 3690 9770
rect 3940 9840 4010 9850
rect 3940 9760 4010 9770
rect 4250 9840 4320 9850
rect 4250 9760 4320 9770
rect 4570 9840 4640 9850
rect 4570 9760 4640 9770
rect 4860 9840 4990 9850
rect 4860 9770 4890 9840
rect 4960 9770 4990 9840
rect -1150 9530 -1120 9600
rect -1050 9530 -1020 9600
rect -1150 9230 -1020 9530
rect -810 9600 -740 9610
rect -810 9520 -740 9530
rect -490 9600 -420 9610
rect -490 9520 -420 9530
rect -170 9600 -100 9610
rect -170 9520 -100 9530
rect 140 9600 210 9610
rect 140 9520 210 9530
rect 460 9600 530 9610
rect 460 9520 530 9530
rect 770 9600 840 9610
rect 770 9520 840 9530
rect 1090 9600 1160 9610
rect 1090 9520 1160 9530
rect 1410 9600 1480 9610
rect 1410 9520 1480 9530
rect 1720 9600 1790 9610
rect 1720 9520 1790 9530
rect 2040 9600 2110 9610
rect 2040 9520 2110 9530
rect 2360 9600 2430 9610
rect 2360 9520 2430 9530
rect 2670 9600 2740 9610
rect 2670 9520 2740 9530
rect 2990 9600 3060 9610
rect 2990 9520 3060 9530
rect 3300 9600 3370 9610
rect 3300 9520 3370 9530
rect 3620 9600 3690 9610
rect 3620 9520 3690 9530
rect 3940 9600 4010 9610
rect 3940 9520 4010 9530
rect 4250 9600 4320 9610
rect 4250 9520 4320 9530
rect 4570 9600 4640 9610
rect 4570 9520 4640 9530
rect 4860 9600 4990 9770
rect 4860 9530 4890 9600
rect 4960 9530 4990 9600
rect -1150 9160 -1120 9230
rect -1050 9160 -1020 9230
rect -1150 2620 -1020 9160
rect -200 9430 -40 9450
rect -200 9350 -160 9430
rect -80 9350 -40 9430
rect -200 8130 -40 9350
rect 3860 9430 4020 9450
rect 3860 9350 3900 9430
rect 3980 9350 4020 9430
rect 1270 9290 1540 9300
rect 1270 9010 1540 9020
rect 2320 9290 2590 9300
rect 2320 9010 2590 9020
rect 220 8780 290 8790
rect 220 8700 290 8710
rect 540 8780 610 8790
rect 540 8700 610 8710
rect 850 8780 920 8790
rect 850 8700 920 8710
rect 1170 8780 1240 8790
rect 1170 8700 1240 8710
rect 1490 8780 1560 8790
rect 1490 8700 1560 8710
rect 1800 8780 1870 8790
rect 1800 8700 1870 8710
rect 2120 8780 2190 8790
rect 2120 8700 2190 8710
rect 2440 8780 2510 8790
rect 2440 8700 2510 8710
rect 2750 8780 2820 8790
rect 2750 8700 2820 8710
rect 3070 8780 3140 8790
rect 3070 8700 3140 8710
rect 3380 8780 3450 8790
rect 3380 8700 3450 8710
rect 220 8570 290 8580
rect 220 8490 290 8500
rect 540 8570 610 8580
rect 540 8490 610 8500
rect 850 8570 920 8580
rect 850 8490 920 8500
rect 1170 8570 1240 8580
rect 1170 8490 1240 8500
rect 1490 8570 1560 8580
rect 1490 8490 1560 8500
rect 1800 8570 1870 8580
rect 1800 8490 1870 8500
rect 2120 8570 2190 8580
rect 2120 8490 2190 8500
rect 2440 8570 2510 8580
rect 2440 8490 2510 8500
rect 2750 8570 2820 8580
rect 2750 8490 2820 8500
rect 3070 8570 3140 8580
rect 3070 8490 3140 8500
rect 3380 8570 3450 8580
rect 3380 8490 3450 8500
rect -200 8050 -160 8130
rect -80 8050 -40 8130
rect 380 8140 450 8150
rect 380 8060 450 8070
rect 700 8140 770 8150
rect 700 8060 770 8070
rect 1010 8140 1080 8150
rect 1010 8060 1080 8070
rect 1330 8140 1400 8150
rect 1330 8060 1400 8070
rect 1650 8140 1720 8150
rect 1650 8060 1720 8070
rect 1960 8140 2030 8150
rect 1960 8060 2030 8070
rect 2280 8140 2350 8150
rect 2280 8060 2350 8070
rect 2590 8140 2660 8150
rect 2590 8060 2660 8070
rect 2910 8140 2980 8150
rect 2910 8060 2980 8070
rect 3230 8140 3300 8150
rect 3230 8060 3300 8070
rect 3540 8140 3610 8150
rect 3540 8060 3610 8070
rect 3860 8130 4020 9350
rect -200 7950 -40 8050
rect -200 7870 -160 7950
rect -80 7870 -40 7950
rect 3860 8050 3900 8130
rect 3980 8050 4020 8130
rect 3860 7950 4020 8050
rect -200 5660 -40 7870
rect 380 7930 450 7940
rect 380 7850 450 7860
rect 700 7930 770 7940
rect 700 7850 770 7860
rect 1010 7930 1080 7940
rect 1010 7850 1080 7860
rect 1330 7930 1400 7940
rect 1330 7850 1400 7860
rect 1650 7930 1720 7940
rect 1650 7850 1720 7860
rect 1960 7930 2030 7940
rect 1960 7850 2030 7860
rect 2280 7930 2350 7940
rect 2280 7850 2350 7860
rect 2590 7930 2660 7940
rect 2590 7850 2660 7860
rect 2910 7930 2980 7940
rect 2910 7850 2980 7860
rect 3230 7930 3300 7940
rect 3230 7850 3300 7860
rect 3540 7930 3610 7940
rect 3540 7850 3610 7860
rect 3860 7870 3900 7950
rect 3980 7870 4020 7950
rect 1040 7680 1300 7690
rect 1040 7410 1300 7420
rect 2540 7680 2800 7690
rect 2540 7410 2800 7420
rect 220 7230 290 7240
rect 220 7150 290 7160
rect 540 7230 610 7240
rect 540 7150 610 7160
rect 850 7230 920 7240
rect 850 7150 920 7160
rect 1170 7230 1240 7240
rect 1170 7150 1240 7160
rect 1490 7230 1560 7240
rect 1490 7150 1560 7160
rect 1800 7230 1870 7240
rect 1800 7150 1870 7160
rect 2120 7230 2190 7240
rect 2120 7150 2190 7160
rect 2430 7230 2500 7240
rect 2430 7150 2500 7160
rect 2750 7230 2820 7240
rect 2750 7150 2820 7160
rect 3070 7230 3140 7240
rect 3070 7150 3140 7160
rect 3380 7230 3450 7240
rect 3380 7150 3450 7160
rect 220 7020 290 7030
rect 220 6940 290 6950
rect 540 7020 610 7030
rect 540 6940 610 6950
rect 850 7020 920 7030
rect 850 6940 920 6950
rect 1170 7020 1240 7030
rect 1170 6940 1240 6950
rect 1490 7020 1560 7030
rect 1490 6940 1560 6950
rect 1800 7020 1870 7030
rect 1800 6940 1870 6950
rect 2120 7020 2190 7030
rect 2120 6940 2190 6950
rect 2430 7020 2500 7030
rect 2430 6940 2500 6950
rect 2750 7020 2820 7030
rect 2750 6940 2820 6950
rect 3070 7020 3140 7030
rect 3070 6940 3140 6950
rect 3380 7020 3450 7030
rect 3380 6940 3450 6950
rect 380 6600 450 6610
rect 380 6520 450 6530
rect 670 6600 800 6610
rect 670 6530 700 6600
rect 770 6530 800 6600
rect 380 6390 450 6400
rect 380 6310 450 6320
rect 670 6390 800 6530
rect 1010 6600 1080 6610
rect 1010 6520 1080 6530
rect 1330 6600 1400 6610
rect 1330 6520 1400 6530
rect 1640 6600 1710 6610
rect 1640 6520 1710 6530
rect 1960 6600 2030 6610
rect 1960 6520 2030 6530
rect 2280 6600 2350 6610
rect 2280 6520 2350 6530
rect 2590 6600 2660 6610
rect 2590 6520 2660 6530
rect 2910 6600 2980 6610
rect 2910 6520 2980 6530
rect 3190 6600 3320 6610
rect 3190 6530 3220 6600
rect 3290 6530 3320 6600
rect 670 6320 700 6390
rect 770 6320 800 6390
rect -200 5540 -180 5660
rect -60 5540 -40 5660
rect -200 5440 -40 5540
rect -200 5320 -180 5440
rect -60 5320 -40 5440
rect -200 5300 -40 5320
rect 40 5100 200 5120
rect 40 4980 60 5100
rect 180 4980 200 5100
rect 40 4880 200 4980
rect 40 4760 60 4880
rect 180 4760 200 4880
rect 40 4140 200 4760
rect 40 4020 60 4140
rect 180 4020 200 4140
rect 40 3920 200 4020
rect 40 3800 60 3920
rect 180 3800 200 3920
rect -1150 2550 -1120 2620
rect -1050 2550 -1020 2620
rect -1150 2460 -1020 2550
rect -1150 2390 -1120 2460
rect -1050 2390 -1020 2460
rect -1150 2370 -1020 2390
rect -500 2780 -100 2900
rect -500 2670 -480 2780
rect -370 2670 -230 2780
rect -120 2670 -100 2780
rect -500 1670 -100 2670
rect -500 1560 -480 1670
rect -370 1560 -230 1670
rect -120 1560 -100 1670
rect -1350 1270 -760 1280
rect -1350 840 -760 850
rect -500 1260 -100 1560
rect -500 1150 -480 1260
rect -370 1150 -230 1260
rect -120 1150 -100 1260
rect -500 150 -100 1150
rect 40 1110 200 3800
rect 670 3570 800 6320
rect 1010 6390 1080 6400
rect 1010 6310 1080 6320
rect 1330 6390 1400 6400
rect 1330 6310 1400 6320
rect 1640 6390 1710 6400
rect 1640 6310 1710 6320
rect 1960 6390 2030 6400
rect 1960 6310 2030 6320
rect 2280 6390 2350 6400
rect 2280 6310 2350 6320
rect 2590 6390 2660 6400
rect 2590 6310 2660 6320
rect 2910 6390 2980 6400
rect 2910 6310 2980 6320
rect 3190 6390 3320 6530
rect 3540 6600 3610 6610
rect 3540 6520 3610 6530
rect 3190 6320 3220 6390
rect 3290 6320 3320 6390
rect 1320 5670 1390 5680
rect 1320 5590 1390 5600
rect 1640 5670 1710 5680
rect 1640 5590 1710 5600
rect 1950 5670 2020 5680
rect 1950 5590 2020 5600
rect 2270 5670 2340 5680
rect 2270 5590 2340 5600
rect 1320 5380 1390 5390
rect 1320 5300 1390 5310
rect 1640 5380 1710 5390
rect 1640 5300 1710 5310
rect 1950 5380 2020 5390
rect 1950 5300 2020 5310
rect 2270 5380 2340 5390
rect 2270 5300 2340 5310
rect 1480 5110 1550 5120
rect 1480 5030 1550 5040
rect 1790 5110 1860 5120
rect 1790 5030 1860 5040
rect 2110 5110 2180 5120
rect 2110 5030 2180 5040
rect 2430 5110 2500 5120
rect 2430 5030 2500 5040
rect 1480 4820 1550 4830
rect 1480 4740 1550 4750
rect 1790 4820 1860 4830
rect 1790 4740 1860 4750
rect 2110 4820 2180 4830
rect 2110 4740 2180 4750
rect 2430 4820 2500 4830
rect 2430 4740 2500 4750
rect 1780 4580 2040 4590
rect 1780 4310 2040 4320
rect 1320 4150 1390 4160
rect 1320 4070 1390 4080
rect 1640 4150 1710 4160
rect 1640 4070 1710 4080
rect 1950 4150 2020 4160
rect 1950 4070 2020 4080
rect 2270 4150 2340 4160
rect 2270 4070 2340 4080
rect 1320 3860 1390 3870
rect 1320 3780 1390 3790
rect 1640 3860 1710 3870
rect 1640 3780 1710 3790
rect 1950 3860 2020 3870
rect 1950 3780 2020 3790
rect 2270 3860 2340 3870
rect 2270 3780 2340 3790
rect 670 3500 700 3570
rect 770 3500 800 3570
rect 1480 3590 1550 3600
rect 1480 3510 1550 3520
rect 1790 3590 1860 3600
rect 1790 3510 1860 3520
rect 2110 3590 2180 3600
rect 2110 3510 2180 3520
rect 2430 3590 2500 3600
rect 2430 3510 2500 3520
rect 3190 3570 3320 6320
rect 3540 6390 3610 6400
rect 3540 6310 3610 6320
rect 3860 5660 4020 7870
rect 3860 5540 3880 5660
rect 4000 5540 4020 5660
rect 3860 5440 4020 5540
rect 3860 5320 3880 5440
rect 4000 5320 4020 5440
rect 3860 5300 4020 5320
rect 4860 9230 4990 9530
rect 4860 9160 4890 9230
rect 4960 9160 4990 9230
rect 670 3320 800 3500
rect 670 3250 700 3320
rect 770 3250 800 3320
rect 3190 3500 3220 3570
rect 3290 3500 3320 3570
rect 3190 3320 3320 3500
rect 670 3220 800 3250
rect 1480 3300 1550 3310
rect 1480 3220 1550 3230
rect 1790 3300 1860 3310
rect 1790 3220 1860 3230
rect 2110 3300 2180 3310
rect 2110 3220 2180 3230
rect 2430 3300 2500 3310
rect 2430 3220 2500 3230
rect 3190 3250 3220 3320
rect 3290 3250 3320 3320
rect 3190 3220 3320 3250
rect 3620 5100 3780 5120
rect 3620 4980 3640 5100
rect 3760 4980 3780 5100
rect 3620 4880 3780 4980
rect 3620 4760 3640 4880
rect 3760 4760 3780 4880
rect 3620 4140 3780 4760
rect 3620 4020 3640 4140
rect 3760 4020 3780 4140
rect 3620 3920 3780 4020
rect 3620 3800 3640 3920
rect 3760 3800 3780 3920
rect 1780 3060 2040 3070
rect 1780 2790 2040 2800
rect 330 2630 400 2640
rect 330 2550 400 2560
rect 850 2630 920 2640
rect 850 2550 920 2560
rect 1360 2630 1430 2640
rect 1360 2550 1430 2560
rect 1880 2630 1950 2640
rect 1880 2550 1950 2560
rect 2390 2630 2460 2640
rect 2390 2550 2460 2560
rect 2910 2630 2980 2640
rect 2910 2550 2980 2560
rect 3430 2630 3500 2640
rect 3430 2550 3500 2560
rect 330 2450 400 2460
rect 330 2370 400 2380
rect 850 2450 920 2460
rect 850 2370 920 2380
rect 1360 2450 1430 2460
rect 1360 2370 1430 2380
rect 1880 2450 1950 2460
rect 1880 2370 1950 2380
rect 2390 2450 2460 2460
rect 2390 2370 2460 2380
rect 2910 2450 2980 2460
rect 2910 2370 2980 2380
rect 3430 2450 3500 2460
rect 3430 2370 3500 2380
rect 590 1960 660 1970
rect 590 1880 660 1890
rect 1100 1960 1170 1970
rect 1100 1880 1170 1890
rect 1620 1960 1690 1970
rect 1620 1880 1690 1890
rect 2140 1960 2210 1970
rect 2140 1880 2210 1890
rect 2650 1960 2720 1970
rect 2650 1880 2720 1890
rect 3170 1960 3240 1970
rect 3170 1880 3240 1890
rect 590 1780 660 1790
rect 590 1700 660 1710
rect 1100 1780 1170 1790
rect 1100 1700 1170 1710
rect 1620 1780 1690 1790
rect 1620 1700 1690 1710
rect 2140 1780 2210 1790
rect 2140 1700 2210 1710
rect 2650 1780 2720 1790
rect 2650 1700 2720 1710
rect 3170 1780 3240 1790
rect 3170 1700 3240 1710
rect 1790 1540 2040 1550
rect 1790 1280 2040 1290
rect 40 1040 70 1110
rect 140 1040 200 1110
rect 40 930 200 1040
rect 590 1110 660 1120
rect 590 1030 660 1040
rect 1100 1110 1170 1120
rect 1100 1030 1170 1040
rect 1620 1110 1690 1120
rect 1620 1030 1690 1040
rect 2130 1110 2200 1120
rect 2130 1030 2200 1040
rect 2650 1110 2720 1120
rect 2650 1030 2720 1040
rect 3170 1110 3240 1120
rect 3170 1030 3240 1040
rect 3620 1110 3780 3800
rect 3620 1040 3680 1110
rect 3750 1040 3780 1110
rect 40 860 70 930
rect 140 860 200 930
rect 40 850 200 860
rect 590 930 660 940
rect 590 850 660 860
rect 1100 930 1170 940
rect 1100 850 1170 860
rect 1620 930 1690 940
rect 1620 850 1690 860
rect 2130 930 2200 940
rect 2130 850 2200 860
rect 2650 930 2720 940
rect 2650 850 2720 860
rect 3170 930 3240 940
rect 3170 850 3240 860
rect 3620 930 3780 1040
rect 3620 860 3680 930
rect 3750 860 3780 930
rect 3620 850 3780 860
rect 3900 2780 4300 2900
rect 3900 2670 3920 2780
rect 4030 2670 4170 2780
rect 4280 2670 4300 2780
rect 3900 1670 4300 2670
rect 4860 2620 4990 9160
rect 4860 2550 4890 2620
rect 4960 2550 4990 2620
rect 4860 2460 4990 2550
rect 4860 2390 4890 2460
rect 4960 2390 4990 2460
rect 4860 2370 4990 2390
rect 3900 1560 3920 1670
rect 4030 1560 4170 1670
rect 4280 1560 4300 1670
rect 3900 1260 4300 1560
rect 3900 1150 3920 1260
rect 4030 1150 4170 1260
rect 4280 1150 4300 1260
rect 330 440 400 450
rect 330 360 400 370
rect 840 440 910 450
rect 840 360 910 370
rect 1360 440 1430 450
rect 1360 360 1430 370
rect 1880 440 1950 450
rect 1880 360 1950 370
rect 2390 440 2460 450
rect 2390 360 2460 370
rect 2910 440 2980 450
rect 2910 360 2980 370
rect 3420 440 3490 450
rect 3420 360 3490 370
rect 330 260 400 270
rect 330 180 400 190
rect 840 260 910 270
rect 840 180 910 190
rect 1360 260 1430 270
rect 1360 180 1430 190
rect 1880 260 1950 270
rect 1880 180 1950 190
rect 2390 260 2460 270
rect 2390 180 2460 190
rect 2910 260 2980 270
rect 2910 180 2980 190
rect 3420 260 3490 270
rect 3420 180 3490 190
rect -500 40 -480 150
rect -370 40 -230 150
rect -120 40 -100 150
rect -500 -100 -100 40
rect 3900 150 4300 1150
rect 4610 1200 5100 1210
rect 4610 930 5100 940
rect 3900 40 3920 150
rect 4030 40 4170 150
rect 4280 40 4300 150
rect 1790 10 2040 20
rect 3900 -100 4300 40
rect 1790 -250 2040 -240
<< via2 >>
rect -6510 16330 -6420 16440
rect -5390 11820 -5320 11890
rect 9200 11820 9270 11890
rect -5390 11700 -5320 11770
rect 9200 11700 9270 11770
rect -5390 11580 -5320 11650
rect 9200 11580 9270 11650
rect -5390 11460 -5320 11530
rect 9200 11460 9270 11530
rect 1270 10660 1540 10930
rect 2320 10660 2590 10930
rect -1280 10380 -1210 10450
rect -960 10380 -890 10450
rect -650 10380 -580 10450
rect -330 10380 -260 10450
rect -20 10380 50 10450
rect 300 10380 370 10450
rect 620 10380 690 10450
rect 930 10380 1000 10450
rect 1250 10380 1320 10450
rect 1570 10380 1640 10450
rect 1880 10380 1950 10450
rect 2200 10380 2270 10450
rect 2510 10380 2580 10450
rect 2830 10380 2900 10450
rect 3150 10380 3220 10450
rect 3460 10380 3530 10450
rect 3780 10380 3850 10450
rect 4090 10380 4160 10450
rect 4410 10380 4480 10450
rect 4730 10380 4800 10450
rect 5040 10380 5110 10450
rect -1280 10140 -1210 10210
rect -960 10140 -890 10210
rect -650 10140 -580 10210
rect -330 10140 -260 10210
rect -20 10140 50 10210
rect 300 10140 370 10210
rect 620 10140 690 10210
rect 930 10140 1000 10210
rect 1250 10140 1320 10210
rect 1570 10140 1640 10210
rect 1880 10140 1950 10210
rect 2200 10140 2270 10210
rect 2510 10140 2580 10210
rect 2830 10140 2900 10210
rect 3150 10140 3220 10210
rect 3460 10140 3530 10210
rect 3780 10140 3850 10210
rect 4090 10140 4160 10210
rect 4410 10140 4480 10210
rect 4730 10140 4800 10210
rect 5040 10140 5110 10210
rect -1120 9770 -1050 9840
rect -810 9770 -740 9840
rect -490 9770 -420 9840
rect -170 9770 -100 9840
rect 140 9770 210 9840
rect 460 9770 530 9840
rect 770 9770 840 9840
rect 1090 9770 1160 9840
rect 1410 9770 1480 9840
rect 1720 9770 1790 9840
rect 2040 9770 2110 9840
rect 2360 9770 2430 9840
rect 2670 9770 2740 9840
rect 2990 9770 3060 9840
rect 3300 9770 3370 9840
rect 3620 9770 3690 9840
rect 3940 9770 4010 9840
rect 4250 9770 4320 9840
rect 4570 9770 4640 9840
rect 4890 9770 4960 9840
rect -1120 9530 -1050 9600
rect -810 9530 -740 9600
rect -490 9530 -420 9600
rect -170 9530 -100 9600
rect 140 9530 210 9600
rect 460 9530 530 9600
rect 770 9530 840 9600
rect 1090 9530 1160 9600
rect 1410 9530 1480 9600
rect 1720 9530 1790 9600
rect 2040 9530 2110 9600
rect 2360 9530 2430 9600
rect 2670 9530 2740 9600
rect 2990 9530 3060 9600
rect 3300 9530 3370 9600
rect 3620 9530 3690 9600
rect 3940 9530 4010 9600
rect 4250 9530 4320 9600
rect 4570 9530 4640 9600
rect 4890 9530 4960 9600
rect -1120 9160 -1050 9230
rect 1270 9020 1540 9290
rect 2320 9020 2590 9290
rect 220 8710 290 8780
rect 540 8710 610 8780
rect 850 8710 920 8780
rect 1170 8710 1240 8780
rect 1490 8710 1560 8780
rect 1800 8710 1870 8780
rect 2120 8710 2190 8780
rect 2440 8710 2510 8780
rect 2750 8710 2820 8780
rect 3070 8710 3140 8780
rect 3380 8710 3450 8780
rect 220 8500 290 8570
rect 540 8500 610 8570
rect 850 8500 920 8570
rect 1170 8500 1240 8570
rect 1490 8500 1560 8570
rect 1800 8500 1870 8570
rect 2120 8500 2190 8570
rect 2440 8500 2510 8570
rect 2750 8500 2820 8570
rect 3070 8500 3140 8570
rect 3380 8500 3450 8570
rect -160 8050 -80 8130
rect 380 8070 450 8140
rect 700 8070 770 8140
rect 1010 8070 1080 8140
rect 1330 8070 1400 8140
rect 1650 8070 1720 8140
rect 1960 8070 2030 8140
rect 2280 8070 2350 8140
rect 2590 8070 2660 8140
rect 2910 8070 2980 8140
rect 3230 8070 3300 8140
rect 3540 8070 3610 8140
rect -160 7870 -80 7950
rect 3900 8050 3980 8130
rect 380 7860 450 7930
rect 700 7860 770 7930
rect 1010 7860 1080 7930
rect 1330 7860 1400 7930
rect 1650 7860 1720 7930
rect 1960 7860 2030 7930
rect 2280 7860 2350 7930
rect 2590 7860 2660 7930
rect 2910 7860 2980 7930
rect 3230 7860 3300 7930
rect 3540 7860 3610 7930
rect 3900 7870 3980 7950
rect 1040 7420 1300 7680
rect 2540 7420 2800 7680
rect 220 7160 290 7230
rect 540 7160 610 7230
rect 850 7160 920 7230
rect 1170 7160 1240 7230
rect 1490 7160 1560 7230
rect 1800 7160 1870 7230
rect 2120 7160 2190 7230
rect 2430 7160 2500 7230
rect 2750 7160 2820 7230
rect 3070 7160 3140 7230
rect 3380 7160 3450 7230
rect 220 6950 290 7020
rect 540 6950 610 7020
rect 850 6950 920 7020
rect 1170 6950 1240 7020
rect 1490 6950 1560 7020
rect 1800 6950 1870 7020
rect 2120 6950 2190 7020
rect 2430 6950 2500 7020
rect 2750 6950 2820 7020
rect 3070 6950 3140 7020
rect 3380 6950 3450 7020
rect 380 6530 450 6600
rect 700 6530 770 6600
rect 380 6320 450 6390
rect 1010 6530 1080 6600
rect 1330 6530 1400 6600
rect 1640 6530 1710 6600
rect 1960 6530 2030 6600
rect 2280 6530 2350 6600
rect 2590 6530 2660 6600
rect 2910 6530 2980 6600
rect 3220 6530 3290 6600
rect 700 6320 770 6390
rect -180 5540 -60 5660
rect -180 5320 -60 5440
rect 60 4980 180 5100
rect 60 4760 180 4880
rect 60 4020 180 4140
rect 60 3800 180 3920
rect -1120 2550 -1050 2620
rect -1120 2390 -1050 2460
rect -1350 850 -760 1270
rect 1010 6320 1080 6390
rect 1330 6320 1400 6390
rect 1640 6320 1710 6390
rect 1960 6320 2030 6390
rect 2280 6320 2350 6390
rect 2590 6320 2660 6390
rect 2910 6320 2980 6390
rect 3540 6530 3610 6600
rect 3220 6320 3290 6390
rect 1320 5600 1390 5670
rect 1640 5600 1710 5670
rect 1950 5600 2020 5670
rect 2270 5600 2340 5670
rect 1320 5310 1390 5380
rect 1640 5310 1710 5380
rect 1950 5310 2020 5380
rect 2270 5310 2340 5380
rect 1480 5040 1550 5110
rect 1790 5040 1860 5110
rect 2110 5040 2180 5110
rect 2430 5040 2500 5110
rect 1480 4750 1550 4820
rect 1790 4750 1860 4820
rect 2110 4750 2180 4820
rect 2430 4750 2500 4820
rect 1780 4320 2040 4580
rect 1320 4080 1390 4150
rect 1640 4080 1710 4150
rect 1950 4080 2020 4150
rect 2270 4080 2340 4150
rect 1320 3790 1390 3860
rect 1640 3790 1710 3860
rect 1950 3790 2020 3860
rect 2270 3790 2340 3860
rect 700 3500 770 3570
rect 1480 3520 1550 3590
rect 1790 3520 1860 3590
rect 2110 3520 2180 3590
rect 2430 3520 2500 3590
rect 3540 6320 3610 6390
rect 3880 5540 4000 5660
rect 3880 5320 4000 5440
rect 4890 9160 4960 9230
rect 700 3250 770 3320
rect 3220 3500 3290 3570
rect 1480 3230 1550 3300
rect 1790 3230 1860 3300
rect 2110 3230 2180 3300
rect 2430 3230 2500 3300
rect 3220 3250 3290 3320
rect 3640 4980 3760 5100
rect 3640 4760 3760 4880
rect 3640 4020 3760 4140
rect 3640 3800 3760 3920
rect 1780 2800 2040 3060
rect 330 2560 400 2630
rect 850 2560 920 2630
rect 1360 2560 1430 2630
rect 1880 2560 1950 2630
rect 2390 2560 2460 2630
rect 2910 2560 2980 2630
rect 3430 2560 3500 2630
rect 330 2380 400 2450
rect 850 2380 920 2450
rect 1360 2380 1430 2450
rect 1880 2380 1950 2450
rect 2390 2380 2460 2450
rect 2910 2380 2980 2450
rect 3430 2380 3500 2450
rect 590 1890 660 1960
rect 1100 1890 1170 1960
rect 1620 1890 1690 1960
rect 2140 1890 2210 1960
rect 2650 1890 2720 1960
rect 3170 1890 3240 1960
rect 590 1710 660 1780
rect 1100 1710 1170 1780
rect 1620 1710 1690 1780
rect 2140 1710 2210 1780
rect 2650 1710 2720 1780
rect 3170 1710 3240 1780
rect 1790 1290 2040 1540
rect 70 1040 140 1110
rect 590 1040 660 1110
rect 1100 1040 1170 1110
rect 1620 1040 1690 1110
rect 2130 1040 2200 1110
rect 2650 1040 2720 1110
rect 3170 1040 3240 1110
rect 3680 1040 3750 1110
rect 70 860 140 930
rect 590 860 660 930
rect 1100 860 1170 930
rect 1620 860 1690 930
rect 2130 860 2200 930
rect 2650 860 2720 930
rect 3170 860 3240 930
rect 3680 860 3750 930
rect 4890 2550 4960 2620
rect 4890 2390 4960 2460
rect 330 370 400 440
rect 840 370 910 440
rect 1360 370 1430 440
rect 1880 370 1950 440
rect 2390 370 2460 440
rect 2910 370 2980 440
rect 3420 370 3490 440
rect 330 190 400 260
rect 840 190 910 260
rect 1360 190 1430 260
rect 1880 190 1950 260
rect 2390 190 2460 260
rect 2910 190 2980 260
rect 3420 190 3490 260
rect 4610 940 5100 1200
rect 1790 -240 2040 10
<< metal3 >>
rect 9890 16490 10100 16550
rect -6530 16440 -6020 16470
rect -6530 16330 -6510 16440
rect -6420 16330 -6250 16440
rect -6160 16330 -6020 16440
rect -6530 12360 -6020 16330
rect -5490 16399 -2090 16419
rect -5490 16335 -5462 16399
rect -2118 16335 -2090 16399
rect -5490 12920 -2090 16335
rect -1690 16399 1710 16419
rect -1690 16335 -1662 16399
rect 1682 16335 1710 16399
rect -1690 12920 1710 16335
rect 2110 16399 5510 16419
rect 2110 16335 2138 16399
rect 5482 16335 5510 16399
rect 2110 12920 5510 16335
rect 5910 16399 9310 16419
rect 5910 16335 5938 16399
rect 9282 16335 9310 16399
rect 5910 12920 9310 16335
rect 9890 16400 9910 16490
rect 9980 16400 10020 16490
rect 10090 16400 10100 16490
rect -6530 12000 -5100 12360
rect 9890 12120 10100 16400
rect -5540 11890 -5100 12000
rect -5540 11820 -5390 11890
rect -5320 11820 -5100 11890
rect -5540 11770 -5100 11820
rect -5540 11700 -5390 11770
rect -5320 11700 -5100 11770
rect -5540 11650 -5100 11700
rect -5540 11580 -5390 11650
rect -5320 11580 -5100 11650
rect -5540 11530 -5100 11580
rect -5540 11460 -5390 11530
rect -5320 11460 -5100 11530
rect -5540 11410 -5100 11460
rect 9080 11930 10100 12120
rect 9080 11890 9450 11930
rect 9080 11820 9200 11890
rect 9270 11820 9450 11890
rect 9080 11770 9450 11820
rect 9080 11700 9200 11770
rect 9270 11700 9450 11770
rect 9080 11650 9450 11700
rect 9080 11580 9200 11650
rect 9270 11580 9450 11650
rect 9080 11530 9450 11580
rect 9080 11460 9200 11530
rect 9270 11460 9450 11530
rect 9080 11410 9450 11460
rect 1260 10930 1550 10935
rect 1260 10660 1270 10930
rect 1540 10660 1550 10930
rect 1260 10655 1550 10660
rect 2310 10930 2600 10935
rect 2310 10660 2320 10930
rect 2590 10660 2600 10930
rect 2310 10655 2600 10660
rect -1280 10455 5110 10460
rect -1290 10450 5120 10455
rect -1290 10380 -1280 10450
rect -1210 10380 -960 10450
rect -890 10430 -650 10450
rect -580 10380 -330 10450
rect -260 10380 -20 10450
rect 50 10380 300 10450
rect 370 10380 620 10450
rect 690 10380 930 10450
rect 1000 10420 1250 10450
rect -1290 10375 -900 10380
rect -1280 10215 -900 10375
rect -1290 10210 -900 10215
rect -650 10210 1000 10380
rect -1290 10140 -1280 10210
rect -1210 10140 -960 10210
rect -890 10140 -650 10180
rect -580 10140 -330 10210
rect -260 10140 -20 10210
rect 50 10140 300 10210
rect 370 10140 620 10210
rect 690 10140 930 10210
rect 1320 10380 1570 10450
rect 1640 10380 1880 10450
rect 1950 10380 2200 10450
rect 2270 10380 2510 10450
rect 2580 10420 2830 10450
rect 1250 10210 2580 10380
rect 1000 10140 1250 10170
rect 1320 10140 1570 10210
rect 1640 10140 1880 10210
rect 1950 10140 2200 10210
rect 2270 10140 2510 10210
rect 2900 10380 3150 10450
rect 3220 10380 3460 10450
rect 3530 10380 3780 10450
rect 3850 10380 4090 10450
rect 4160 10380 4410 10450
rect 4480 10420 4730 10450
rect 2830 10210 4480 10380
rect 2580 10140 2830 10170
rect 2900 10140 3150 10210
rect 3220 10140 3460 10210
rect 3530 10140 3780 10210
rect 3850 10140 4090 10210
rect 4160 10140 4410 10210
rect 4800 10380 5040 10450
rect 5110 10380 5120 10450
rect 4730 10375 5120 10380
rect 4730 10215 5110 10375
rect 4730 10210 5120 10215
rect 4480 10140 4730 10170
rect 4800 10140 5040 10210
rect 5110 10140 5120 10210
rect -1290 10135 5120 10140
rect -1280 10130 5110 10135
rect -1280 9840 5110 9850
rect -1280 9770 -1120 9840
rect -1050 9770 -810 9840
rect -740 9770 -490 9840
rect -420 9770 -170 9840
rect -100 9770 140 9840
rect 210 9770 460 9840
rect 530 9770 770 9840
rect 840 9770 1090 9840
rect 1160 9770 1410 9840
rect 1480 9770 1720 9840
rect 1790 9770 2040 9840
rect 2110 9770 2360 9840
rect 2430 9770 2670 9840
rect 2740 9770 2990 9840
rect 3060 9770 3300 9840
rect 3370 9770 3620 9840
rect 3690 9770 3940 9840
rect 4010 9770 4250 9840
rect 4320 9770 4570 9840
rect 4640 9770 4890 9840
rect 4960 9770 5110 9840
rect -1280 9600 5110 9770
rect -1280 9530 -1120 9600
rect -1050 9530 -810 9600
rect -740 9530 -490 9600
rect -420 9530 -170 9600
rect -100 9530 140 9600
rect 210 9530 460 9600
rect 530 9530 770 9600
rect 840 9530 1090 9600
rect 1160 9530 1410 9600
rect 1480 9530 1720 9600
rect 1790 9530 2040 9600
rect 2110 9530 2360 9600
rect 2430 9530 2670 9600
rect 2740 9530 2990 9600
rect 3060 9530 3300 9600
rect 3370 9530 3620 9600
rect 3690 9530 3940 9600
rect 4010 9530 4250 9600
rect 4320 9530 4570 9600
rect 4640 9530 4890 9600
rect 4960 9530 5110 9600
rect -1280 9520 5110 9530
rect 1260 9290 1550 9295
rect -1790 9230 -1020 9260
rect -1790 9160 -1760 9230
rect -1690 9160 -1120 9230
rect -1050 9160 -1020 9230
rect -1790 9130 -1020 9160
rect 1260 9020 1270 9290
rect 1540 9020 1550 9290
rect 1260 9015 1550 9020
rect 2310 9290 2600 9295
rect 2310 9020 2320 9290
rect 2590 9020 2600 9290
rect 4860 9230 5390 9260
rect 4860 9160 4890 9230
rect 4960 9160 5290 9230
rect 5360 9160 5390 9230
rect 4860 9130 5390 9160
rect 2310 9015 2600 9020
rect 220 8785 3610 8790
rect 210 8780 3610 8785
rect 210 8710 220 8780
rect 290 8710 540 8780
rect 610 8770 850 8780
rect 920 8710 1170 8780
rect 1240 8710 1490 8780
rect 1560 8710 1800 8780
rect 1870 8770 2120 8780
rect 2190 8710 2440 8780
rect 2510 8710 2750 8780
rect 2820 8710 3070 8780
rect 3140 8770 3380 8780
rect 3450 8710 3610 8780
rect 210 8705 600 8710
rect 220 8575 600 8705
rect 210 8570 600 8575
rect 860 8570 1870 8710
rect 2130 8570 3130 8710
rect 3390 8570 3610 8710
rect 210 8500 220 8570
rect 290 8500 540 8570
rect 610 8500 850 8510
rect 920 8500 1170 8570
rect 1240 8500 1490 8570
rect 1560 8500 1800 8570
rect 1870 8500 2120 8510
rect 2190 8500 2440 8570
rect 2510 8500 2750 8570
rect 2820 8500 3070 8570
rect 3140 8500 3380 8510
rect 3450 8500 3610 8570
rect 210 8495 3610 8500
rect 220 8490 3610 8495
rect -200 8140 4020 8150
rect -200 8130 380 8140
rect -200 8050 -160 8130
rect -80 8070 380 8130
rect 450 8070 700 8140
rect 770 8070 1010 8140
rect 1080 8070 1330 8140
rect 1400 8070 1650 8140
rect 1720 8070 1960 8140
rect 2030 8070 2280 8140
rect 2350 8070 2590 8140
rect 2660 8070 2910 8140
rect 2980 8070 3230 8140
rect 3300 8070 3540 8140
rect 3610 8130 4020 8140
rect 3610 8070 3900 8130
rect -80 8050 3900 8070
rect 3980 8050 4020 8130
rect -200 7950 4020 8050
rect -200 7870 -160 7950
rect -80 7930 3900 7950
rect -80 7870 380 7930
rect -200 7860 380 7870
rect 450 7860 700 7930
rect 770 7860 1010 7930
rect 1080 7860 1330 7930
rect 1400 7860 1650 7930
rect 1720 7860 1960 7930
rect 2030 7860 2280 7930
rect 2350 7860 2590 7930
rect 2660 7860 2910 7930
rect 2980 7860 3230 7930
rect 3300 7860 3540 7930
rect 3610 7870 3900 7930
rect 3980 7870 4020 7950
rect 3610 7860 4020 7870
rect -200 7850 4020 7860
rect 1030 7680 1310 7685
rect 1030 7420 1040 7680
rect 1300 7420 1310 7680
rect 1030 7415 1310 7420
rect 2530 7680 2810 7685
rect 2530 7420 2540 7680
rect 2800 7420 2810 7680
rect 2530 7415 2810 7420
rect 220 7235 3610 7240
rect 210 7230 3610 7235
rect 210 7160 220 7230
rect 290 7160 540 7230
rect 610 7220 850 7230
rect 920 7160 1170 7230
rect 1240 7160 1490 7230
rect 1560 7160 1800 7230
rect 1870 7220 2120 7230
rect 2190 7160 2430 7230
rect 2500 7160 2750 7230
rect 2820 7160 3070 7230
rect 3140 7220 3380 7230
rect 3450 7160 3610 7230
rect 210 7155 600 7160
rect 220 7025 600 7155
rect 210 7020 600 7025
rect 860 7020 1870 7160
rect 2130 7020 3130 7160
rect 3390 7020 3610 7160
rect 210 6950 220 7020
rect 290 6950 540 7020
rect 610 6950 850 6960
rect 920 6950 1170 7020
rect 1240 6950 1490 7020
rect 1560 6950 1800 7020
rect 1870 6950 2120 6960
rect 2190 6950 2430 7020
rect 2500 6950 2750 7020
rect 2820 6950 3070 7020
rect 3140 6950 3380 6960
rect 3450 6950 3610 7020
rect 210 6945 3610 6950
rect 220 6940 3610 6945
rect 220 6605 3610 6610
rect 220 6600 3620 6605
rect 220 6530 380 6600
rect 450 6530 700 6600
rect 770 6530 1010 6600
rect 1080 6530 1330 6600
rect 1400 6530 1640 6600
rect 1710 6530 1960 6600
rect 2030 6530 2280 6600
rect 2350 6530 2590 6600
rect 2660 6530 2910 6600
rect 2980 6530 3220 6600
rect 3290 6530 3540 6600
rect 3610 6530 3620 6600
rect 220 6525 3620 6530
rect 220 6395 3610 6525
rect 220 6390 3620 6395
rect 220 6320 380 6390
rect 450 6320 700 6390
rect 770 6320 1010 6390
rect 1080 6320 1330 6390
rect 1400 6320 1640 6390
rect 1710 6320 1960 6390
rect 2030 6320 2280 6390
rect 2350 6320 2590 6390
rect 2660 6320 2910 6390
rect 2980 6320 3220 6390
rect 3290 6320 3540 6390
rect 3610 6320 3620 6390
rect 220 6315 3620 6320
rect 220 6310 3610 6315
rect -200 5670 4020 5680
rect -200 5660 1320 5670
rect -200 5540 -180 5660
rect -60 5600 1320 5660
rect 1390 5600 1640 5670
rect 1710 5600 1950 5670
rect 2020 5600 2270 5670
rect 2340 5660 4020 5670
rect 2340 5600 3880 5660
rect -60 5540 3880 5600
rect 4000 5540 4020 5660
rect -200 5440 4020 5540
rect -200 5320 -180 5440
rect -60 5380 3880 5440
rect -60 5320 1320 5380
rect -200 5310 1320 5320
rect 1390 5310 1640 5380
rect 1710 5310 1950 5380
rect 2020 5310 2270 5380
rect 2340 5320 3880 5380
rect 4000 5320 4020 5440
rect 2340 5310 4020 5320
rect -200 5300 4020 5310
rect 40 5110 3780 5120
rect 40 5100 1480 5110
rect 40 4980 60 5100
rect 180 5040 1480 5100
rect 1550 5040 1790 5110
rect 1860 5040 2110 5110
rect 2180 5040 2430 5110
rect 2500 5100 3780 5110
rect 2500 5040 3640 5100
rect 180 4980 3640 5040
rect 3760 4980 3780 5100
rect 40 4880 3780 4980
rect 40 4760 60 4880
rect 180 4820 3640 4880
rect 180 4760 1480 4820
rect 40 4750 1480 4760
rect 1550 4750 1790 4820
rect 1860 4750 2110 4820
rect 2180 4750 2430 4820
rect 2500 4760 3640 4820
rect 3760 4760 3780 4880
rect 2500 4750 3780 4760
rect 40 4740 3780 4750
rect 1770 4580 2050 4585
rect 1770 4320 1780 4580
rect 2040 4320 2050 4580
rect 1770 4315 2050 4320
rect 40 4150 3780 4160
rect 40 4140 1320 4150
rect 40 4020 60 4140
rect 180 4080 1320 4140
rect 1390 4080 1640 4150
rect 1710 4080 1950 4150
rect 2020 4080 2270 4150
rect 2340 4140 3780 4150
rect 2340 4080 3640 4140
rect 180 4020 3640 4080
rect 3760 4020 3780 4140
rect 40 3920 3780 4020
rect 40 3800 60 3920
rect 180 3860 3640 3920
rect 180 3800 1320 3860
rect 40 3790 1320 3800
rect 1390 3790 1640 3860
rect 1710 3790 1950 3860
rect 2020 3790 2270 3860
rect 2340 3800 3640 3860
rect 3760 3800 3780 3920
rect 2340 3790 3780 3800
rect 40 3780 3780 3790
rect 670 3590 3320 3600
rect 670 3570 1480 3590
rect 670 3500 700 3570
rect 770 3520 1480 3570
rect 1550 3520 1790 3590
rect 1860 3520 2110 3590
rect 2180 3520 2430 3590
rect 2500 3570 3320 3590
rect 2500 3520 3220 3570
rect 770 3500 3220 3520
rect 3290 3500 3320 3570
rect 670 3320 3320 3500
rect 670 3250 700 3320
rect 770 3300 3220 3320
rect 770 3250 1480 3300
rect 670 3230 1480 3250
rect 1550 3230 1790 3300
rect 1860 3230 2110 3300
rect 2180 3230 2430 3300
rect 2500 3250 3220 3300
rect 3290 3250 3320 3320
rect 2500 3230 3320 3250
rect 670 3220 3320 3230
rect 1770 3060 2050 3065
rect 1770 2800 1780 3060
rect 2040 2800 2050 3060
rect 1770 2795 2050 2800
rect -1150 2630 4990 2640
rect -1150 2620 330 2630
rect -1150 2550 -1120 2620
rect -1050 2560 330 2620
rect 400 2560 850 2630
rect 920 2560 1360 2630
rect 1430 2560 1880 2630
rect 1950 2560 2390 2630
rect 2460 2560 2910 2630
rect 2980 2560 3430 2630
rect 3500 2620 4990 2630
rect 3500 2560 4890 2620
rect -1050 2550 4890 2560
rect 4960 2550 4990 2620
rect -1150 2460 4990 2550
rect -1150 2390 -1120 2460
rect -1050 2450 4890 2460
rect -1050 2390 330 2450
rect -1150 2380 330 2390
rect 400 2380 850 2450
rect 920 2380 1360 2450
rect 1430 2380 1880 2450
rect 1950 2380 2390 2450
rect 2460 2380 2910 2450
rect 2980 2380 3430 2450
rect 3500 2390 4890 2450
rect 4960 2390 4990 2460
rect 3500 2380 4990 2390
rect -1150 2370 4990 2380
rect 330 1960 3500 1970
rect 330 1890 590 1960
rect 660 1890 760 1960
rect 330 1780 760 1890
rect 330 1710 590 1780
rect 660 1710 760 1780
rect 1010 1890 1100 1960
rect 1170 1890 1620 1960
rect 1690 1890 2140 1960
rect 2210 1890 2650 1960
rect 2720 1890 2820 1960
rect 1010 1780 2820 1890
rect 1010 1710 1100 1780
rect 1170 1710 1620 1780
rect 1690 1710 2140 1780
rect 2210 1710 2650 1780
rect 2720 1710 2820 1780
rect 3070 1890 3170 1960
rect 3240 1890 3500 1960
rect 3070 1780 3500 1890
rect 3070 1710 3170 1780
rect 3240 1710 3500 1780
rect 330 1700 3500 1710
rect 1780 1540 2050 1545
rect 1780 1290 1790 1540
rect 2040 1290 2050 1540
rect 1780 1285 2050 1290
rect -1360 1270 -750 1275
rect -1360 850 -1350 1270
rect -760 850 -750 1270
rect 4600 1200 5110 1205
rect 70 1115 3750 1120
rect 60 1110 3760 1115
rect 60 1040 70 1110
rect 140 1040 590 1110
rect 660 1040 1100 1110
rect 1170 1040 1620 1110
rect 1690 1040 2130 1110
rect 2200 1040 2650 1110
rect 2720 1040 3170 1110
rect 3240 1040 3680 1110
rect 3750 1040 3760 1110
rect 60 1035 3760 1040
rect 70 935 3750 1035
rect 4600 940 4610 1200
rect 5100 940 5110 1200
rect 4600 935 5110 940
rect 60 930 3760 935
rect 60 860 70 930
rect 140 860 590 930
rect 660 860 1100 930
rect 1170 860 1620 930
rect 1690 860 2130 930
rect 2200 860 2650 930
rect 2720 860 3170 930
rect 3240 860 3680 930
rect 3750 860 3760 930
rect 60 855 3760 860
rect 70 850 3750 855
rect -1360 845 -750 850
rect 70 440 3750 450
rect 70 370 330 440
rect 400 370 500 440
rect 70 260 500 370
rect 70 190 330 260
rect 400 190 500 260
rect 750 370 840 440
rect 910 370 1360 440
rect 1430 370 1880 440
rect 1950 370 2390 440
rect 2460 370 2910 440
rect 2980 370 3080 440
rect 750 260 3080 370
rect 750 190 840 260
rect 910 190 1360 260
rect 1430 190 1880 260
rect 1950 190 2390 260
rect 2460 190 2910 260
rect 2980 190 3080 260
rect 3330 370 3420 440
rect 3490 370 3750 440
rect 3330 260 3750 370
rect 3330 190 3420 260
rect 3490 190 3750 260
rect 70 180 3750 190
rect 1780 10 2050 15
rect 1780 -240 1790 10
rect 2040 -240 2050 10
rect 1780 -245 2050 -240
<< via3 >>
rect -6510 16330 -6420 16440
rect -6250 16330 -6160 16440
rect -5462 16335 -2118 16399
rect -1662 16335 1682 16399
rect 2138 16335 5482 16399
rect 5938 16335 9282 16399
rect 9910 16400 9980 16490
rect 10020 16400 10090 16490
rect 1270 10660 1540 10930
rect 2320 10660 2590 10930
rect -900 10380 -890 10430
rect -890 10380 -650 10430
rect -900 10210 -650 10380
rect -900 10180 -890 10210
rect -890 10180 -650 10210
rect 1000 10170 1250 10420
rect 2580 10170 2830 10420
rect 4480 10170 4730 10420
rect -1760 9160 -1690 9230
rect 1270 9020 1540 9290
rect 2320 9020 2590 9290
rect 5290 9160 5360 9230
rect 600 8710 610 8770
rect 610 8710 850 8770
rect 850 8710 860 8770
rect 1870 8710 2120 8770
rect 2120 8710 2130 8770
rect 3130 8710 3140 8770
rect 3140 8710 3380 8770
rect 3380 8710 3390 8770
rect 600 8570 860 8710
rect 1870 8570 2130 8710
rect 3130 8570 3390 8710
rect 600 8510 610 8570
rect 610 8510 850 8570
rect 850 8510 860 8570
rect 1870 8510 2120 8570
rect 2120 8510 2130 8570
rect 3130 8510 3140 8570
rect 3140 8510 3380 8570
rect 3380 8510 3390 8570
rect 1040 7420 1300 7680
rect 2540 7420 2800 7680
rect 600 7160 610 7220
rect 610 7160 850 7220
rect 850 7160 860 7220
rect 1870 7160 2120 7220
rect 2120 7160 2130 7220
rect 3130 7160 3140 7220
rect 3140 7160 3380 7220
rect 3380 7160 3390 7220
rect 600 7020 860 7160
rect 1870 7020 2130 7160
rect 3130 7020 3390 7160
rect 600 6960 610 7020
rect 610 6960 850 7020
rect 850 6960 860 7020
rect 1870 6960 2120 7020
rect 2120 6960 2130 7020
rect 3130 6960 3140 7020
rect 3140 6960 3380 7020
rect 3380 6960 3390 7020
rect 1780 4320 2040 4580
rect 1780 2800 2040 3060
rect 760 1710 1010 1960
rect 2820 1710 3070 1960
rect 1790 1290 2040 1540
rect -1350 850 -760 1270
rect 4610 940 5100 1200
rect 500 190 750 440
rect 3080 190 3330 440
rect 1790 -240 2040 10
<< mimcap >>
rect -5390 16180 -2190 16220
rect -5390 13060 -5350 16180
rect -2230 13060 -2190 16180
rect -5390 13020 -2190 13060
rect -1590 16180 1610 16220
rect -1590 13060 -1550 16180
rect 1570 13060 1610 16180
rect -1590 13020 1610 13060
rect 2210 16180 5410 16220
rect 2210 13060 2250 16180
rect 5370 13060 5410 16180
rect 2210 13020 5410 13060
rect 6010 16180 9210 16220
rect 6010 13060 6050 16180
rect 9170 13060 9210 16180
rect 6010 13020 9210 13060
<< mimcapcontact >>
rect -5350 13060 -2230 16180
rect -1550 13060 1570 16180
rect 2250 13060 5370 16180
rect 6050 13060 9170 16180
<< metal4 >>
rect -6530 16490 10100 16550
rect -6530 16440 9910 16490
rect -6530 16330 -6510 16440
rect -6420 16330 -6250 16440
rect -6160 16400 9910 16440
rect 9980 16400 10020 16490
rect 10090 16400 10100 16490
rect -6160 16399 10100 16400
rect -6160 16335 -5462 16399
rect -2118 16335 -1662 16399
rect 1682 16335 2138 16399
rect 5482 16335 5938 16399
rect 9282 16335 10100 16399
rect -6160 16330 10100 16335
rect -6530 16310 10100 16330
rect -5351 16180 -2229 16181
rect -5351 13060 -5350 16180
rect -2230 14840 -2229 16180
rect -1551 16180 1571 16181
rect -1551 14840 -1550 16180
rect -2230 14480 -1550 14840
rect -2230 13060 -2229 14480
rect -5351 13059 -2229 13060
rect -1970 11350 -1820 14480
rect -1551 13060 -1550 14480
rect 1570 14840 1571 16180
rect 2249 16180 5371 16181
rect 2249 14840 2250 16180
rect 1570 14480 2250 14840
rect 1570 13060 1571 14480
rect -1551 13059 1571 13060
rect 2249 13060 2250 14480
rect 5370 14840 5371 16180
rect 6049 16180 9171 16181
rect 6049 14840 6050 16180
rect 5370 14480 6050 14840
rect 5370 13060 5371 14480
rect 2249 13059 5371 13060
rect 5560 11410 5880 14480
rect 6049 13060 6050 14480
rect 9170 13060 9171 16180
rect 6049 13059 9171 13060
rect -1970 11220 -1650 11350
rect -1790 9230 -1650 11220
rect 5250 11210 5880 11410
rect 1269 10930 1541 10931
rect 1269 10660 1270 10930
rect 1540 10660 1541 10930
rect 1269 10659 1541 10660
rect 2319 10930 2591 10931
rect 2319 10660 2320 10930
rect 2590 10660 2591 10930
rect 2319 10659 2591 10660
rect -901 10430 -649 10431
rect -901 10180 -900 10430
rect -650 10180 -649 10430
rect -901 10179 -649 10180
rect 999 10420 1251 10421
rect 999 10170 1000 10420
rect 1250 10170 1251 10420
rect 999 10169 1251 10170
rect 2579 10420 2831 10421
rect 2579 10170 2580 10420
rect 2830 10170 2831 10420
rect 2579 10169 2831 10170
rect 4479 10420 4731 10421
rect 4479 10170 4480 10420
rect 4730 10170 4731 10420
rect 4479 10169 4731 10170
rect -1790 9160 -1760 9230
rect -1690 9160 -1650 9230
rect -1790 9130 -1650 9160
rect 1269 9290 1541 9291
rect 1269 9020 1270 9290
rect 1540 9020 1541 9290
rect 1269 9019 1541 9020
rect 2319 9290 2591 9291
rect 2319 9020 2320 9290
rect 2590 9020 2591 9290
rect 5250 9230 5390 11210
rect 5250 9160 5290 9230
rect 5360 9160 5390 9230
rect 5250 9130 5390 9160
rect 2319 9019 2591 9020
rect 599 8770 861 8771
rect 599 8510 600 8770
rect 860 8510 861 8770
rect 599 8509 861 8510
rect 1869 8770 2131 8771
rect 1869 8510 1870 8770
rect 2130 8510 2131 8770
rect 1869 8509 2131 8510
rect 3129 8770 3391 8771
rect 3129 8510 3130 8770
rect 3390 8510 3391 8770
rect 3129 8509 3391 8510
rect 1039 7680 1301 7681
rect 1039 7420 1040 7680
rect 1300 7420 1301 7680
rect 1039 7419 1301 7420
rect 2539 7680 2801 7681
rect 2539 7420 2540 7680
rect 2800 7420 2801 7680
rect 2539 7419 2801 7420
rect 599 7220 861 7221
rect 599 6960 600 7220
rect 860 6960 861 7220
rect 599 6959 861 6960
rect 1869 7220 2131 7221
rect 1869 6960 1870 7220
rect 2130 6960 2131 7220
rect 1869 6959 2131 6960
rect 3129 7220 3391 7221
rect 3129 6960 3130 7220
rect 3390 6960 3391 7220
rect 3129 6959 3391 6960
rect 1779 4580 2041 4581
rect 1779 4320 1780 4580
rect 2040 4320 2041 4580
rect 1779 4319 2041 4320
rect 1779 3060 2041 3061
rect 1779 2800 1780 3060
rect 2040 2800 2041 3060
rect 1779 2799 2041 2800
rect 759 1960 1011 1961
rect 759 1710 760 1960
rect 1010 1710 1011 1960
rect 759 1709 1011 1710
rect 2819 1960 3071 1961
rect 2819 1710 2820 1960
rect 3070 1710 3071 1960
rect 2819 1709 3071 1710
rect 1789 1540 2041 1541
rect 1789 1290 1790 1540
rect 2040 1290 2041 1540
rect 1789 1289 2041 1290
rect -1351 1270 -759 1271
rect -1351 850 -1350 1270
rect -760 850 -759 1270
rect 4609 1200 5101 1201
rect 4609 940 4610 1200
rect 5100 940 5101 1200
rect 4609 939 5101 940
rect -1351 849 -759 850
rect 499 440 751 441
rect 499 190 500 440
rect 750 190 751 440
rect 499 189 751 190
rect 3079 440 3331 441
rect 3079 190 3080 440
rect 3330 190 3331 440
rect 3079 189 3331 190
rect 1789 10 2041 11
rect 1789 -240 1790 10
rect 2040 -240 2041 10
rect 1789 -241 2041 -240
<< via4 >>
rect 1270 10660 1540 10930
rect 2320 10660 2590 10930
rect -900 10180 -650 10430
rect 1000 10170 1250 10420
rect 2580 10170 2830 10420
rect 4480 10170 4730 10420
rect 1270 9020 1540 9290
rect 2320 9020 2590 9290
rect 600 8510 860 8770
rect 1870 8510 2130 8770
rect 3130 8510 3390 8770
rect 1040 7420 1300 7680
rect 2540 7420 2800 7680
rect 600 6960 860 7220
rect 1870 6960 2130 7220
rect 3130 6960 3390 7220
rect 1780 4320 2040 4580
rect 1780 2800 2040 3060
rect 760 1710 1010 1960
rect 2820 1710 3070 1960
rect 1790 1290 2040 1540
rect -1350 850 -760 1270
rect 4610 940 5100 1200
rect 500 190 750 440
rect 3080 190 3330 440
rect 1790 -240 2040 10
<< metal5 >>
rect 1240 10930 2620 10980
rect 1240 10660 1270 10930
rect 1540 10660 2320 10930
rect 2590 10660 2620 10930
rect 1240 10460 2620 10660
rect -930 10430 4770 10460
rect -930 10180 -900 10430
rect -650 10420 4770 10430
rect -650 10180 1000 10420
rect -930 10170 1000 10180
rect 1250 10170 2580 10420
rect 2830 10170 4480 10420
rect 4730 10170 4770 10420
rect -930 10130 4770 10170
rect 1240 9290 2620 10130
rect 1240 9020 1270 9290
rect 1540 9020 2320 9290
rect 2590 9020 2620 9290
rect 1240 8800 2620 9020
rect 450 8770 3430 8800
rect 450 8510 600 8770
rect 860 8510 1870 8770
rect 2130 8510 3130 8770
rect 3390 8510 3430 8770
rect 450 8480 3430 8510
rect 1240 7710 2620 8480
rect 1010 7680 2830 7710
rect 1010 7420 1040 7680
rect 1300 7420 2540 7680
rect 2800 7420 2830 7680
rect 1010 7250 2830 7420
rect 560 7220 3430 7250
rect 560 6960 600 7220
rect 860 6960 1870 7220
rect 2130 6960 3130 7220
rect 3390 6960 3430 7220
rect 560 6930 3430 6960
rect 1690 4580 2130 4620
rect 1690 4320 1780 4580
rect 2040 4320 2130 4580
rect 1690 3060 2130 4320
rect 1690 2800 1780 3060
rect 2040 2800 2130 3060
rect 1690 2000 2130 2800
rect -920 1960 4720 2000
rect -920 1710 760 1960
rect 1010 1710 2820 1960
rect 3070 1710 4720 1960
rect -920 1540 4720 1710
rect -920 1410 1790 1540
rect -1350 1294 1790 1410
rect -1374 1290 1790 1294
rect 2040 1290 4720 1540
rect -1374 1270 5130 1290
rect -1374 850 -1350 1270
rect -760 1200 5130 1270
rect -760 940 4610 1200
rect 5100 940 5130 1200
rect -760 880 5130 940
rect -760 850 4720 880
rect -1374 826 4720 850
rect -1350 610 4720 826
rect -920 440 4720 610
rect -920 190 500 440
rect 750 190 3080 440
rect 3330 190 4720 440
rect -920 150 4720 190
rect 1700 10 2140 150
rect 1700 -240 1790 10
rect 2040 -240 2140 10
rect 1700 -310 2140 -240
<< res5p73 >>
rect -4617 10271 -2613 11421
rect 7113 10271 9117 11421
rect -4617 8811 -2613 9961
rect 7113 8811 9117 9961
<< labels >>
rlabel metal5 4480 1040 4480 1040 1 Vss
port 1 n
rlabel metal5 1900 10860 1900 10860 1 Vdd
port 2 n
rlabel metal2 -330 2180 -330 2180 1 Vmirror
port 3 n
rlabel metal1 2660 5760 2660 5760 1 Vp
port 4 n
rlabel metal1 2670 4230 2670 4230 1 Vn
port 5 n
rlabel metal1 5890 10060 5890 10060 1 Vmid
port 6 n
rlabel metal2 4910 9070 4910 9070 1 Vout
port 7 n
<< end >>
