magic
tech sky130A
magscale 1 2
timestamp 1683391037
<< nwell >>
rect -1826 -719 1826 719
<< pmos >>
rect -1630 -500 -1530 500
rect -1472 -500 -1372 500
rect -1314 -500 -1214 500
rect -1156 -500 -1056 500
rect -998 -500 -898 500
rect -840 -500 -740 500
rect -682 -500 -582 500
rect -524 -500 -424 500
rect -366 -500 -266 500
rect -208 -500 -108 500
rect -50 -500 50 500
rect 108 -500 208 500
rect 266 -500 366 500
rect 424 -500 524 500
rect 582 -500 682 500
rect 740 -500 840 500
rect 898 -500 998 500
rect 1056 -500 1156 500
rect 1214 -500 1314 500
rect 1372 -500 1472 500
rect 1530 -500 1630 500
<< pdiff >>
rect -1688 488 -1630 500
rect -1688 -488 -1676 488
rect -1642 -488 -1630 488
rect -1688 -500 -1630 -488
rect -1530 488 -1472 500
rect -1530 -488 -1518 488
rect -1484 -488 -1472 488
rect -1530 -500 -1472 -488
rect -1372 488 -1314 500
rect -1372 -488 -1360 488
rect -1326 -488 -1314 488
rect -1372 -500 -1314 -488
rect -1214 488 -1156 500
rect -1214 -488 -1202 488
rect -1168 -488 -1156 488
rect -1214 -500 -1156 -488
rect -1056 488 -998 500
rect -1056 -488 -1044 488
rect -1010 -488 -998 488
rect -1056 -500 -998 -488
rect -898 488 -840 500
rect -898 -488 -886 488
rect -852 -488 -840 488
rect -898 -500 -840 -488
rect -740 488 -682 500
rect -740 -488 -728 488
rect -694 -488 -682 488
rect -740 -500 -682 -488
rect -582 488 -524 500
rect -582 -488 -570 488
rect -536 -488 -524 488
rect -582 -500 -524 -488
rect -424 488 -366 500
rect -424 -488 -412 488
rect -378 -488 -366 488
rect -424 -500 -366 -488
rect -266 488 -208 500
rect -266 -488 -254 488
rect -220 -488 -208 488
rect -266 -500 -208 -488
rect -108 488 -50 500
rect -108 -488 -96 488
rect -62 -488 -50 488
rect -108 -500 -50 -488
rect 50 488 108 500
rect 50 -488 62 488
rect 96 -488 108 488
rect 50 -500 108 -488
rect 208 488 266 500
rect 208 -488 220 488
rect 254 -488 266 488
rect 208 -500 266 -488
rect 366 488 424 500
rect 366 -488 378 488
rect 412 -488 424 488
rect 366 -500 424 -488
rect 524 488 582 500
rect 524 -488 536 488
rect 570 -488 582 488
rect 524 -500 582 -488
rect 682 488 740 500
rect 682 -488 694 488
rect 728 -488 740 488
rect 682 -500 740 -488
rect 840 488 898 500
rect 840 -488 852 488
rect 886 -488 898 488
rect 840 -500 898 -488
rect 998 488 1056 500
rect 998 -488 1010 488
rect 1044 -488 1056 488
rect 998 -500 1056 -488
rect 1156 488 1214 500
rect 1156 -488 1168 488
rect 1202 -488 1214 488
rect 1156 -500 1214 -488
rect 1314 488 1372 500
rect 1314 -488 1326 488
rect 1360 -488 1372 488
rect 1314 -500 1372 -488
rect 1472 488 1530 500
rect 1472 -488 1484 488
rect 1518 -488 1530 488
rect 1472 -500 1530 -488
rect 1630 488 1688 500
rect 1630 -488 1642 488
rect 1676 -488 1688 488
rect 1630 -500 1688 -488
<< pdiffc >>
rect -1676 -488 -1642 488
rect -1518 -488 -1484 488
rect -1360 -488 -1326 488
rect -1202 -488 -1168 488
rect -1044 -488 -1010 488
rect -886 -488 -852 488
rect -728 -488 -694 488
rect -570 -488 -536 488
rect -412 -488 -378 488
rect -254 -488 -220 488
rect -96 -488 -62 488
rect 62 -488 96 488
rect 220 -488 254 488
rect 378 -488 412 488
rect 536 -488 570 488
rect 694 -488 728 488
rect 852 -488 886 488
rect 1010 -488 1044 488
rect 1168 -488 1202 488
rect 1326 -488 1360 488
rect 1484 -488 1518 488
rect 1642 -488 1676 488
<< nsubdiff >>
rect -1790 649 -1694 683
rect 1694 649 1790 683
rect -1790 587 -1756 649
rect 1756 587 1790 649
rect -1790 -649 -1756 -587
rect 1756 -649 1790 -587
rect -1790 -683 -1694 -649
rect 1694 -683 1790 -649
<< nsubdiffcont >>
rect -1694 649 1694 683
rect -1790 -587 -1756 587
rect 1756 -587 1790 587
rect -1694 -683 1694 -649
<< poly >>
rect -1630 581 -1530 597
rect -1630 547 -1614 581
rect -1546 547 -1530 581
rect -1630 500 -1530 547
rect -1472 581 -1372 597
rect -1472 547 -1456 581
rect -1388 547 -1372 581
rect -1472 500 -1372 547
rect -1314 581 -1214 597
rect -1314 547 -1298 581
rect -1230 547 -1214 581
rect -1314 500 -1214 547
rect -1156 581 -1056 597
rect -1156 547 -1140 581
rect -1072 547 -1056 581
rect -1156 500 -1056 547
rect -998 581 -898 597
rect -998 547 -982 581
rect -914 547 -898 581
rect -998 500 -898 547
rect -840 581 -740 597
rect -840 547 -824 581
rect -756 547 -740 581
rect -840 500 -740 547
rect -682 581 -582 597
rect -682 547 -666 581
rect -598 547 -582 581
rect -682 500 -582 547
rect -524 581 -424 597
rect -524 547 -508 581
rect -440 547 -424 581
rect -524 500 -424 547
rect -366 581 -266 597
rect -366 547 -350 581
rect -282 547 -266 581
rect -366 500 -266 547
rect -208 581 -108 597
rect -208 547 -192 581
rect -124 547 -108 581
rect -208 500 -108 547
rect -50 581 50 597
rect -50 547 -34 581
rect 34 547 50 581
rect -50 500 50 547
rect 108 581 208 597
rect 108 547 124 581
rect 192 547 208 581
rect 108 500 208 547
rect 266 581 366 597
rect 266 547 282 581
rect 350 547 366 581
rect 266 500 366 547
rect 424 581 524 597
rect 424 547 440 581
rect 508 547 524 581
rect 424 500 524 547
rect 582 581 682 597
rect 582 547 598 581
rect 666 547 682 581
rect 582 500 682 547
rect 740 581 840 597
rect 740 547 756 581
rect 824 547 840 581
rect 740 500 840 547
rect 898 581 998 597
rect 898 547 914 581
rect 982 547 998 581
rect 898 500 998 547
rect 1056 581 1156 597
rect 1056 547 1072 581
rect 1140 547 1156 581
rect 1056 500 1156 547
rect 1214 581 1314 597
rect 1214 547 1230 581
rect 1298 547 1314 581
rect 1214 500 1314 547
rect 1372 581 1472 597
rect 1372 547 1388 581
rect 1456 547 1472 581
rect 1372 500 1472 547
rect 1530 581 1630 597
rect 1530 547 1546 581
rect 1614 547 1630 581
rect 1530 500 1630 547
rect -1630 -547 -1530 -500
rect -1630 -581 -1614 -547
rect -1546 -581 -1530 -547
rect -1630 -597 -1530 -581
rect -1472 -547 -1372 -500
rect -1472 -581 -1456 -547
rect -1388 -581 -1372 -547
rect -1472 -597 -1372 -581
rect -1314 -547 -1214 -500
rect -1314 -581 -1298 -547
rect -1230 -581 -1214 -547
rect -1314 -597 -1214 -581
rect -1156 -547 -1056 -500
rect -1156 -581 -1140 -547
rect -1072 -581 -1056 -547
rect -1156 -597 -1056 -581
rect -998 -547 -898 -500
rect -998 -581 -982 -547
rect -914 -581 -898 -547
rect -998 -597 -898 -581
rect -840 -547 -740 -500
rect -840 -581 -824 -547
rect -756 -581 -740 -547
rect -840 -597 -740 -581
rect -682 -547 -582 -500
rect -682 -581 -666 -547
rect -598 -581 -582 -547
rect -682 -597 -582 -581
rect -524 -547 -424 -500
rect -524 -581 -508 -547
rect -440 -581 -424 -547
rect -524 -597 -424 -581
rect -366 -547 -266 -500
rect -366 -581 -350 -547
rect -282 -581 -266 -547
rect -366 -597 -266 -581
rect -208 -547 -108 -500
rect -208 -581 -192 -547
rect -124 -581 -108 -547
rect -208 -597 -108 -581
rect -50 -547 50 -500
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -50 -597 50 -581
rect 108 -547 208 -500
rect 108 -581 124 -547
rect 192 -581 208 -547
rect 108 -597 208 -581
rect 266 -547 366 -500
rect 266 -581 282 -547
rect 350 -581 366 -547
rect 266 -597 366 -581
rect 424 -547 524 -500
rect 424 -581 440 -547
rect 508 -581 524 -547
rect 424 -597 524 -581
rect 582 -547 682 -500
rect 582 -581 598 -547
rect 666 -581 682 -547
rect 582 -597 682 -581
rect 740 -547 840 -500
rect 740 -581 756 -547
rect 824 -581 840 -547
rect 740 -597 840 -581
rect 898 -547 998 -500
rect 898 -581 914 -547
rect 982 -581 998 -547
rect 898 -597 998 -581
rect 1056 -547 1156 -500
rect 1056 -581 1072 -547
rect 1140 -581 1156 -547
rect 1056 -597 1156 -581
rect 1214 -547 1314 -500
rect 1214 -581 1230 -547
rect 1298 -581 1314 -547
rect 1214 -597 1314 -581
rect 1372 -547 1472 -500
rect 1372 -581 1388 -547
rect 1456 -581 1472 -547
rect 1372 -597 1472 -581
rect 1530 -547 1630 -500
rect 1530 -581 1546 -547
rect 1614 -581 1630 -547
rect 1530 -597 1630 -581
<< polycont >>
rect -1614 547 -1546 581
rect -1456 547 -1388 581
rect -1298 547 -1230 581
rect -1140 547 -1072 581
rect -982 547 -914 581
rect -824 547 -756 581
rect -666 547 -598 581
rect -508 547 -440 581
rect -350 547 -282 581
rect -192 547 -124 581
rect -34 547 34 581
rect 124 547 192 581
rect 282 547 350 581
rect 440 547 508 581
rect 598 547 666 581
rect 756 547 824 581
rect 914 547 982 581
rect 1072 547 1140 581
rect 1230 547 1298 581
rect 1388 547 1456 581
rect 1546 547 1614 581
rect -1614 -581 -1546 -547
rect -1456 -581 -1388 -547
rect -1298 -581 -1230 -547
rect -1140 -581 -1072 -547
rect -982 -581 -914 -547
rect -824 -581 -756 -547
rect -666 -581 -598 -547
rect -508 -581 -440 -547
rect -350 -581 -282 -547
rect -192 -581 -124 -547
rect -34 -581 34 -547
rect 124 -581 192 -547
rect 282 -581 350 -547
rect 440 -581 508 -547
rect 598 -581 666 -547
rect 756 -581 824 -547
rect 914 -581 982 -547
rect 1072 -581 1140 -547
rect 1230 -581 1298 -547
rect 1388 -581 1456 -547
rect 1546 -581 1614 -547
<< locali >>
rect -1790 649 -1694 683
rect 1694 649 1790 683
rect -1790 587 -1756 649
rect 1756 587 1790 649
rect -1630 547 -1614 581
rect -1546 547 -1530 581
rect -1472 547 -1456 581
rect -1388 547 -1372 581
rect -1314 547 -1298 581
rect -1230 547 -1214 581
rect -1156 547 -1140 581
rect -1072 547 -1056 581
rect -998 547 -982 581
rect -914 547 -898 581
rect -840 547 -824 581
rect -756 547 -740 581
rect -682 547 -666 581
rect -598 547 -582 581
rect -524 547 -508 581
rect -440 547 -424 581
rect -366 547 -350 581
rect -282 547 -266 581
rect -208 547 -192 581
rect -124 547 -108 581
rect -50 547 -34 581
rect 34 547 50 581
rect 108 547 124 581
rect 192 547 208 581
rect 266 547 282 581
rect 350 547 366 581
rect 424 547 440 581
rect 508 547 524 581
rect 582 547 598 581
rect 666 547 682 581
rect 740 547 756 581
rect 824 547 840 581
rect 898 547 914 581
rect 982 547 998 581
rect 1056 547 1072 581
rect 1140 547 1156 581
rect 1214 547 1230 581
rect 1298 547 1314 581
rect 1372 547 1388 581
rect 1456 547 1472 581
rect 1530 547 1546 581
rect 1614 547 1630 581
rect -1676 488 -1642 504
rect -1676 -504 -1642 -488
rect -1518 488 -1484 504
rect -1518 -504 -1484 -488
rect -1360 488 -1326 504
rect -1360 -504 -1326 -488
rect -1202 488 -1168 504
rect -1202 -504 -1168 -488
rect -1044 488 -1010 504
rect -1044 -504 -1010 -488
rect -886 488 -852 504
rect -886 -504 -852 -488
rect -728 488 -694 504
rect -728 -504 -694 -488
rect -570 488 -536 504
rect -570 -504 -536 -488
rect -412 488 -378 504
rect -412 -504 -378 -488
rect -254 488 -220 504
rect -254 -504 -220 -488
rect -96 488 -62 504
rect -96 -504 -62 -488
rect 62 488 96 504
rect 62 -504 96 -488
rect 220 488 254 504
rect 220 -504 254 -488
rect 378 488 412 504
rect 378 -504 412 -488
rect 536 488 570 504
rect 536 -504 570 -488
rect 694 488 728 504
rect 694 -504 728 -488
rect 852 488 886 504
rect 852 -504 886 -488
rect 1010 488 1044 504
rect 1010 -504 1044 -488
rect 1168 488 1202 504
rect 1168 -504 1202 -488
rect 1326 488 1360 504
rect 1326 -504 1360 -488
rect 1484 488 1518 504
rect 1484 -504 1518 -488
rect 1642 488 1676 504
rect 1642 -504 1676 -488
rect -1630 -581 -1614 -547
rect -1546 -581 -1530 -547
rect -1472 -581 -1456 -547
rect -1388 -581 -1372 -547
rect -1314 -581 -1298 -547
rect -1230 -581 -1214 -547
rect -1156 -581 -1140 -547
rect -1072 -581 -1056 -547
rect -998 -581 -982 -547
rect -914 -581 -898 -547
rect -840 -581 -824 -547
rect -756 -581 -740 -547
rect -682 -581 -666 -547
rect -598 -581 -582 -547
rect -524 -581 -508 -547
rect -440 -581 -424 -547
rect -366 -581 -350 -547
rect -282 -581 -266 -547
rect -208 -581 -192 -547
rect -124 -581 -108 -547
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect 108 -581 124 -547
rect 192 -581 208 -547
rect 266 -581 282 -547
rect 350 -581 366 -547
rect 424 -581 440 -547
rect 508 -581 524 -547
rect 582 -581 598 -547
rect 666 -581 682 -547
rect 740 -581 756 -547
rect 824 -581 840 -547
rect 898 -581 914 -547
rect 982 -581 998 -547
rect 1056 -581 1072 -547
rect 1140 -581 1156 -547
rect 1214 -581 1230 -547
rect 1298 -581 1314 -547
rect 1372 -581 1388 -547
rect 1456 -581 1472 -547
rect 1530 -581 1546 -547
rect 1614 -581 1630 -547
rect -1790 -649 -1756 -587
rect 1756 -649 1790 -587
rect -1790 -683 -1694 -649
rect 1694 -683 1790 -649
<< viali >>
rect -1614 547 -1546 581
rect -1456 547 -1388 581
rect -1298 547 -1230 581
rect -1140 547 -1072 581
rect -982 547 -914 581
rect -824 547 -756 581
rect -666 547 -598 581
rect -508 547 -440 581
rect -350 547 -282 581
rect -192 547 -124 581
rect -34 547 34 581
rect 124 547 192 581
rect 282 547 350 581
rect 440 547 508 581
rect 598 547 666 581
rect 756 547 824 581
rect 914 547 982 581
rect 1072 547 1140 581
rect 1230 547 1298 581
rect 1388 547 1456 581
rect 1546 547 1614 581
rect -1676 -488 -1642 488
rect -1518 -488 -1484 488
rect -1360 -488 -1326 488
rect -1202 -488 -1168 488
rect -1044 -488 -1010 488
rect -886 -488 -852 488
rect -728 -488 -694 488
rect -570 -488 -536 488
rect -412 -488 -378 488
rect -254 -488 -220 488
rect -96 -488 -62 488
rect 62 -488 96 488
rect 220 -488 254 488
rect 378 -488 412 488
rect 536 -488 570 488
rect 694 -488 728 488
rect 852 -488 886 488
rect 1010 -488 1044 488
rect 1168 -488 1202 488
rect 1326 -488 1360 488
rect 1484 -488 1518 488
rect 1642 -488 1676 488
rect -1614 -581 -1546 -547
rect -1456 -581 -1388 -547
rect -1298 -581 -1230 -547
rect -1140 -581 -1072 -547
rect -982 -581 -914 -547
rect -824 -581 -756 -547
rect -666 -581 -598 -547
rect -508 -581 -440 -547
rect -350 -581 -282 -547
rect -192 -581 -124 -547
rect -34 -581 34 -547
rect 124 -581 192 -547
rect 282 -581 350 -547
rect 440 -581 508 -547
rect 598 -581 666 -547
rect 756 -581 824 -547
rect 914 -581 982 -547
rect 1072 -581 1140 -547
rect 1230 -581 1298 -547
rect 1388 -581 1456 -547
rect 1546 -581 1614 -547
<< metal1 >>
rect -1626 581 -1534 587
rect -1626 547 -1614 581
rect -1546 547 -1534 581
rect -1626 541 -1534 547
rect -1468 581 -1376 587
rect -1468 547 -1456 581
rect -1388 547 -1376 581
rect -1468 541 -1376 547
rect -1310 581 -1218 587
rect -1310 547 -1298 581
rect -1230 547 -1218 581
rect -1310 541 -1218 547
rect -1152 581 -1060 587
rect -1152 547 -1140 581
rect -1072 547 -1060 581
rect -1152 541 -1060 547
rect -994 581 -902 587
rect -994 547 -982 581
rect -914 547 -902 581
rect -994 541 -902 547
rect -836 581 -744 587
rect -836 547 -824 581
rect -756 547 -744 581
rect -836 541 -744 547
rect -678 581 -586 587
rect -678 547 -666 581
rect -598 547 -586 581
rect -678 541 -586 547
rect -520 581 -428 587
rect -520 547 -508 581
rect -440 547 -428 581
rect -520 541 -428 547
rect -362 581 -270 587
rect -362 547 -350 581
rect -282 547 -270 581
rect -362 541 -270 547
rect -204 581 -112 587
rect -204 547 -192 581
rect -124 547 -112 581
rect -204 541 -112 547
rect -46 581 46 587
rect -46 547 -34 581
rect 34 547 46 581
rect -46 541 46 547
rect 112 581 204 587
rect 112 547 124 581
rect 192 547 204 581
rect 112 541 204 547
rect 270 581 362 587
rect 270 547 282 581
rect 350 547 362 581
rect 270 541 362 547
rect 428 581 520 587
rect 428 547 440 581
rect 508 547 520 581
rect 428 541 520 547
rect 586 581 678 587
rect 586 547 598 581
rect 666 547 678 581
rect 586 541 678 547
rect 744 581 836 587
rect 744 547 756 581
rect 824 547 836 581
rect 744 541 836 547
rect 902 581 994 587
rect 902 547 914 581
rect 982 547 994 581
rect 902 541 994 547
rect 1060 581 1152 587
rect 1060 547 1072 581
rect 1140 547 1152 581
rect 1060 541 1152 547
rect 1218 581 1310 587
rect 1218 547 1230 581
rect 1298 547 1310 581
rect 1218 541 1310 547
rect 1376 581 1468 587
rect 1376 547 1388 581
rect 1456 547 1468 581
rect 1376 541 1468 547
rect 1534 581 1626 587
rect 1534 547 1546 581
rect 1614 547 1626 581
rect 1534 541 1626 547
rect -1682 488 -1636 500
rect -1682 -488 -1676 488
rect -1642 -488 -1636 488
rect -1682 -500 -1636 -488
rect -1524 488 -1478 500
rect -1524 -488 -1518 488
rect -1484 -488 -1478 488
rect -1524 -500 -1478 -488
rect -1366 488 -1320 500
rect -1366 -488 -1360 488
rect -1326 -488 -1320 488
rect -1366 -500 -1320 -488
rect -1208 488 -1162 500
rect -1208 -488 -1202 488
rect -1168 -488 -1162 488
rect -1208 -500 -1162 -488
rect -1050 488 -1004 500
rect -1050 -488 -1044 488
rect -1010 -488 -1004 488
rect -1050 -500 -1004 -488
rect -892 488 -846 500
rect -892 -488 -886 488
rect -852 -488 -846 488
rect -892 -500 -846 -488
rect -734 488 -688 500
rect -734 -488 -728 488
rect -694 -488 -688 488
rect -734 -500 -688 -488
rect -576 488 -530 500
rect -576 -488 -570 488
rect -536 -488 -530 488
rect -576 -500 -530 -488
rect -418 488 -372 500
rect -418 -488 -412 488
rect -378 -488 -372 488
rect -418 -500 -372 -488
rect -260 488 -214 500
rect -260 -488 -254 488
rect -220 -488 -214 488
rect -260 -500 -214 -488
rect -102 488 -56 500
rect -102 -488 -96 488
rect -62 -488 -56 488
rect -102 -500 -56 -488
rect 56 488 102 500
rect 56 -488 62 488
rect 96 -488 102 488
rect 56 -500 102 -488
rect 214 488 260 500
rect 214 -488 220 488
rect 254 -488 260 488
rect 214 -500 260 -488
rect 372 488 418 500
rect 372 -488 378 488
rect 412 -488 418 488
rect 372 -500 418 -488
rect 530 488 576 500
rect 530 -488 536 488
rect 570 -488 576 488
rect 530 -500 576 -488
rect 688 488 734 500
rect 688 -488 694 488
rect 728 -488 734 488
rect 688 -500 734 -488
rect 846 488 892 500
rect 846 -488 852 488
rect 886 -488 892 488
rect 846 -500 892 -488
rect 1004 488 1050 500
rect 1004 -488 1010 488
rect 1044 -488 1050 488
rect 1004 -500 1050 -488
rect 1162 488 1208 500
rect 1162 -488 1168 488
rect 1202 -488 1208 488
rect 1162 -500 1208 -488
rect 1320 488 1366 500
rect 1320 -488 1326 488
rect 1360 -488 1366 488
rect 1320 -500 1366 -488
rect 1478 488 1524 500
rect 1478 -488 1484 488
rect 1518 -488 1524 488
rect 1478 -500 1524 -488
rect 1636 488 1682 500
rect 1636 -488 1642 488
rect 1676 -488 1682 488
rect 1636 -500 1682 -488
rect -1626 -547 -1534 -541
rect -1626 -581 -1614 -547
rect -1546 -581 -1534 -547
rect -1626 -587 -1534 -581
rect -1468 -547 -1376 -541
rect -1468 -581 -1456 -547
rect -1388 -581 -1376 -547
rect -1468 -587 -1376 -581
rect -1310 -547 -1218 -541
rect -1310 -581 -1298 -547
rect -1230 -581 -1218 -547
rect -1310 -587 -1218 -581
rect -1152 -547 -1060 -541
rect -1152 -581 -1140 -547
rect -1072 -581 -1060 -547
rect -1152 -587 -1060 -581
rect -994 -547 -902 -541
rect -994 -581 -982 -547
rect -914 -581 -902 -547
rect -994 -587 -902 -581
rect -836 -547 -744 -541
rect -836 -581 -824 -547
rect -756 -581 -744 -547
rect -836 -587 -744 -581
rect -678 -547 -586 -541
rect -678 -581 -666 -547
rect -598 -581 -586 -547
rect -678 -587 -586 -581
rect -520 -547 -428 -541
rect -520 -581 -508 -547
rect -440 -581 -428 -547
rect -520 -587 -428 -581
rect -362 -547 -270 -541
rect -362 -581 -350 -547
rect -282 -581 -270 -547
rect -362 -587 -270 -581
rect -204 -547 -112 -541
rect -204 -581 -192 -547
rect -124 -581 -112 -547
rect -204 -587 -112 -581
rect -46 -547 46 -541
rect -46 -581 -34 -547
rect 34 -581 46 -547
rect -46 -587 46 -581
rect 112 -547 204 -541
rect 112 -581 124 -547
rect 192 -581 204 -547
rect 112 -587 204 -581
rect 270 -547 362 -541
rect 270 -581 282 -547
rect 350 -581 362 -547
rect 270 -587 362 -581
rect 428 -547 520 -541
rect 428 -581 440 -547
rect 508 -581 520 -547
rect 428 -587 520 -581
rect 586 -547 678 -541
rect 586 -581 598 -547
rect 666 -581 678 -547
rect 586 -587 678 -581
rect 744 -547 836 -541
rect 744 -581 756 -547
rect 824 -581 836 -547
rect 744 -587 836 -581
rect 902 -547 994 -541
rect 902 -581 914 -547
rect 982 -581 994 -547
rect 902 -587 994 -581
rect 1060 -547 1152 -541
rect 1060 -581 1072 -547
rect 1140 -581 1152 -547
rect 1060 -587 1152 -581
rect 1218 -547 1310 -541
rect 1218 -581 1230 -547
rect 1298 -581 1310 -547
rect 1218 -587 1310 -581
rect 1376 -547 1468 -541
rect 1376 -581 1388 -547
rect 1456 -581 1468 -547
rect 1376 -587 1468 -581
rect 1534 -547 1626 -541
rect 1534 -581 1546 -547
rect 1614 -581 1626 -547
rect 1534 -587 1626 -581
<< properties >>
string FIXED_BBOX -1773 -666 1773 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 0.5 m 1 nf 21 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
