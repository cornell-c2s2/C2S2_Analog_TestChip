magic
tech sky130A
magscale 1 2
timestamp 1683899510
<< metal4 >>
rect -2750 480 2750 537
rect -2750 -537 2750 -480
<< rmetal4 >>
rect -2750 -480 2750 480
<< properties >>
string gencell sky130_fd_pr__res_generic_m4
string library sky130
string parameters w 27.5 l 4.8 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 8.203m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
