magic
tech sky130A
magscale 1 2
timestamp 1682777243
<< nwell >>
rect -2138 -2138 2138 2138
<< pwell >>
rect -2276 2138 2276 2276
rect -2276 -2138 -2138 2138
rect 2138 -2138 2276 2138
rect -2276 -2276 2276 -2138
<< psubdiff >>
rect -2240 2206 -2144 2240
rect 2144 2206 2240 2240
rect -2240 2144 -2206 2206
rect 2206 2144 2240 2206
rect -2240 -2206 -2206 -2144
rect 2206 -2206 2240 -2144
rect -2240 -2240 -2144 -2206
rect 2144 -2240 2240 -2206
<< nsubdiff >>
rect -2102 2068 -2006 2102
rect 2006 2068 2102 2102
rect -2102 2006 -2068 2068
rect 2068 2006 2102 2068
rect -2102 -2068 -2068 -2006
rect 2068 -2068 2102 -2006
rect -2102 -2102 -2006 -2068
rect 2006 -2102 2102 -2068
<< psubdiffcont >>
rect -2144 2206 2144 2240
rect -2240 -2144 -2206 2144
rect 2206 -2144 2240 2144
rect -2144 -2240 2144 -2206
<< nsubdiffcont >>
rect -2006 2068 2006 2102
rect -2102 -2006 -2068 2006
rect 2068 -2006 2102 2006
rect -2006 -2102 2006 -2068
<< pdiode >>
rect -2000 1988 2000 2000
rect -2000 -1988 -1988 1988
rect 1988 -1988 2000 1988
rect -2000 -2000 2000 -1988
<< pdiodec >>
rect -1988 -1988 1988 1988
<< locali >>
rect -2240 2206 -2144 2240
rect 2144 2206 2240 2240
rect -2240 2144 -2206 2206
rect 2206 2144 2240 2206
rect -2102 2068 -2006 2102
rect 2006 2068 2102 2102
rect -2102 2006 -2068 2068
rect 2068 2006 2102 2068
rect -2004 -1988 -1988 1988
rect 1988 -1988 2004 1988
rect -2102 -2068 -2068 -2006
rect 2068 -2068 2102 -2006
rect -2102 -2102 -2006 -2068
rect 2006 -2102 2102 -2068
rect -2240 -2206 -2206 -2144
rect 2206 -2206 2240 -2144
rect -2240 -2240 -2144 -2206
rect 2144 -2240 2240 -2206
<< viali >>
rect -552 2206 552 2240
rect -2240 -552 -2206 552
rect -517 2068 517 2102
rect -2102 -517 -2068 517
rect -1988 -1988 1988 1988
rect 2068 -517 2102 517
rect -517 -2102 517 -2068
rect 2206 -552 2240 552
rect -552 -2240 552 -2206
<< metal1 >>
rect -564 2240 564 2246
rect -564 2206 -552 2240
rect 552 2206 564 2240
rect -564 2200 564 2206
rect -529 2102 529 2108
rect -529 2068 -517 2102
rect 517 2068 529 2102
rect -529 2062 529 2068
rect -2000 1988 2000 1994
rect -2246 552 -2200 564
rect -2246 -552 -2240 552
rect -2206 -552 -2200 552
rect -2108 517 -2062 529
rect -2108 -517 -2102 517
rect -2068 -517 -2062 517
rect -2108 -529 -2062 -517
rect -2246 -564 -2200 -552
rect -2000 -1988 -1988 1988
rect 1988 -1988 2000 1988
rect 2200 552 2246 564
rect 2062 517 2108 529
rect 2062 -517 2068 517
rect 2102 -517 2108 517
rect 2062 -529 2108 -517
rect 2200 -552 2206 552
rect 2240 -552 2246 552
rect 2200 -564 2246 -552
rect -2000 -1994 2000 -1988
rect -529 -2068 529 -2062
rect -529 -2102 -517 -2068
rect 517 -2102 529 -2068
rect -529 -2108 529 -2102
rect -564 -2206 564 -2200
rect -564 -2240 -552 -2206
rect 552 -2240 564 -2206
rect -564 -2246 564 -2240
<< properties >>
string FIXED_BBOX -2085 -2085 2085 2085
string gencell sky130_fd_pr__diode_pd2nw_05v5
string library sky130
string parameters w 20 l 20 area 400.0 peri 80.0 nx 1 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 25 viagt 25 viagl 25 viagr 25
<< end >>
