magic
tech sky130A
magscale 1 2
timestamp 1676748949
<< nwell >>
rect -4170 1941 4040 3182
<< pwell >>
rect -835 1575 240 1625
<< metal1 >>
rect -3590 2960 3588 3030
rect -3678 2860 3670 2870
rect -3678 2790 -1720 2860
rect -1650 2790 -1500 2860
rect -1430 2790 1460 2860
rect 1530 2790 1700 2860
rect 1770 2790 3670 2860
rect -3678 2658 3670 2790
rect -3590 2370 3580 2450
rect -3680 2270 3676 2280
rect -3680 2200 -1720 2270
rect -1650 2200 -1500 2270
rect -1430 2200 1460 2270
rect 1530 2200 1700 2270
rect 1770 2200 3676 2270
rect -3680 2190 3676 2200
rect -3600 2110 -3590 2130
rect 3570 2110 3594 2130
rect -3600 2040 -560 2110
rect -490 2040 -450 2110
rect -380 2040 380 2110
rect 450 2040 490 2110
rect 560 2040 3594 2110
rect -3600 2030 3594 2040
rect -920 1550 900 1620
rect -920 1540 380 1550
rect -920 1470 -560 1540
rect -490 1470 -450 1540
rect -380 1480 380 1540
rect 450 1480 490 1550
rect 560 1480 900 1550
rect -380 1470 900 1480
rect -900 1390 900 1470
rect -550 1350 -390 1390
rect -80 1350 75 1390
rect 390 1350 545 1390
rect -840 1265 830 1320
rect 1440 1030 1790 1050
rect -1740 1010 1460 1030
rect -1740 940 -1720 1010
rect -1650 940 -1510 1010
rect -1440 960 1460 1010
rect 1530 960 1700 1030
rect 1770 960 1790 1030
rect -1440 940 1790 960
rect -1740 920 1460 940
rect -1740 850 -1720 920
rect -1650 850 -1510 920
rect -1440 870 1460 920
rect 1530 870 1700 940
rect 1770 870 1790 940
rect -1440 850 1790 870
rect -1740 820 -1410 850
rect -615 790 620 795
rect -615 780 -560 790
rect -620 720 -560 780
rect -490 720 -450 790
rect -380 720 380 790
rect 450 720 490 790
rect 560 780 620 790
rect 560 720 630 780
rect -620 710 630 720
rect -3550 490 3540 495
rect -3550 420 -1720 490
rect -1650 420 -1500 490
rect -1430 420 1460 490
rect 1530 420 1700 490
rect 1770 420 3540 490
rect -3620 340 3615 345
rect -3620 270 -560 340
rect -490 270 -450 340
rect -380 270 380 340
rect 450 270 490 340
rect 560 270 3615 340
rect -3620 260 3615 270
rect -3550 95 3540 170
rect -2060 -290 -1830 95
rect -750 -290 -520 95
rect 530 -290 760 95
rect 1790 -290 2020 95
rect -2500 -720 2540 -290
rect -2540 -18130 2540 -17640
<< via1 >>
rect -1720 2790 -1650 2860
rect -1500 2790 -1430 2860
rect 1460 2790 1530 2860
rect 1700 2790 1770 2860
rect -1720 2200 -1650 2270
rect -1500 2200 -1430 2270
rect 1460 2200 1530 2270
rect 1700 2200 1770 2270
rect -560 2040 -490 2110
rect -450 2040 -380 2110
rect 380 2040 450 2110
rect 490 2040 560 2110
rect -560 1470 -490 1540
rect -450 1470 -380 1540
rect 380 1480 450 1550
rect 490 1480 560 1550
rect -1720 940 -1650 1010
rect -1510 940 -1440 1010
rect 1460 960 1530 1030
rect 1700 960 1770 1030
rect -1720 850 -1650 920
rect -1510 850 -1440 920
rect 1460 870 1530 940
rect 1700 870 1770 940
rect -560 720 -490 790
rect -450 720 -380 790
rect 380 720 450 790
rect 490 720 560 790
rect -1720 420 -1650 490
rect -1500 420 -1430 490
rect 1460 420 1530 490
rect 1700 420 1770 490
rect -560 270 -490 340
rect -450 270 -380 340
rect 380 270 450 340
rect 490 270 560 340
<< metal2 >>
rect 1440 2860 1790 2870
rect -1740 2790 -1720 2860
rect -1650 2790 -1500 2860
rect -1430 2790 -1410 2860
rect -1740 2270 -1410 2790
rect -1740 2200 -1720 2270
rect -1650 2200 -1500 2270
rect -1430 2200 -1410 2270
rect -1740 1010 -1410 2200
rect 1440 2790 1460 2860
rect 1530 2790 1700 2860
rect 1770 2790 1790 2860
rect 1440 2270 1790 2790
rect 1440 2200 1460 2270
rect 1530 2200 1700 2270
rect 1770 2200 1790 2270
rect -1740 940 -1720 1010
rect -1650 940 -1510 1010
rect -1440 940 -1410 1010
rect -1740 920 -1410 940
rect -1740 850 -1720 920
rect -1650 850 -1510 920
rect -1440 850 -1410 920
rect -1740 490 -1410 850
rect -1740 420 -1720 490
rect -1650 420 -1500 490
rect -1430 420 -1410 490
rect -1740 410 -1410 420
rect -580 2110 -360 2120
rect -580 2040 -560 2110
rect -490 2040 -450 2110
rect -380 2040 -360 2110
rect -580 1540 -360 2040
rect -580 1470 -560 1540
rect -490 1470 -450 1540
rect -380 1470 -360 1540
rect -580 790 -360 1470
rect -580 720 -560 790
rect -490 720 -450 790
rect -380 720 -360 790
rect -580 340 -360 720
rect -580 270 -560 340
rect -490 270 -450 340
rect -380 270 -360 340
rect -580 200 -360 270
rect 360 2110 580 2130
rect 360 2040 380 2110
rect 450 2040 490 2110
rect 560 2040 580 2110
rect 360 1550 580 2040
rect 360 1480 380 1550
rect 450 1480 490 1550
rect 560 1480 580 1550
rect 360 790 580 1480
rect 360 720 380 790
rect 450 720 490 790
rect 560 720 580 790
rect 360 340 580 720
rect 1440 1030 1790 2200
rect 1440 960 1460 1030
rect 1530 960 1700 1030
rect 1770 960 1790 1030
rect 1440 940 1790 960
rect 1440 870 1460 940
rect 1530 870 1700 940
rect 1770 870 1790 940
rect 1440 490 1790 870
rect 1440 420 1460 490
rect 1530 420 1700 490
rect 1770 420 1790 490
rect 1440 390 1790 420
rect 360 270 380 340
rect 450 270 490 340
rect 560 270 580 340
rect 360 210 580 270
use sky130_fd_pr__nfet_01v8_GG6QWW  sky130_fd_pr__nfet_01v8_GG6QWW_0
timestamp 1676503286
transform 0 1 0 -1 0 296
box -296 -3755 296 3755
use sky130_fd_pr__nfet_01v8_JTC45A  sky130_fd_pr__nfet_01v8_JTC45A_0
timestamp 1676503286
transform 0 1 -3 -1 0 1446
box -296 -1037 296 1037
use sky130_fd_pr__nfet_01v8_N53VJN  sky130_fd_pr__nfet_01v8_N53VJN_0
timestamp 1676503286
transform 0 1 -1 -1 0 871
box -246 -819 246 819
use sky130_fd_pr__pfet_01v8_MKLXZC  sky130_fd_pr__pfet_01v8_MKLXZC_0
timestamp 1676746197
transform 0 1 -1 -1 0 2236
box -296 -3809 296 3809
use sky130_fd_pr__pfet_01v8_MKLXZC  sky130_fd_pr__pfet_01v8_MKLXZC_1
timestamp 1676746197
transform 0 1 -1 -1 0 2826
box -296 -3809 296 3809
use sky130_fd_pr__res_xhigh_po_5p73_EG97HE  sky130_fd_pr__res_xhigh_po_5p73_EG97HE_0
timestamp 1676748949
transform -1 0 1970 0 -1 -9192
box -575 -8902 575 8902
use sky130_fd_pr__res_xhigh_po_5p73_EG97HE  sky130_fd_pr__res_xhigh_po_5p73_EG97HE_1
timestamp 1676748949
transform -1 0 660 0 -1 -9192
box -575 -8902 575 8902
use sky130_fd_pr__res_xhigh_po_5p73_EG97HE  sky130_fd_pr__res_xhigh_po_5p73_EG97HE_2
timestamp 1676748949
transform -1 0 -650 0 -1 -9198
box -575 -8902 575 8902
use sky130_fd_pr__res_xhigh_po_5p73_EG97HE  sky130_fd_pr__res_xhigh_po_5p73_EG97HE_3
timestamp 1676748949
transform -1 0 -1920 0 -1 -9198
box -575 -8902 575 8902
<< end >>
