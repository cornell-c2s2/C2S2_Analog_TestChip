magic
tech sky130A
magscale 1 2
timestamp 1683899510
<< metal4 >>
rect -480 2750 480 2807
rect -480 -2807 480 -2750
<< rmetal4 >>
rect -480 -2750 480 2750
<< properties >>
string gencell sky130_fd_pr__res_generic_m4
string library sky130
string parameters w 4.8 l 27.5 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 269.27m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
