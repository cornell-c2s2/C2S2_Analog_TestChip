magic
tech sky130A
magscale 1 2
timestamp 1683391037
<< nwell >>
rect -6280 3640 6340 9080
<< locali >>
rect -2600 8050 -2340 8090
rect -2600 7980 -2590 8050
rect -2500 7980 -2450 8050
rect -2360 7980 -2340 8050
rect -2600 7940 -2340 7980
rect -130 8060 160 8090
rect -130 8050 50 8060
rect -130 7980 -110 8050
rect -20 7990 50 8050
rect 140 7990 160 8060
rect -20 7980 160 7990
rect -130 7940 160 7980
rect 2330 8060 2620 8090
rect 2330 7990 2350 8060
rect 2430 7990 2520 8060
rect 2600 7990 2620 8060
rect 2330 7950 2620 7990
rect -2610 7520 -2320 7540
rect -2610 7440 -2590 7520
rect -2510 7440 -2420 7520
rect -2340 7440 -2320 7520
rect -2610 7410 -2320 7440
rect -130 7520 160 7560
rect -130 7440 -110 7520
rect -30 7440 60 7520
rect 140 7440 160 7520
rect -130 7390 160 7440
rect 2330 7520 2620 7540
rect 2330 7440 2350 7520
rect 2430 7440 2520 7520
rect 2600 7440 2620 7520
rect 2330 7410 2620 7440
rect -2610 6360 -2320 6430
rect -2610 6280 -2590 6360
rect -2500 6280 -2430 6360
rect -2340 6280 -2320 6360
rect -2610 6250 -2320 6280
rect -130 6350 160 6450
rect -130 6280 -110 6350
rect -30 6280 60 6350
rect 140 6280 160 6350
rect -130 6250 160 6280
rect 2330 6350 2620 6450
rect 2330 6280 2350 6350
rect 2430 6280 2520 6350
rect 2600 6280 2620 6350
rect 2330 6250 2620 6280
rect -4470 5280 -4160 5330
rect -4470 5200 -4450 5280
rect -4360 5200 -4270 5280
rect -4180 5200 -4160 5280
rect -4470 5160 -4160 5200
rect -1940 5280 -1650 5300
rect -1940 5200 -1920 5280
rect -1830 5200 -1760 5280
rect -1670 5200 -1650 5280
rect -1940 5170 -1650 5200
rect 530 5280 820 5300
rect 530 5200 550 5280
rect 640 5200 710 5280
rect 800 5200 820 5280
rect 530 5170 820 5200
rect 2980 5280 3270 5300
rect 2980 5200 3000 5280
rect 3090 5200 3160 5280
rect 3250 5200 3270 5280
rect 2980 5170 3270 5200
rect 5480 5280 5770 5300
rect 5480 5200 5500 5280
rect 5590 5200 5660 5280
rect 5750 5200 5770 5280
rect 5480 5170 5770 5200
rect -8790 4750 -8700 4880
rect 8460 4740 8600 4850
rect -4470 4210 -4160 4240
rect -4470 4200 -4270 4210
rect -4470 4120 -4450 4200
rect -4360 4130 -4270 4200
rect -4180 4130 -4160 4210
rect -4360 4120 -4160 4130
rect -4470 4070 -4160 4120
rect -1940 4200 -1650 4220
rect -1940 4120 -1920 4200
rect -1830 4120 -1760 4200
rect -1670 4120 -1650 4200
rect -1940 4090 -1650 4120
rect 530 4200 820 4220
rect 530 4120 550 4200
rect 640 4120 710 4200
rect 800 4120 820 4200
rect 530 4090 820 4120
rect 2980 4200 3270 4220
rect 2980 4120 3000 4200
rect 3090 4120 3160 4200
rect 3250 4120 3270 4200
rect 2980 4090 3270 4120
rect 5480 4200 5770 4220
rect 5480 4120 5500 4200
rect 5590 4120 5660 4200
rect 5750 4120 5770 4200
rect 5480 4090 5770 4120
rect -3030 1790 -2860 1820
rect -3030 1700 -3000 1790
rect -2890 1700 -2860 1790
rect -3030 1670 -2860 1700
rect 1880 1790 2050 1830
rect 1880 1700 1910 1790
rect 2020 1700 2050 1790
rect 1880 1670 2050 1700
<< viali >>
rect -2600 9030 -2510 9100
rect -2430 9030 -2340 9100
rect -110 9030 -20 9100
rect 60 9030 150 9100
rect 2350 9030 2430 9110
rect 2520 9030 2600 9110
rect -2590 7980 -2500 8050
rect -2450 7980 -2360 8050
rect -110 7980 -20 8050
rect 50 7990 140 8060
rect 2350 7990 2430 8060
rect 2520 7990 2600 8060
rect -2590 7440 -2510 7520
rect -2420 7440 -2340 7520
rect -110 7440 -30 7520
rect 60 7440 140 7520
rect 2350 7440 2430 7520
rect 2520 7440 2600 7520
rect -2590 6280 -2500 6360
rect -2430 6280 -2340 6360
rect -110 6280 -30 6350
rect 60 6280 140 6350
rect 2350 6280 2430 6350
rect 2520 6280 2600 6350
rect -4450 5200 -4360 5280
rect -4270 5200 -4180 5280
rect -1920 5200 -1830 5280
rect -1760 5200 -1670 5280
rect 550 5200 640 5280
rect 710 5200 800 5280
rect 3000 5200 3090 5280
rect 3160 5200 3250 5280
rect 5500 5200 5590 5280
rect 5660 5200 5750 5280
rect -4450 4120 -4360 4200
rect -4270 4130 -4180 4210
rect -1920 4120 -1830 4200
rect -1760 4120 -1670 4200
rect 550 4120 640 4200
rect 710 4120 800 4200
rect 3000 4120 3090 4200
rect 3160 4120 3250 4200
rect 5500 4120 5590 4200
rect 5660 4120 5750 4200
rect -8810 3260 -8720 3390
rect -8600 3260 -8510 3390
rect 8500 3290 8570 3380
rect 8660 3290 8730 3380
rect -2290 2800 -2180 2910
rect -1430 2800 -1320 2910
rect -220 2800 -110 2910
rect 630 2800 740 2910
rect 2200 2800 2310 2910
rect 3080 2800 3190 2910
rect -3000 1700 -2890 1790
rect 1910 1700 2020 1790
rect -3060 490 -2940 590
rect -1840 490 -1720 590
rect -630 490 -510 590
rect 590 490 710 590
rect 1820 480 1940 580
rect 3030 490 3150 590
<< metal1 >>
rect 2338 9110 2442 9116
rect -2612 9100 -2498 9106
rect -2612 9030 -2600 9100
rect -2510 9030 -2498 9100
rect -2612 9024 -2498 9030
rect -2442 9100 -2328 9106
rect -2442 9030 -2430 9100
rect -2340 9030 -2328 9100
rect -2442 9024 -2328 9030
rect -122 9100 -8 9106
rect -122 9030 -110 9100
rect -20 9030 -8 9100
rect -122 9024 -8 9030
rect 48 9100 162 9106
rect 48 9030 60 9100
rect 150 9030 162 9100
rect 48 9024 162 9030
rect 2338 9030 2350 9110
rect 2430 9030 2442 9110
rect 2338 9024 2442 9030
rect 2508 9110 2612 9116
rect 2508 9030 2520 9110
rect 2600 9030 2612 9110
rect 2508 9024 2612 9030
rect -2610 8940 -2600 8990
rect -4210 8910 -2600 8940
rect -2520 8940 -2510 8990
rect -2440 8940 -2430 8990
rect -2520 8910 -2430 8940
rect -2350 8940 -2340 8990
rect -120 8940 -110 8990
rect -2350 8910 -110 8940
rect -30 8940 -20 8990
rect 50 8940 60 8990
rect -30 8910 60 8940
rect 140 8940 150 8990
rect 2340 8940 2350 8980
rect 140 8910 2350 8940
rect -4210 8900 2350 8910
rect 2430 8940 2440 8980
rect 2510 8940 2520 8980
rect 2430 8900 2520 8940
rect 2600 8940 2610 8980
rect 2600 8900 4230 8940
rect -3160 8850 -3150 8860
rect -4280 8820 -3150 8850
rect -4280 8810 -3480 8820
rect -4300 8750 -3480 8810
rect -4300 8710 -3870 8750
rect -3880 8670 -3870 8710
rect -3790 8710 -3700 8750
rect -3790 8670 -3780 8710
rect -3710 8670 -3700 8710
rect -3620 8740 -3480 8750
rect -3400 8740 -3330 8820
rect -3250 8790 -3150 8820
rect -3020 8850 -3010 8860
rect -1920 8850 -1910 8860
rect -3020 8790 -1910 8850
rect -1780 8850 -1770 8860
rect -690 8850 -680 8860
rect -1780 8820 -680 8850
rect -1780 8790 -990 8820
rect -3250 8750 -990 8790
rect -3250 8740 -1350 8750
rect -3620 8710 -1350 8740
rect -3620 8670 -3610 8710
rect -1360 8670 -1350 8710
rect -1270 8710 -1180 8750
rect -1270 8670 -1260 8710
rect -1190 8670 -1180 8710
rect -1100 8740 -990 8750
rect -910 8740 -840 8820
rect -760 8790 -680 8820
rect -550 8850 -540 8860
rect 550 8850 560 8860
rect -550 8790 560 8850
rect 690 8850 700 8860
rect 1790 8850 1800 8860
rect 690 8820 1800 8850
rect 690 8790 1490 8820
rect -760 8750 1490 8790
rect -760 8740 1140 8750
rect -1100 8710 1140 8740
rect -1100 8670 -1090 8710
rect 1130 8670 1140 8710
rect 1220 8710 1310 8750
rect 1220 8670 1230 8710
rect 1300 8670 1310 8710
rect 1390 8740 1490 8750
rect 1570 8740 1640 8820
rect 1720 8790 1800 8820
rect 1930 8850 1940 8860
rect 3020 8850 3030 8860
rect 1930 8790 3030 8850
rect 3160 8850 3170 8860
rect 3160 8810 4300 8850
rect 3160 8790 4310 8810
rect 1720 8750 4310 8790
rect 1720 8740 3590 8750
rect 1390 8710 3590 8740
rect 1390 8670 1400 8710
rect 3580 8670 3590 8710
rect 3670 8710 3760 8750
rect 3670 8670 3680 8710
rect 3750 8670 3760 8710
rect 3840 8710 4310 8750
rect 3840 8670 3850 8710
rect -2610 8400 -2600 8450
rect -4210 8370 -2600 8400
rect -2520 8400 -2510 8450
rect -2440 8400 -2430 8450
rect -2520 8370 -2430 8400
rect -2350 8400 -2340 8450
rect -120 8400 -110 8450
rect -2350 8370 -110 8400
rect -30 8400 -20 8450
rect 50 8400 60 8450
rect -30 8370 60 8400
rect 140 8400 150 8450
rect 2340 8400 2350 8440
rect 140 8370 2350 8400
rect -4210 8360 2350 8370
rect 2430 8400 2440 8440
rect 2510 8400 2520 8440
rect 2430 8360 2520 8400
rect 2600 8400 2610 8440
rect 2600 8360 4230 8400
rect -3160 8310 -3150 8320
rect -4280 8280 -3150 8310
rect -4280 8270 -3480 8280
rect -4290 8210 -3480 8270
rect -4290 8170 -3870 8210
rect -3880 8130 -3870 8170
rect -3790 8170 -3700 8210
rect -3790 8130 -3780 8170
rect -3710 8130 -3700 8170
rect -3620 8200 -3480 8210
rect -3400 8200 -3330 8280
rect -3250 8250 -3150 8280
rect -3020 8310 -3010 8320
rect -1920 8310 -1910 8320
rect -3020 8250 -1910 8310
rect -1780 8310 -1770 8320
rect -690 8310 -680 8320
rect -1780 8280 -680 8310
rect -1780 8250 -990 8280
rect -3250 8210 -990 8250
rect -3250 8200 -1350 8210
rect -3620 8170 -1350 8200
rect -3620 8130 -3610 8170
rect -1360 8130 -1350 8170
rect -1270 8170 -1180 8210
rect -1270 8130 -1260 8170
rect -1190 8130 -1180 8170
rect -1100 8200 -990 8210
rect -910 8200 -840 8280
rect -760 8250 -680 8280
rect -550 8310 -540 8320
rect 550 8310 560 8320
rect -550 8250 560 8310
rect 690 8310 700 8320
rect 1790 8310 1800 8320
rect 690 8280 1800 8310
rect 690 8250 1490 8280
rect -760 8210 1490 8250
rect -760 8200 1140 8210
rect -1100 8170 1140 8200
rect -1100 8130 -1090 8170
rect 1130 8130 1140 8170
rect 1220 8170 1310 8210
rect 1220 8130 1230 8170
rect 1300 8130 1310 8170
rect 1390 8200 1490 8210
rect 1570 8200 1640 8280
rect 1720 8250 1800 8280
rect 1930 8310 1940 8320
rect 3020 8310 3030 8320
rect 1930 8250 3030 8310
rect 3160 8310 3170 8320
rect 3160 8260 4300 8310
rect 3160 8250 4290 8260
rect 1720 8200 4290 8250
rect 1390 8170 3590 8200
rect 1390 8130 1400 8170
rect 3580 8120 3590 8170
rect 3670 8170 3760 8200
rect 3670 8120 3680 8170
rect 3750 8120 3760 8170
rect 3840 8170 4290 8200
rect 3840 8120 3850 8170
rect -2600 8056 -2340 8090
rect 38 8060 152 8066
rect -2602 8050 -2340 8056
rect -2602 7980 -2590 8050
rect -2500 7980 -2450 8050
rect -2360 7980 -2340 8050
rect -2602 7974 -2340 7980
rect -122 8050 -8 8056
rect -122 7980 -110 8050
rect -20 7980 -8 8050
rect 38 7990 50 8060
rect 140 7990 152 8060
rect 38 7984 152 7990
rect 2338 8060 2442 8066
rect 2338 7990 2350 8060
rect 2430 7990 2442 8060
rect 2338 7984 2442 7990
rect 2508 8060 2612 8066
rect 2508 7990 2520 8060
rect 2600 7990 2612 8060
rect 2508 7984 2612 7990
rect -122 7974 -8 7980
rect -2600 7940 -2340 7974
rect -2610 7860 -2600 7910
rect -4210 7830 -2600 7860
rect -2520 7860 -2510 7910
rect -2440 7860 -2430 7910
rect -2520 7830 -2430 7860
rect -2350 7860 -2340 7910
rect -120 7860 -110 7920
rect -2350 7840 -110 7860
rect -30 7860 -20 7920
rect 50 7860 60 7920
rect -30 7840 60 7860
rect 140 7860 150 7920
rect 2340 7860 2350 7900
rect 140 7840 2350 7860
rect -2350 7830 2350 7840
rect -4210 7820 2350 7830
rect 2430 7860 2440 7900
rect 2510 7860 2520 7900
rect 2430 7820 2520 7860
rect 2600 7860 2610 7900
rect 2600 7820 4230 7860
rect -3160 7770 -3150 7780
rect -4280 7740 -3150 7770
rect -4280 7670 -3480 7740
rect -4280 7630 -3870 7670
rect -3880 7590 -3870 7630
rect -3790 7630 -3700 7670
rect -3790 7590 -3780 7630
rect -3710 7590 -3700 7630
rect -3620 7660 -3480 7670
rect -3400 7660 -3330 7740
rect -3250 7710 -3150 7740
rect -3020 7770 -3010 7780
rect -1920 7770 -1910 7780
rect -3020 7710 -1910 7770
rect -1780 7770 -1770 7780
rect -690 7770 -680 7780
rect -1780 7740 -680 7770
rect -1780 7710 -990 7740
rect -3250 7670 -990 7710
rect -3250 7660 -1350 7670
rect -3620 7630 -1350 7660
rect -3620 7590 -3610 7630
rect -1360 7590 -1350 7630
rect -1270 7630 -1180 7670
rect -1270 7590 -1260 7630
rect -1190 7590 -1180 7630
rect -1100 7660 -990 7670
rect -910 7660 -840 7740
rect -760 7710 -680 7740
rect -550 7770 -540 7780
rect 550 7770 560 7780
rect -550 7710 560 7770
rect 690 7770 700 7780
rect 1790 7770 1800 7780
rect 690 7740 1800 7770
rect 690 7710 1500 7740
rect -760 7660 1500 7710
rect 1580 7660 1640 7740
rect 1720 7710 1800 7740
rect 1930 7770 1940 7780
rect 3020 7770 3030 7780
rect 1930 7710 3030 7770
rect 3160 7770 3170 7780
rect 3160 7710 4300 7770
rect 1720 7670 4300 7710
rect 1720 7660 3590 7670
rect -1100 7630 1140 7660
rect -1100 7590 -1090 7630
rect 1130 7580 1140 7630
rect 1220 7630 1310 7660
rect 1220 7580 1230 7630
rect 1300 7580 1310 7630
rect 1390 7630 3590 7660
rect 1390 7580 1400 7630
rect 3580 7590 3590 7630
rect 3670 7630 3760 7670
rect 3670 7590 3680 7630
rect 3750 7590 3760 7630
rect 3840 7630 4300 7670
rect 3840 7590 3850 7630
rect -2602 7520 -2498 7526
rect -2602 7440 -2590 7520
rect -2510 7440 -2498 7520
rect -2602 7434 -2498 7440
rect -2432 7520 -2328 7526
rect -2432 7440 -2420 7520
rect -2340 7440 -2328 7520
rect -2432 7434 -2328 7440
rect -122 7520 -18 7526
rect -122 7440 -110 7520
rect -30 7440 -18 7520
rect -122 7434 -18 7440
rect 48 7520 152 7526
rect 48 7440 60 7520
rect 140 7440 152 7520
rect 48 7434 152 7440
rect 2338 7520 2442 7526
rect 2338 7440 2350 7520
rect 2430 7440 2442 7520
rect 2338 7434 2442 7440
rect 2508 7520 2612 7526
rect 2508 7440 2520 7520
rect 2600 7440 2612 7520
rect 2508 7434 2612 7440
rect -2600 7330 -2590 7390
rect -4200 7310 -2590 7330
rect -2510 7330 -2500 7390
rect -2430 7330 -2420 7390
rect -2510 7310 -2420 7330
rect -2340 7330 -2330 7390
rect -120 7330 -110 7400
rect -2340 7320 -110 7330
rect -30 7330 -20 7400
rect 50 7330 60 7400
rect -30 7320 60 7330
rect 140 7330 150 7400
rect 2340 7330 2350 7390
rect 140 7320 2350 7330
rect -2340 7310 2350 7320
rect 2430 7330 2440 7390
rect 2510 7330 2520 7390
rect 2430 7310 2520 7330
rect 2600 7330 2610 7390
rect 2600 7310 4240 7330
rect -4200 7290 4240 7310
rect -3160 7230 -3150 7240
rect -4280 7180 -3150 7230
rect -3160 7170 -3150 7180
rect -3020 7230 -3010 7240
rect -1920 7230 -1910 7240
rect -3020 7180 -1910 7230
rect -3020 7170 -3010 7180
rect -1920 7170 -1910 7180
rect -1780 7230 -1770 7240
rect -690 7230 -680 7240
rect -1780 7180 -680 7230
rect -1780 7170 -1770 7180
rect -690 7170 -680 7180
rect -550 7230 -540 7240
rect 550 7230 560 7240
rect -550 7180 560 7230
rect -550 7170 -540 7180
rect 550 7170 560 7180
rect 690 7230 700 7240
rect 1780 7230 1790 7240
rect 690 7180 1790 7230
rect 690 7170 700 7180
rect 1780 7170 1790 7180
rect 1920 7230 1930 7240
rect 3020 7230 3030 7240
rect 1920 7180 3030 7230
rect 1920 7170 1930 7180
rect 3020 7170 3030 7180
rect 3160 7230 3170 7240
rect 3160 7180 4300 7230
rect 3160 7170 3170 7180
rect 200 7140 430 7150
rect -2200 7130 -2190 7140
rect -4210 7090 -3870 7130
rect -3880 7050 -3870 7090
rect -3790 7090 -3700 7130
rect -3790 7050 -3780 7090
rect -3710 7050 -3700 7090
rect -3620 7090 -2190 7130
rect -3620 7050 -3610 7090
rect -2210 7060 -2190 7090
rect -2110 7130 -2100 7140
rect -2090 7130 -2080 7140
rect -2110 7060 -2080 7130
rect -2000 7130 -1990 7140
rect 200 7130 220 7140
rect -2000 7090 -1360 7130
rect -2000 7060 -1980 7090
rect -2210 7030 -1980 7060
rect -1370 7050 -1360 7090
rect -1280 7090 -1190 7130
rect -1280 7050 -1270 7090
rect -1200 7050 -1190 7090
rect -1110 7090 220 7130
rect -1110 7050 -1100 7090
rect 200 7060 220 7090
rect 300 7060 330 7140
rect 410 7130 430 7140
rect 2660 7130 2890 7140
rect 410 7090 1130 7130
rect 410 7060 430 7090
rect 200 7050 430 7060
rect 1120 7050 1130 7090
rect 1210 7090 1300 7130
rect 1210 7050 1220 7090
rect 1290 7050 1300 7090
rect 1380 7090 2680 7130
rect 1380 7050 1390 7090
rect 2660 7050 2680 7090
rect 2760 7050 2790 7130
rect 2870 7090 3620 7130
rect 2870 7050 2890 7090
rect 3610 7050 3620 7090
rect 3700 7090 3790 7130
rect 3700 7050 3710 7090
rect 3780 7050 3790 7090
rect 3870 7090 4230 7130
rect 3870 7050 3880 7090
rect 2660 7030 2890 7050
rect -2600 6750 -2590 6810
rect -4210 6730 -2590 6750
rect -2510 6750 -2500 6810
rect -2430 6750 -2420 6810
rect -2510 6730 -2420 6750
rect -2340 6750 -2330 6810
rect -120 6750 -110 6820
rect -2340 6740 -110 6750
rect -30 6750 -20 6820
rect 50 6750 60 6820
rect -30 6740 60 6750
rect 140 6750 150 6820
rect 2340 6750 2350 6810
rect 140 6740 2350 6750
rect -2340 6730 2350 6740
rect 2430 6750 2440 6810
rect 2510 6750 2520 6810
rect 2430 6730 2520 6750
rect 2600 6750 2610 6810
rect 2600 6730 4230 6750
rect -4210 6710 4230 6730
rect -3160 6650 -3150 6660
rect -4280 6600 -3150 6650
rect -3160 6590 -3150 6600
rect -3020 6650 -3010 6660
rect -1920 6650 -1910 6660
rect -3020 6600 -1910 6650
rect -3020 6590 -3010 6600
rect -1920 6590 -1910 6600
rect -1780 6650 -1770 6660
rect -680 6650 -670 6660
rect -1780 6600 -670 6650
rect -1780 6590 -1770 6600
rect -680 6590 -670 6600
rect -540 6650 -530 6660
rect 550 6650 560 6660
rect -540 6600 560 6650
rect -540 6590 -530 6600
rect 550 6590 560 6600
rect 690 6650 700 6660
rect 1780 6650 1790 6660
rect 690 6600 1790 6650
rect 690 6590 700 6600
rect 1780 6590 1790 6600
rect 1920 6650 1930 6660
rect 3020 6650 3030 6660
rect 1920 6600 3030 6650
rect 1920 6590 1930 6600
rect 3020 6590 3030 6600
rect 3160 6650 3170 6660
rect 3160 6600 4300 6650
rect 3160 6590 3170 6600
rect 200 6550 430 6560
rect 2660 6550 2890 6560
rect -4210 6510 -3870 6550
rect -3880 6470 -3870 6510
rect -3790 6510 -3700 6550
rect -3790 6470 -3780 6510
rect -3710 6470 -3700 6510
rect -3620 6530 -1360 6550
rect -3620 6510 -2190 6530
rect -3620 6470 -3610 6510
rect -2210 6450 -2190 6510
rect -2110 6450 -2080 6530
rect -2000 6510 -1360 6530
rect -2000 6450 -1980 6510
rect -1370 6470 -1360 6510
rect -1280 6510 -1190 6550
rect -1280 6470 -1270 6510
rect -1200 6470 -1190 6510
rect -1110 6510 220 6550
rect -1110 6470 -1100 6510
rect 200 6470 220 6510
rect 300 6470 330 6550
rect 410 6540 2680 6550
rect 410 6510 1130 6540
rect 410 6470 430 6510
rect 200 6450 430 6470
rect 1120 6460 1130 6510
rect 1210 6510 1300 6540
rect 1210 6460 1220 6510
rect 1290 6460 1300 6510
rect 1380 6510 2680 6540
rect 1380 6460 1390 6510
rect 2660 6470 2680 6510
rect 2760 6470 2790 6550
rect 2870 6510 3620 6550
rect 2870 6470 2890 6510
rect 3610 6470 3620 6510
rect 3700 6510 3790 6550
rect 3700 6470 3710 6510
rect 3780 6470 3790 6510
rect 3870 6510 4230 6550
rect 3870 6470 3880 6510
rect 2660 6450 2890 6470
rect -2210 6440 -1980 6450
rect 9540 6440 9970 6560
rect -9960 6270 -9530 6390
rect -2602 6360 -2488 6366
rect -2602 6280 -2590 6360
rect -2500 6280 -2488 6360
rect -2602 6274 -2488 6280
rect -2442 6360 -2328 6366
rect -2442 6280 -2430 6360
rect -2340 6280 -2328 6360
rect -2442 6274 -2328 6280
rect -122 6350 -18 6356
rect -122 6280 -110 6350
rect -30 6280 -18 6350
rect -122 6274 -18 6280
rect 48 6350 152 6356
rect 48 6280 60 6350
rect 140 6280 152 6350
rect 48 6274 152 6280
rect 2338 6350 2442 6356
rect 2338 6280 2350 6350
rect 2430 6280 2442 6350
rect 2338 6274 2442 6280
rect 2508 6350 2612 6356
rect 2508 6280 2520 6350
rect 2600 6280 2612 6350
rect 2508 6274 2612 6280
rect 9540 6300 9560 6440
rect 9690 6300 9820 6440
rect 9950 6300 9970 6440
rect -9960 6130 -9940 6270
rect -9810 6130 -9690 6270
rect -9560 6130 -9530 6270
rect -2600 6170 -2590 6230
rect -4210 6150 -2590 6170
rect -2510 6170 -2500 6230
rect -2430 6170 -2420 6230
rect -2510 6150 -2420 6170
rect -2340 6170 -2330 6230
rect -120 6170 -110 6240
rect -2340 6160 -110 6170
rect -30 6170 -20 6240
rect 50 6170 60 6240
rect -30 6160 60 6170
rect 140 6170 150 6240
rect 2340 6170 2350 6230
rect 140 6160 2350 6170
rect -2340 6150 2350 6160
rect 2430 6170 2440 6230
rect 2510 6170 2520 6230
rect 2430 6150 2520 6170
rect 2600 6170 2610 6230
rect 2600 6150 4230 6170
rect -4210 6130 4230 6150
rect -9960 3530 -9530 6130
rect -3160 6070 -3150 6080
rect -4280 6020 -3150 6070
rect -3160 6010 -3150 6020
rect -3020 6070 -3010 6080
rect -1920 6070 -1910 6080
rect -3020 6020 -1910 6070
rect -3020 6010 -3010 6020
rect -1920 6010 -1910 6020
rect -1780 6070 -1770 6080
rect -690 6070 -680 6080
rect -1780 6020 -680 6070
rect -1780 6010 -1770 6020
rect -690 6010 -680 6020
rect -550 6070 -540 6080
rect 550 6070 560 6080
rect -550 6020 560 6070
rect -550 6010 -540 6020
rect 550 6010 560 6020
rect 690 6070 700 6080
rect 1780 6070 1790 6080
rect 690 6020 1790 6070
rect 690 6010 700 6020
rect 1780 6010 1790 6020
rect 1920 6070 1930 6080
rect 3020 6070 3030 6080
rect 1920 6020 3030 6070
rect 1920 6010 1930 6020
rect 3020 6010 3030 6020
rect 3160 6070 3170 6080
rect 3160 6020 4300 6070
rect 3160 6010 3170 6020
rect -7530 5560 -7100 6000
rect -2210 5960 -1980 5990
rect 200 5970 430 5980
rect 2660 5970 2890 5980
rect -1370 5960 -1360 5970
rect -4210 5940 -1360 5960
rect -4210 5920 -3890 5940
rect -3900 5860 -3890 5920
rect -3810 5920 -3680 5940
rect -3810 5860 -3800 5920
rect -3690 5860 -3680 5920
rect -3600 5920 -1360 5940
rect -3600 5860 -3590 5920
rect -2210 5870 -1980 5920
rect -1370 5890 -1360 5920
rect -1280 5960 -1270 5970
rect -1200 5960 -1190 5970
rect -1280 5920 -1190 5960
rect -1280 5890 -1270 5920
rect -1200 5890 -1190 5920
rect -1110 5960 -1100 5970
rect 200 5960 220 5970
rect -1110 5920 220 5960
rect -1110 5890 -1100 5920
rect 200 5890 220 5920
rect 300 5890 330 5970
rect 410 5960 430 5970
rect 1120 5960 1130 5970
rect 410 5920 1130 5960
rect 410 5890 430 5920
rect 1120 5890 1130 5920
rect 1210 5960 1220 5970
rect 1290 5960 1300 5970
rect 1210 5920 1300 5960
rect 1210 5890 1220 5920
rect 1290 5890 1300 5920
rect 1380 5960 1390 5970
rect 2660 5960 2680 5970
rect 1380 5920 2680 5960
rect 1380 5890 1390 5920
rect 2660 5890 2680 5920
rect 2760 5890 2790 5970
rect 2870 5960 2890 5970
rect 3610 5960 3620 5970
rect 2870 5920 3620 5960
rect 2870 5890 2890 5920
rect 3610 5890 3620 5920
rect 3700 5960 3710 5970
rect 3780 5960 3790 5970
rect 3700 5920 3790 5960
rect 3700 5890 3710 5920
rect 3780 5890 3790 5920
rect 3870 5960 3880 5970
rect 3870 5920 4230 5960
rect 3870 5890 3880 5920
rect 200 5870 430 5890
rect 2660 5870 2890 5890
rect -4480 5630 -4470 5700
rect -6050 5620 -4470 5630
rect -4390 5630 -4380 5700
rect -4250 5630 -4240 5700
rect -4390 5620 -4240 5630
rect -4160 5630 -4150 5700
rect -1930 5630 -1920 5690
rect -4160 5620 -1920 5630
rect -6050 5610 -1920 5620
rect -1840 5630 -1830 5690
rect -1760 5630 -1750 5690
rect -1840 5610 -1750 5630
rect -1670 5630 -1660 5690
rect 530 5630 540 5690
rect -1670 5610 540 5630
rect 620 5630 630 5690
rect 720 5630 730 5690
rect 620 5610 730 5630
rect 810 5630 820 5690
rect 2980 5630 2990 5690
rect 810 5610 2990 5630
rect 3070 5630 3080 5690
rect 3170 5630 3180 5690
rect 3070 5610 3180 5630
rect 3260 5630 3270 5690
rect 5490 5630 5500 5690
rect 3260 5610 5500 5630
rect 5580 5630 5590 5690
rect 5660 5630 5670 5690
rect 5580 5610 5670 5630
rect 5750 5630 5760 5690
rect 5750 5610 6100 5630
rect -6050 5580 6100 5610
rect 7100 5560 7530 6000
rect -7530 5530 -6090 5560
rect -5000 5530 -4990 5540
rect -7530 5490 -4990 5530
rect -7530 5460 -6090 5490
rect -5000 5470 -4990 5490
rect -4860 5530 -4850 5540
rect -3760 5530 -3750 5540
rect -4860 5490 -3750 5530
rect -4860 5470 -4850 5490
rect -3760 5470 -3750 5490
rect -3620 5530 -3610 5540
rect -2530 5530 -2520 5540
rect -3620 5490 -2520 5530
rect -3620 5470 -3610 5490
rect -2530 5470 -2520 5490
rect -2390 5530 -2380 5540
rect -1290 5530 -1280 5540
rect -2390 5490 -1280 5530
rect -2390 5470 -2380 5490
rect -1290 5470 -1280 5490
rect -1150 5530 -1140 5540
rect -50 5530 -40 5540
rect -1150 5490 -40 5530
rect -1150 5470 -1140 5490
rect -50 5470 -40 5490
rect 90 5530 100 5540
rect 1180 5530 1190 5540
rect 90 5490 1190 5530
rect 90 5470 100 5490
rect 1180 5470 1190 5490
rect 1320 5530 1330 5540
rect 2420 5530 2430 5540
rect 1320 5490 2430 5530
rect 1320 5470 1330 5490
rect 2420 5470 2430 5490
rect 2560 5530 2570 5540
rect 3650 5530 3660 5540
rect 2560 5490 3660 5530
rect 2560 5470 2570 5490
rect 3650 5470 3660 5490
rect 3790 5530 3800 5540
rect 4890 5530 4900 5540
rect 3790 5490 4900 5530
rect 3790 5470 3800 5490
rect 4890 5470 4900 5490
rect 5030 5530 5040 5540
rect 6130 5530 7530 5560
rect 5030 5490 7530 5530
rect 5030 5470 5040 5490
rect 6130 5460 7530 5490
rect -7530 5020 -7100 5460
rect -6050 5420 6100 5430
rect -6050 5380 -5720 5420
rect -5730 5340 -5720 5380
rect -5640 5380 -5510 5420
rect -5640 5340 -5630 5380
rect -5520 5340 -5510 5380
rect -5430 5380 -3240 5420
rect -5430 5340 -5420 5380
rect -3250 5340 -3240 5380
rect -3160 5380 -3020 5420
rect -3160 5340 -3150 5380
rect -3030 5340 -3020 5380
rect -2940 5380 -710 5420
rect -2940 5340 -2930 5380
rect -720 5340 -710 5380
rect -630 5380 -530 5420
rect -630 5340 -620 5380
rect -540 5340 -530 5380
rect -450 5410 6100 5420
rect -450 5380 1750 5410
rect -450 5340 -440 5380
rect 1740 5330 1750 5380
rect 1830 5380 1930 5410
rect 1830 5330 1840 5380
rect 1920 5330 1930 5380
rect 2010 5380 4230 5410
rect 2010 5330 2020 5380
rect 4220 5330 4230 5380
rect 4310 5380 4400 5410
rect 4310 5330 4320 5380
rect 4390 5330 4400 5380
rect 4480 5380 6100 5410
rect 4480 5330 4490 5380
rect -4462 5280 -4348 5286
rect -4462 5200 -4450 5280
rect -4360 5200 -4348 5280
rect -4462 5194 -4348 5200
rect -4282 5280 -4168 5286
rect -4282 5200 -4270 5280
rect -4180 5200 -4168 5280
rect -4282 5194 -4168 5200
rect -1932 5280 -1818 5286
rect -1932 5200 -1920 5280
rect -1830 5200 -1818 5280
rect -1932 5194 -1818 5200
rect -1772 5280 -1658 5286
rect -1772 5200 -1760 5280
rect -1670 5200 -1658 5280
rect -1772 5194 -1658 5200
rect 538 5280 652 5286
rect 538 5200 550 5280
rect 640 5200 652 5280
rect 538 5194 652 5200
rect 698 5280 812 5286
rect 698 5200 710 5280
rect 800 5200 812 5280
rect 698 5194 812 5200
rect 2988 5280 3102 5286
rect 2988 5200 3000 5280
rect 3090 5200 3102 5280
rect 2988 5194 3102 5200
rect 3148 5280 3262 5286
rect 3148 5200 3160 5280
rect 3250 5200 3262 5280
rect 3148 5194 3262 5200
rect 5488 5280 5602 5286
rect 5488 5200 5500 5280
rect 5590 5200 5602 5280
rect 5488 5194 5602 5200
rect 5648 5280 5762 5286
rect 5648 5200 5660 5280
rect 5750 5200 5762 5280
rect 5648 5194 5762 5200
rect -4480 5100 -4470 5160
rect -6050 5080 -4470 5100
rect -4390 5100 -4380 5160
rect -4250 5100 -4240 5160
rect -4390 5080 -4240 5100
rect -4160 5100 -4150 5160
rect -1930 5100 -1920 5150
rect -4160 5080 -1920 5100
rect -6050 5070 -1920 5080
rect -1840 5100 -1830 5150
rect -1760 5100 -1750 5160
rect -1840 5080 -1750 5100
rect -1670 5100 -1660 5160
rect 530 5100 540 5160
rect -1670 5080 540 5100
rect 620 5100 630 5160
rect 720 5100 730 5160
rect 620 5080 730 5100
rect 810 5100 820 5160
rect 2980 5100 2990 5150
rect 810 5080 2990 5100
rect -1840 5070 2990 5080
rect 3070 5100 3080 5150
rect 3170 5100 3180 5150
rect 3070 5070 3180 5100
rect 3260 5100 3270 5150
rect 5490 5100 5500 5150
rect 3260 5070 5500 5100
rect 5580 5100 5590 5150
rect 5660 5100 5670 5150
rect 5580 5070 5670 5100
rect 5750 5100 5760 5150
rect 5750 5070 6100 5100
rect -6050 5050 6100 5070
rect -7530 4990 -6090 5020
rect 7100 5010 7530 5460
rect -5000 4990 -4990 5010
rect -7530 4950 -4990 4990
rect -7530 4910 -6090 4950
rect -5000 4940 -4990 4950
rect -4860 4990 -4850 5010
rect -3760 4990 -3750 5000
rect -4860 4950 -3750 4990
rect -4860 4940 -4850 4950
rect -3760 4930 -3750 4950
rect -3620 4990 -3610 5000
rect -2530 4990 -2520 5000
rect -3620 4950 -2520 4990
rect -3620 4930 -3610 4950
rect -2530 4930 -2520 4950
rect -2390 4990 -2380 5000
rect -1290 4990 -1280 5000
rect -2390 4950 -1280 4990
rect -2390 4930 -2380 4950
rect -1290 4930 -1280 4950
rect -1150 4990 -1140 5000
rect -50 4990 -40 5000
rect -1150 4950 -40 4990
rect -1150 4930 -1140 4950
rect -50 4930 -40 4950
rect 90 4990 100 5000
rect 1180 4990 1190 5000
rect 90 4950 1190 4990
rect 90 4930 100 4950
rect 1180 4930 1190 4950
rect 1320 4990 1330 5000
rect 2420 4990 2430 5000
rect 1320 4950 2430 4990
rect 1320 4930 1330 4950
rect 2420 4930 2430 4950
rect 2560 4990 2570 5000
rect 3650 4990 3660 5000
rect 2560 4950 3660 4990
rect 2560 4930 2570 4950
rect 3650 4930 3660 4950
rect 3790 4990 3800 5000
rect 4890 4990 4900 5000
rect 3790 4950 4900 4990
rect 3790 4930 3800 4950
rect 4890 4930 4900 4950
rect 5030 4990 5040 5000
rect 6130 4990 7530 5010
rect 5030 4950 7530 4990
rect 5030 4930 5040 4950
rect 6130 4910 7530 4950
rect -7530 4480 -7100 4910
rect -6050 4880 6100 4890
rect -6050 4840 -5720 4880
rect -5730 4800 -5720 4840
rect -5640 4840 -5510 4880
rect -5640 4800 -5630 4840
rect -5520 4800 -5510 4840
rect -5430 4840 -3240 4880
rect -5430 4800 -5420 4840
rect -3250 4800 -3240 4840
rect -3160 4840 -3020 4880
rect -3160 4800 -3150 4840
rect -3030 4800 -3020 4840
rect -2940 4840 -710 4880
rect -2940 4800 -2930 4840
rect -720 4800 -710 4840
rect -630 4840 -520 4880
rect -630 4800 -620 4840
rect -530 4800 -520 4840
rect -440 4870 6100 4880
rect -440 4840 1750 4870
rect -440 4800 -430 4840
rect 1740 4790 1750 4840
rect 1830 4840 1930 4870
rect 1830 4790 1840 4840
rect 1920 4790 1930 4840
rect 2010 4840 4230 4870
rect 2010 4790 2020 4840
rect 4220 4790 4230 4840
rect 4310 4840 4400 4870
rect 4310 4790 4320 4840
rect 4390 4790 4400 4840
rect 4480 4840 6100 4870
rect 4480 4790 4490 4840
rect -4480 4560 -4470 4620
rect -6050 4540 -4470 4560
rect -4390 4560 -4380 4620
rect -4250 4560 -4240 4620
rect -4390 4540 -4240 4560
rect -4160 4560 -4150 4620
rect -1940 4560 -1930 4610
rect -4160 4540 -1930 4560
rect -6050 4530 -1930 4540
rect -1850 4560 -1840 4610
rect -1770 4560 -1760 4610
rect -1850 4530 -1760 4560
rect -1680 4560 -1670 4610
rect 530 4560 540 4610
rect -1680 4530 540 4560
rect 620 4560 630 4610
rect 710 4560 720 4610
rect 620 4530 720 4560
rect 800 4560 810 4610
rect 2980 4560 2990 4610
rect 800 4530 2990 4560
rect 3070 4560 3080 4610
rect 3170 4560 3180 4610
rect 3070 4530 3180 4560
rect 3260 4560 3270 4610
rect 5490 4560 5500 4610
rect 3260 4530 5500 4560
rect 5580 4560 5590 4610
rect 5660 4560 5670 4610
rect 5580 4530 5670 4560
rect 5750 4560 5760 4610
rect 5750 4530 6100 4560
rect -6050 4510 6100 4530
rect 7100 4480 7530 4910
rect -7530 4450 -6070 4480
rect -5000 4450 -4990 4460
rect -7530 4410 -4990 4450
rect -7530 4370 -6070 4410
rect -5000 4390 -4990 4410
rect -4860 4450 -4850 4460
rect -3760 4450 -3750 4460
rect -4860 4410 -3750 4450
rect -4860 4390 -4850 4410
rect -3760 4390 -3750 4410
rect -3620 4450 -3610 4460
rect -2530 4450 -2520 4460
rect -3620 4410 -2520 4450
rect -3620 4390 -3610 4410
rect -2530 4390 -2520 4410
rect -2390 4450 -2380 4460
rect -1290 4450 -1280 4460
rect -2390 4410 -1280 4450
rect -2390 4390 -2380 4410
rect -1290 4390 -1280 4410
rect -1150 4450 -1140 4460
rect -50 4450 -40 4460
rect -1150 4410 -40 4450
rect -1150 4390 -1140 4410
rect -50 4390 -40 4410
rect 90 4450 100 4460
rect 1180 4450 1190 4460
rect 90 4410 1190 4450
rect 90 4390 100 4410
rect 1180 4390 1190 4410
rect 1320 4450 1330 4460
rect 2420 4450 2430 4460
rect 1320 4410 2430 4450
rect 1320 4390 1330 4410
rect 2420 4390 2430 4410
rect 2560 4450 2570 4460
rect 3650 4450 3660 4460
rect 2560 4410 3660 4450
rect 2560 4390 2570 4410
rect 3650 4390 3660 4410
rect 3790 4450 3800 4460
rect 4890 4450 4900 4460
rect 3790 4410 4900 4450
rect 3790 4390 3800 4410
rect 4890 4390 4900 4410
rect 5030 4450 5040 4460
rect 6130 4450 7530 4480
rect 5030 4410 7530 4450
rect 5030 4390 5040 4410
rect 6130 4380 7530 4410
rect -7530 3940 -7100 4370
rect -6050 4340 6100 4350
rect -6050 4300 -5720 4340
rect -5730 4260 -5720 4300
rect -5640 4300 -5510 4340
rect -5640 4260 -5630 4300
rect -5520 4260 -5510 4300
rect -5430 4300 -3250 4340
rect -5430 4260 -5420 4300
rect -3260 4260 -3250 4300
rect -3170 4300 -3010 4340
rect -3170 4260 -3160 4300
rect -3020 4260 -3010 4300
rect -2930 4300 -710 4340
rect -2930 4260 -2920 4300
rect -720 4260 -710 4300
rect -630 4300 -530 4340
rect -630 4260 -620 4300
rect -540 4260 -530 4300
rect -450 4330 6100 4340
rect -450 4300 1760 4330
rect -450 4260 -440 4300
rect 1750 4250 1760 4300
rect 1840 4300 1930 4330
rect 1840 4250 1850 4300
rect 1920 4250 1930 4300
rect 2010 4300 4230 4330
rect 2010 4250 2020 4300
rect 4220 4250 4230 4300
rect 4310 4300 4400 4330
rect 4310 4250 4320 4300
rect 4390 4250 4400 4300
rect 4480 4300 6100 4330
rect 4480 4250 4490 4300
rect -4282 4210 -4168 4216
rect -4462 4200 -4348 4206
rect -4462 4120 -4450 4200
rect -4360 4120 -4348 4200
rect -4282 4130 -4270 4210
rect -4180 4130 -4168 4210
rect -4282 4124 -4168 4130
rect -1932 4200 -1818 4206
rect -4462 4114 -4348 4120
rect -1932 4120 -1920 4200
rect -1830 4120 -1818 4200
rect -1932 4114 -1818 4120
rect -1772 4200 -1658 4206
rect -1772 4120 -1760 4200
rect -1670 4120 -1658 4200
rect -1772 4114 -1658 4120
rect 538 4200 652 4206
rect 538 4120 550 4200
rect 640 4120 652 4200
rect 538 4114 652 4120
rect 698 4200 812 4206
rect 698 4120 710 4200
rect 800 4120 812 4200
rect 698 4114 812 4120
rect 2988 4200 3102 4206
rect 2988 4120 3000 4200
rect 3090 4120 3102 4200
rect 2988 4114 3102 4120
rect 3148 4200 3262 4206
rect 3148 4120 3160 4200
rect 3250 4120 3262 4200
rect 3148 4114 3262 4120
rect 5488 4200 5602 4206
rect 5488 4120 5500 4200
rect 5590 4120 5602 4200
rect 5488 4114 5602 4120
rect 5648 4200 5762 4206
rect 5648 4120 5660 4200
rect 5750 4120 5762 4200
rect 5648 4114 5762 4120
rect -4480 4020 -4470 4070
rect -6050 3990 -4470 4020
rect -4390 4020 -4380 4070
rect -4250 4020 -4240 4070
rect -4390 3990 -4240 4020
rect -4160 4020 -4150 4070
rect -1950 4020 -1940 4080
rect -4160 4000 -1940 4020
rect -1860 4020 -1850 4080
rect -1760 4020 -1750 4080
rect -1860 4000 -1750 4020
rect -1670 4020 -1660 4080
rect 530 4020 540 4070
rect -1670 4000 540 4020
rect -4160 3990 540 4000
rect 620 4020 630 4070
rect 720 4020 730 4070
rect 620 3990 730 4020
rect 810 4020 820 4070
rect 2980 4020 2990 4070
rect 810 3990 2990 4020
rect 3070 4020 3080 4070
rect 3170 4020 3180 4070
rect 3070 3990 3180 4020
rect 3260 4020 3270 4070
rect 5490 4020 5500 4060
rect 3260 3990 5500 4020
rect -6050 3980 5500 3990
rect 5580 4020 5590 4060
rect 5660 4020 5670 4060
rect 5580 3980 5670 4020
rect 5750 4020 5760 4060
rect 5750 3980 6100 4020
rect -6050 3970 6100 3980
rect 7100 3940 7530 4380
rect -7530 3910 -6080 3940
rect -5000 3910 -4990 3920
rect -7530 3870 -4990 3910
rect -7530 3830 -6080 3870
rect -5000 3850 -4990 3870
rect -4860 3910 -4850 3920
rect -3760 3910 -3750 3920
rect -4860 3870 -3750 3910
rect -4860 3850 -4850 3870
rect -3760 3850 -3750 3870
rect -3620 3910 -3610 3920
rect -2530 3910 -2520 3920
rect -3620 3870 -2520 3910
rect -3620 3850 -3610 3870
rect -2530 3850 -2520 3870
rect -2390 3910 -2380 3920
rect -1290 3910 -1280 3920
rect -2390 3870 -1280 3910
rect -2390 3850 -2380 3870
rect -1290 3850 -1280 3870
rect -1150 3910 -1140 3920
rect -50 3910 -40 3920
rect -1150 3870 -40 3910
rect -1150 3850 -1140 3870
rect -50 3850 -40 3870
rect 90 3910 100 3920
rect 1180 3910 1190 3920
rect 90 3870 1190 3910
rect 90 3850 100 3870
rect 1180 3850 1190 3870
rect 1320 3910 1330 3920
rect 2420 3910 2430 3920
rect 1320 3870 2430 3910
rect 1320 3850 1330 3870
rect 2420 3850 2430 3870
rect 2560 3910 2570 3920
rect 3650 3910 3660 3920
rect 2560 3870 3660 3910
rect 2560 3850 2570 3870
rect 3650 3850 3660 3870
rect 3790 3910 3800 3920
rect 4890 3910 4900 3920
rect 3790 3870 4900 3910
rect 3790 3850 3800 3870
rect 4890 3850 4900 3870
rect 5030 3910 5040 3920
rect 6130 3910 7530 3940
rect 5030 3870 7530 3910
rect 5030 3850 5040 3870
rect 6130 3840 7530 3870
rect -7530 3520 -7100 3830
rect -6050 3800 6100 3810
rect -6050 3760 -5720 3800
rect -5730 3720 -5720 3760
rect -5640 3760 -5510 3800
rect -5640 3720 -5630 3760
rect -5520 3720 -5510 3760
rect -5430 3790 -710 3800
rect -5430 3760 -3250 3790
rect -5430 3720 -5420 3760
rect -3260 3710 -3250 3760
rect -3170 3760 -3010 3790
rect -3170 3710 -3160 3760
rect -3020 3710 -3010 3760
rect -2930 3760 -710 3790
rect -2930 3710 -2920 3760
rect -720 3720 -710 3760
rect -630 3760 -520 3800
rect -630 3720 -620 3760
rect -530 3720 -520 3760
rect -440 3790 6100 3800
rect -440 3760 1750 3790
rect -440 3720 -430 3760
rect 1740 3710 1750 3760
rect 1830 3760 1940 3790
rect 1830 3710 1840 3760
rect 1930 3710 1940 3760
rect 2020 3780 6100 3790
rect 2020 3760 4230 3780
rect 2020 3710 2030 3760
rect 4220 3700 4230 3760
rect 4310 3760 4400 3780
rect 4310 3700 4320 3760
rect 4390 3700 4400 3760
rect 4480 3760 6100 3780
rect 4480 3700 4490 3760
rect 7100 3520 7530 3840
rect 9540 3500 9970 6300
rect -8816 3390 -8714 3402
rect -8606 3390 -8504 3402
rect -8820 3260 -8810 3390
rect -8720 3260 -8710 3390
rect -8610 3260 -8600 3390
rect -8510 3260 -8500 3390
rect 8494 3380 8576 3392
rect 8654 3380 8736 3392
rect 8490 3290 8500 3380
rect 8570 3290 8580 3380
rect 8650 3290 8660 3380
rect 8730 3290 8740 3380
rect -2210 3270 -1980 3280
rect -8816 3248 -8714 3260
rect -8606 3248 -8504 3260
rect -3760 3220 -3750 3270
rect -4120 3200 -3750 3220
rect -3620 3220 -3610 3270
rect -2440 3260 -2340 3270
rect -2530 3220 -2520 3260
rect -3620 3200 -2520 3220
rect -4120 3190 -2520 3200
rect -2390 3220 -2340 3260
rect -2210 3220 -2190 3270
rect -2390 3190 -2190 3220
rect -2110 3190 -2080 3270
rect -2000 3220 -1980 3270
rect -20 3260 80 3290
rect 200 3270 430 3290
rect 2660 3280 2890 3290
rect -1290 3220 -1280 3260
rect -2000 3190 -1280 3220
rect -1150 3220 -1140 3260
rect -50 3220 -40 3260
rect -1150 3190 -40 3220
rect 90 3220 100 3260
rect 200 3220 220 3270
rect 90 3190 220 3220
rect 300 3190 330 3270
rect 410 3220 430 3270
rect 1180 3220 1190 3260
rect 410 3190 1190 3220
rect 1320 3220 1330 3260
rect 2410 3220 2430 3280
rect 1320 3210 2430 3220
rect 2560 3220 2570 3280
rect 2660 3220 2680 3280
rect 2560 3210 2680 3220
rect 1320 3200 2680 3210
rect 2760 3200 2790 3280
rect 2870 3220 2890 3280
rect 8494 3278 8576 3290
rect 8654 3278 8736 3290
rect 3650 3220 3660 3260
rect 2870 3200 3660 3220
rect 1320 3190 3660 3200
rect 3790 3220 3800 3260
rect 3790 3190 4210 3220
rect -4120 3180 4210 3190
rect -1860 3130 -1710 3140
rect -640 3130 -490 3140
rect 580 3130 730 3140
rect 1800 3130 1950 3140
rect 3010 3130 3160 3140
rect -4190 3090 4270 3130
rect -1860 3070 -1710 3090
rect -640 3070 -490 3090
rect 580 3070 730 3090
rect 1800 3070 1950 3090
rect 3010 3070 3160 3090
rect -4120 3020 4210 3030
rect -4120 3000 1200 3020
rect -4120 2990 -3810 3000
rect -3820 2920 -3810 2990
rect -3720 2920 -3670 3000
rect -3580 2990 1200 3000
rect -3580 2920 -3570 2990
rect -1230 2940 -1130 2990
rect 1190 2940 1200 2990
rect 1290 2940 1340 3020
rect 1430 2990 4210 3020
rect 1430 2940 1440 2990
rect -3810 2770 -3580 2920
rect -2302 2910 -2168 2916
rect -2302 2800 -2290 2910
rect -2180 2800 -2168 2910
rect -2302 2794 -2168 2800
rect -1442 2910 -1308 2916
rect -1442 2800 -1430 2910
rect -1320 2800 -1308 2910
rect -1442 2794 -1308 2800
rect -232 2910 -98 2916
rect -232 2800 -220 2910
rect -110 2800 -98 2910
rect -232 2794 -98 2800
rect 618 2910 752 2916
rect 618 2800 630 2910
rect 740 2800 752 2910
rect 618 2794 752 2800
rect -3820 2720 -3810 2770
rect -4120 2690 -3810 2720
rect -3720 2690 -3670 2770
rect -3580 2720 -3570 2770
rect -2440 2720 -2340 2770
rect -20 2720 80 2790
rect 1200 2760 1430 2940
rect 3650 2930 3750 2990
rect 2188 2910 2322 2916
rect 2188 2800 2200 2910
rect 2310 2800 2322 2910
rect 2188 2794 2322 2800
rect 3068 2910 3202 2916
rect 3068 2800 3080 2910
rect 3190 2800 3202 2910
rect 3068 2794 3202 2800
rect 1190 2720 1200 2760
rect -3580 2690 1200 2720
rect -4120 2680 1200 2690
rect 1290 2680 1340 2760
rect 1430 2720 1440 2760
rect 2410 2720 2510 2780
rect 1430 2680 4210 2720
rect -1860 2630 -1710 2640
rect -640 2630 -490 2640
rect 580 2630 730 2640
rect 1800 2630 1950 2640
rect 3010 2630 3160 2640
rect -4180 2590 4280 2630
rect -1860 2570 -1710 2590
rect -640 2570 -490 2590
rect 580 2570 730 2590
rect 1800 2570 1950 2590
rect 3010 2570 3160 2590
rect -2530 2530 -2380 2540
rect -4120 2510 -990 2530
rect -4120 2490 -3480 2510
rect -3680 2440 -3580 2490
rect -3490 2430 -3480 2490
rect -3400 2490 -3330 2510
rect -3400 2430 -3390 2490
rect -3340 2430 -3330 2490
rect -3250 2490 -990 2510
rect -3250 2430 -3240 2490
rect -2530 2470 -2380 2490
rect -1290 2460 -1130 2490
rect -1230 2440 -1130 2460
rect -1000 2450 -990 2490
rect -910 2490 -840 2530
rect -910 2450 -900 2490
rect -850 2450 -840 2490
rect -760 2490 1490 2530
rect -760 2450 -750 2490
rect -50 2460 100 2490
rect 1210 2430 1310 2490
rect 1480 2450 1490 2490
rect 1570 2490 1630 2530
rect 1570 2450 1580 2490
rect 1620 2450 1630 2490
rect 1710 2490 4210 2530
rect 1710 2450 1720 2490
rect 2420 2460 2570 2490
rect 3650 2460 3800 2490
rect 3650 2430 3750 2460
rect -3120 2280 -2810 2310
rect -3240 2220 -3030 2280
rect -3560 2200 -3030 2220
rect -2950 2200 -2920 2280
rect -2840 2220 -2810 2280
rect 1820 2270 2040 2280
rect -630 2220 -620 2250
rect -2840 2200 -620 2220
rect -3560 2180 -620 2200
rect -630 2170 -620 2180
rect -540 2220 -530 2250
rect 1820 2220 1830 2270
rect -540 2190 1830 2220
rect 1910 2190 1950 2270
rect 2030 2220 2040 2270
rect 3020 2220 3030 2260
rect 2030 2190 3030 2220
rect -540 2180 3030 2190
rect 3110 2220 3120 2260
rect 3110 2180 3560 2220
rect -540 2170 -530 2180
rect -3640 2100 3600 2120
rect -3640 2020 -1850 2100
rect -1770 2020 560 2100
rect 640 2020 3600 2100
rect -3640 2000 3600 2020
rect -3560 1880 -3110 1920
rect -3120 1840 -3110 1880
rect -3030 1880 1780 1920
rect -3030 1840 -3020 1880
rect 1770 1840 1780 1880
rect 1860 1880 3560 1920
rect 1860 1840 1870 1880
rect -3012 1790 -2878 1796
rect -3012 1700 -3000 1790
rect -2890 1700 -2878 1790
rect -3012 1694 -2878 1700
rect 1898 1790 2032 1796
rect 1898 1700 1910 1790
rect 2020 1700 2032 1790
rect 1898 1694 2032 1700
rect -630 1600 -620 1630
rect -3560 1560 -620 1600
rect -630 1550 -620 1560
rect -540 1600 -530 1630
rect 3020 1600 3030 1640
rect -540 1560 3030 1600
rect 3110 1600 3120 1640
rect 3110 1560 3560 1600
rect -540 1550 -530 1560
rect -3620 1490 3620 1500
rect -3660 1480 3620 1490
rect -3660 1400 -2460 1480
rect -2370 1400 -2340 1480
rect -2250 1400 -1850 1480
rect -1770 1400 -10 1480
rect 80 1400 110 1480
rect 200 1400 560 1480
rect 640 1400 2420 1480
rect 2510 1400 2540 1480
rect 2630 1400 3620 1480
rect -3660 1390 3620 1400
rect -3620 1380 3620 1390
rect -3560 1260 -3110 1300
rect -3120 1220 -3110 1260
rect -3030 1260 1780 1300
rect -3030 1220 -3020 1260
rect 1770 1220 1780 1260
rect 1860 1260 3560 1300
rect 1860 1220 1870 1260
rect -1240 1020 -1230 1050
rect -4120 980 -1230 1020
rect -1240 970 -1230 980
rect -1140 1020 -1130 1050
rect 3640 1020 3650 1070
rect -1140 990 3650 1020
rect 3740 1020 3750 1070
rect 3740 990 4200 1020
rect -1140 980 4200 990
rect -1140 970 -1130 980
rect -4200 880 4280 900
rect -4200 800 -2460 880
rect -2370 800 -2340 880
rect -2250 800 -10 880
rect 80 800 110 880
rect 200 800 2420 880
rect 2510 800 2540 880
rect 2630 800 4280 880
rect -4200 780 4280 800
rect -3820 700 -3810 720
rect -4120 660 -3810 700
rect -3820 640 -3810 660
rect -3720 700 -3710 720
rect -3680 700 -3670 720
rect -3720 660 -3670 700
rect -3720 640 -3710 660
rect -3680 640 -3670 660
rect -3580 700 -3570 720
rect 1190 700 1200 720
rect -3580 660 1200 700
rect -3580 640 -3570 660
rect 1190 640 1200 660
rect 1290 700 1300 720
rect 1330 700 1340 720
rect 1290 660 1340 700
rect 1290 640 1300 660
rect 1330 640 1340 660
rect 1430 700 1440 720
rect 1430 660 4200 700
rect 1430 640 1440 660
rect -3080 590 -2920 600
rect -3080 490 -3060 590
rect -2940 490 -2920 590
rect -3080 420 -2920 490
rect -1860 590 -1700 600
rect -1860 490 -1840 590
rect -1720 490 -1700 590
rect -1860 420 -1700 490
rect -650 590 -490 600
rect 578 590 722 596
rect 3018 590 3162 596
rect -650 490 -630 590
rect -510 490 -490 590
rect -1240 420 -1230 450
rect -4120 380 -1230 420
rect -1240 370 -1230 380
rect -1140 420 -1130 450
rect -650 420 -490 490
rect 570 490 590 590
rect 710 490 730 590
rect 1808 580 1952 586
rect 570 420 730 490
rect 1800 480 1820 580
rect 1940 480 1960 580
rect 1800 420 1960 480
rect 3010 490 3030 590
rect 3150 490 3170 590
rect 3010 420 3170 490
rect 3640 420 3650 470
rect -1140 390 3650 420
rect 3740 420 3750 470
rect 3740 390 4200 420
rect -1140 380 4200 390
rect -1140 370 -1130 380
rect -4180 280 4280 300
rect -4180 200 -2460 280
rect -2370 200 -2340 280
rect -2250 200 -10 280
rect 80 200 110 280
rect 200 200 2420 280
rect 2510 200 2540 280
rect 2630 200 4280 280
rect -4180 180 4280 200
rect 1190 100 1200 120
rect -4120 60 -3810 100
rect -3820 20 -3810 60
rect -3720 60 -3670 100
rect -3720 20 -3710 60
rect -3680 20 -3670 60
rect -3580 60 1200 100
rect -3580 20 -3570 60
rect 1190 40 1200 60
rect 1290 100 1300 120
rect 1330 100 1340 120
rect 1290 60 1340 100
rect 1290 40 1300 60
rect 1330 40 1340 60
rect 1430 100 1440 120
rect 1430 60 4200 100
rect 1430 40 1440 60
<< via1 >>
rect -2600 9030 -2510 9100
rect -2430 9030 -2340 9100
rect -110 9030 -20 9100
rect 60 9030 150 9100
rect 2350 9030 2430 9110
rect 2520 9030 2600 9110
rect -2600 8910 -2520 8990
rect -2430 8910 -2350 8990
rect -110 8910 -30 8990
rect 60 8910 140 8990
rect 2350 8900 2430 8980
rect 2520 8900 2600 8980
rect -3870 8670 -3790 8750
rect -3700 8670 -3620 8750
rect -3480 8740 -3400 8820
rect -3330 8740 -3250 8820
rect -3150 8790 -3020 8860
rect -1910 8790 -1780 8860
rect -1350 8670 -1270 8750
rect -1180 8670 -1100 8750
rect -990 8740 -910 8820
rect -840 8740 -760 8820
rect -680 8790 -550 8860
rect 560 8790 690 8860
rect 1140 8670 1220 8750
rect 1310 8670 1390 8750
rect 1490 8740 1570 8820
rect 1640 8740 1720 8820
rect 1800 8790 1930 8860
rect 3030 8790 3160 8860
rect 3590 8670 3670 8750
rect 3760 8670 3840 8750
rect -2600 8370 -2520 8450
rect -2430 8370 -2350 8450
rect -110 8370 -30 8450
rect 60 8370 140 8450
rect 2350 8360 2430 8440
rect 2520 8360 2600 8440
rect -3870 8130 -3790 8210
rect -3700 8130 -3620 8210
rect -3480 8200 -3400 8280
rect -3330 8200 -3250 8280
rect -3150 8250 -3020 8320
rect -1910 8250 -1780 8320
rect -1350 8130 -1270 8210
rect -1180 8130 -1100 8210
rect -990 8200 -910 8280
rect -840 8200 -760 8280
rect -680 8250 -550 8320
rect 560 8250 690 8320
rect 1140 8130 1220 8210
rect 1310 8130 1390 8210
rect 1490 8200 1570 8280
rect 1640 8200 1720 8280
rect 1800 8250 1930 8320
rect 3030 8250 3160 8320
rect 3590 8120 3670 8200
rect 3760 8120 3840 8200
rect -2590 7980 -2500 8050
rect -2450 7980 -2360 8050
rect -110 7980 -20 8050
rect 50 7990 140 8060
rect 2350 7990 2430 8060
rect 2520 7990 2600 8060
rect -2600 7830 -2520 7910
rect -2430 7830 -2350 7910
rect -110 7840 -30 7920
rect 60 7840 140 7920
rect 2350 7820 2430 7900
rect 2520 7820 2600 7900
rect -3870 7590 -3790 7670
rect -3700 7590 -3620 7670
rect -3480 7660 -3400 7740
rect -3330 7660 -3250 7740
rect -3150 7710 -3020 7780
rect -1910 7710 -1780 7780
rect -1350 7590 -1270 7670
rect -1180 7590 -1100 7670
rect -990 7660 -910 7740
rect -840 7660 -760 7740
rect -680 7710 -550 7780
rect 560 7710 690 7780
rect 1500 7660 1580 7740
rect 1640 7660 1720 7740
rect 1800 7710 1930 7780
rect 3030 7710 3160 7780
rect 1140 7580 1220 7660
rect 1310 7580 1390 7660
rect 3590 7590 3670 7670
rect 3760 7590 3840 7670
rect -2590 7440 -2510 7520
rect -2420 7440 -2340 7520
rect -110 7440 -30 7520
rect 60 7440 140 7520
rect 2350 7440 2430 7520
rect 2520 7440 2600 7520
rect -2590 7310 -2510 7390
rect -2420 7310 -2340 7390
rect -110 7320 -30 7400
rect 60 7320 140 7400
rect 2350 7310 2430 7390
rect 2520 7310 2600 7390
rect -3150 7170 -3020 7240
rect -1910 7170 -1780 7240
rect -680 7170 -550 7240
rect 560 7170 690 7240
rect 1790 7170 1920 7240
rect 3030 7170 3160 7240
rect -3870 7050 -3790 7130
rect -3700 7050 -3620 7130
rect -2190 7060 -2110 7140
rect -2080 7060 -2000 7140
rect -1360 7050 -1280 7130
rect -1190 7050 -1110 7130
rect 220 7060 300 7140
rect 330 7060 410 7140
rect 1130 7050 1210 7130
rect 1300 7050 1380 7130
rect 2680 7050 2760 7130
rect 2790 7050 2870 7130
rect 3620 7050 3700 7130
rect 3790 7050 3870 7130
rect -2590 6730 -2510 6810
rect -2420 6730 -2340 6810
rect -110 6740 -30 6820
rect 60 6740 140 6820
rect 2350 6730 2430 6810
rect 2520 6730 2600 6810
rect -3150 6590 -3020 6660
rect -1910 6590 -1780 6660
rect -670 6590 -540 6660
rect 560 6590 690 6660
rect 1790 6590 1920 6660
rect 3030 6590 3160 6660
rect -3870 6470 -3790 6550
rect -3700 6470 -3620 6550
rect -2190 6450 -2110 6530
rect -2080 6450 -2000 6530
rect -1360 6470 -1280 6550
rect -1190 6470 -1110 6550
rect 220 6470 300 6550
rect 330 6470 410 6550
rect 1130 6460 1210 6540
rect 1300 6460 1380 6540
rect 2680 6470 2760 6550
rect 2790 6470 2870 6550
rect 3620 6470 3700 6550
rect 3790 6470 3870 6550
rect -2590 6280 -2500 6360
rect -2430 6280 -2340 6360
rect -110 6280 -30 6350
rect 60 6280 140 6350
rect 2350 6280 2430 6350
rect 2520 6280 2600 6350
rect 9560 6300 9690 6440
rect 9820 6300 9950 6440
rect -9940 6130 -9810 6270
rect -9690 6130 -9560 6270
rect -2590 6150 -2510 6230
rect -2420 6150 -2340 6230
rect -110 6160 -30 6240
rect 60 6160 140 6240
rect 2350 6150 2430 6230
rect 2520 6150 2600 6230
rect -3150 6010 -3020 6080
rect -1910 6010 -1780 6080
rect -680 6010 -550 6080
rect 560 6010 690 6080
rect 1790 6010 1920 6080
rect 3030 6010 3160 6080
rect -3890 5860 -3810 5940
rect -3680 5860 -3600 5940
rect -1360 5890 -1280 5970
rect -1190 5890 -1110 5970
rect 220 5890 300 5970
rect 330 5890 410 5970
rect 1130 5890 1210 5970
rect 1300 5890 1380 5970
rect 2680 5890 2760 5970
rect 2790 5890 2870 5970
rect 3620 5890 3700 5970
rect 3790 5890 3870 5970
rect -4470 5620 -4390 5700
rect -4240 5620 -4160 5700
rect -1920 5610 -1840 5690
rect -1750 5610 -1670 5690
rect 540 5610 620 5690
rect 730 5610 810 5690
rect 2990 5610 3070 5690
rect 3180 5610 3260 5690
rect 5500 5610 5580 5690
rect 5670 5610 5750 5690
rect -4990 5470 -4860 5540
rect -3750 5470 -3620 5540
rect -2520 5470 -2390 5540
rect -1280 5470 -1150 5540
rect -40 5470 90 5540
rect 1190 5470 1320 5540
rect 2430 5470 2560 5540
rect 3660 5470 3790 5540
rect 4900 5470 5030 5540
rect -5720 5340 -5640 5420
rect -5510 5340 -5430 5420
rect -3240 5340 -3160 5420
rect -3020 5340 -2940 5420
rect -710 5340 -630 5420
rect -530 5340 -450 5420
rect 1750 5330 1830 5410
rect 1930 5330 2010 5410
rect 4230 5330 4310 5410
rect 4400 5330 4480 5410
rect -4450 5200 -4360 5280
rect -4270 5200 -4180 5280
rect -1920 5200 -1830 5280
rect -1760 5200 -1670 5280
rect 550 5200 640 5280
rect 710 5200 800 5280
rect 3000 5200 3090 5280
rect 3160 5200 3250 5280
rect 5500 5200 5590 5280
rect 5660 5200 5750 5280
rect -4470 5080 -4390 5160
rect -4240 5080 -4160 5160
rect -1920 5070 -1840 5150
rect -1750 5080 -1670 5160
rect 540 5080 620 5160
rect 730 5080 810 5160
rect 2990 5070 3070 5150
rect 3180 5070 3260 5150
rect 5500 5070 5580 5150
rect 5670 5070 5750 5150
rect -4990 4940 -4860 5010
rect -3750 4930 -3620 5000
rect -2520 4930 -2390 5000
rect -1280 4930 -1150 5000
rect -40 4930 90 5000
rect 1190 4930 1320 5000
rect 2430 4930 2560 5000
rect 3660 4930 3790 5000
rect 4900 4930 5030 5000
rect -5720 4800 -5640 4880
rect -5510 4800 -5430 4880
rect -3240 4800 -3160 4880
rect -3020 4800 -2940 4880
rect -710 4800 -630 4880
rect -520 4800 -440 4880
rect 1750 4790 1830 4870
rect 1930 4790 2010 4870
rect 4230 4790 4310 4870
rect 4400 4790 4480 4870
rect -4470 4540 -4390 4620
rect -4240 4540 -4160 4620
rect -1930 4530 -1850 4610
rect -1760 4530 -1680 4610
rect 540 4530 620 4610
rect 720 4530 800 4610
rect 2990 4530 3070 4610
rect 3180 4530 3260 4610
rect 5500 4530 5580 4610
rect 5670 4530 5750 4610
rect -4990 4390 -4860 4460
rect -3750 4390 -3620 4460
rect -2520 4390 -2390 4460
rect -1280 4390 -1150 4460
rect -40 4390 90 4460
rect 1190 4390 1320 4460
rect 2430 4390 2560 4460
rect 3660 4390 3790 4460
rect 4900 4390 5030 4460
rect -5720 4260 -5640 4340
rect -5510 4260 -5430 4340
rect -3250 4260 -3170 4340
rect -3010 4260 -2930 4340
rect -710 4260 -630 4340
rect -530 4260 -450 4340
rect 1760 4250 1840 4330
rect 1930 4250 2010 4330
rect 4230 4250 4310 4330
rect 4400 4250 4480 4330
rect -4450 4120 -4360 4200
rect -4270 4130 -4180 4210
rect -1920 4120 -1830 4200
rect -1760 4120 -1670 4200
rect 550 4120 640 4200
rect 710 4120 800 4200
rect 3000 4120 3090 4200
rect 3160 4120 3250 4200
rect 5500 4120 5590 4200
rect 5660 4120 5750 4200
rect -4470 3990 -4390 4070
rect -4240 3990 -4160 4070
rect -1940 4000 -1860 4080
rect -1750 4000 -1670 4080
rect 540 3990 620 4070
rect 730 3990 810 4070
rect 2990 3990 3070 4070
rect 3180 3990 3260 4070
rect 5500 3980 5580 4060
rect 5670 3980 5750 4060
rect -4990 3850 -4860 3920
rect -3750 3850 -3620 3920
rect -2520 3850 -2390 3920
rect -1280 3850 -1150 3920
rect -40 3850 90 3920
rect 1190 3850 1320 3920
rect 2430 3850 2560 3920
rect 3660 3850 3790 3920
rect 4900 3850 5030 3920
rect -5720 3720 -5640 3800
rect -5510 3720 -5430 3800
rect -3250 3710 -3170 3790
rect -3010 3710 -2930 3790
rect -710 3720 -630 3800
rect -520 3720 -440 3800
rect 1750 3710 1830 3790
rect 1940 3710 2020 3790
rect 4230 3700 4310 3780
rect 4400 3700 4480 3780
rect -8810 3260 -8720 3390
rect -8600 3260 -8510 3390
rect 8500 3290 8570 3380
rect 8660 3290 8730 3380
rect -3750 3200 -3620 3270
rect -2520 3190 -2390 3260
rect -2190 3190 -2110 3270
rect -2080 3190 -2000 3270
rect -1280 3190 -1150 3260
rect -40 3190 90 3260
rect 220 3190 300 3270
rect 330 3190 410 3270
rect 1190 3190 1320 3260
rect 2430 3210 2560 3280
rect 2680 3200 2760 3280
rect 2790 3200 2870 3280
rect 3660 3190 3790 3260
rect -3810 2920 -3720 3000
rect -3670 2920 -3580 3000
rect 1200 2940 1290 3020
rect 1340 2940 1430 3020
rect -2290 2800 -2180 2910
rect -1430 2800 -1320 2910
rect -220 2800 -110 2910
rect 630 2800 740 2910
rect -3810 2690 -3720 2770
rect -3670 2690 -3580 2770
rect 2200 2800 2310 2910
rect 3080 2800 3190 2910
rect 1200 2680 1290 2760
rect 1340 2680 1430 2760
rect -3480 2430 -3400 2510
rect -3330 2430 -3250 2510
rect -990 2450 -910 2530
rect -840 2450 -760 2530
rect 1490 2450 1570 2530
rect 1630 2450 1710 2530
rect -3030 2200 -2950 2280
rect -2920 2200 -2840 2280
rect -620 2170 -540 2250
rect 1830 2190 1910 2270
rect 1950 2190 2030 2270
rect 3030 2180 3110 2260
rect -1850 2020 -1770 2100
rect 560 2020 640 2100
rect -3110 1840 -3030 1920
rect 1780 1840 1860 1920
rect -3000 1700 -2890 1790
rect 1910 1700 2020 1790
rect -620 1550 -540 1630
rect 3030 1560 3110 1640
rect -2460 1400 -2370 1480
rect -2340 1400 -2250 1480
rect -1850 1400 -1770 1480
rect -10 1400 80 1480
rect 110 1400 200 1480
rect 560 1400 640 1480
rect 2420 1400 2510 1480
rect 2540 1400 2630 1480
rect -3110 1220 -3030 1300
rect 1780 1220 1860 1300
rect -1230 970 -1140 1050
rect 3650 990 3740 1070
rect -2460 800 -2370 880
rect -2340 800 -2250 880
rect -10 800 80 880
rect 110 800 200 880
rect 2420 800 2510 880
rect 2540 800 2630 880
rect -3810 640 -3720 720
rect -3670 640 -3580 720
rect 1200 640 1290 720
rect 1340 640 1430 720
rect -3060 490 -2940 590
rect -1840 490 -1720 590
rect -630 490 -510 590
rect -1230 370 -1140 450
rect 590 490 710 590
rect 1820 480 1940 580
rect 3030 490 3150 590
rect 3650 390 3740 470
rect -2460 200 -2370 280
rect -2340 200 -2250 280
rect -10 200 80 280
rect 110 200 200 280
rect 2420 200 2510 280
rect 2540 200 2630 280
rect -3810 20 -3720 100
rect -3670 20 -3580 100
rect 1200 40 1290 120
rect 1340 40 1430 120
<< metal2 >>
rect -2620 9100 -2330 9120
rect -2620 9030 -2600 9100
rect -2510 9030 -2430 9100
rect -2340 9030 -2330 9100
rect -2620 8990 -2330 9030
rect -2620 8910 -2600 8990
rect -2520 8910 -2430 8990
rect -2350 8910 -2330 8990
rect -130 9100 160 9120
rect -130 9030 -110 9100
rect -20 9030 60 9100
rect 150 9030 160 9100
rect -130 8990 160 9030
rect -3890 8750 -3600 8870
rect -3160 8860 -3010 8910
rect -3890 8670 -3870 8750
rect -3790 8670 -3700 8750
rect -3620 8670 -3600 8750
rect -3480 8820 -3400 8830
rect -3480 8730 -3400 8740
rect -3330 8820 -3250 8830
rect -3330 8730 -3250 8740
rect -3160 8790 -3150 8860
rect -3020 8790 -3010 8860
rect -3890 8210 -3600 8670
rect -3160 8320 -3010 8790
rect -3890 8130 -3870 8210
rect -3790 8130 -3700 8210
rect -3620 8130 -3600 8210
rect -3480 8280 -3400 8290
rect -3480 8190 -3400 8200
rect -3330 8280 -3250 8290
rect -3330 8190 -3250 8200
rect -3160 8250 -3150 8320
rect -3020 8250 -3010 8320
rect -3890 7670 -3600 8130
rect -3160 7780 -3010 8250
rect -2620 8450 -2330 8910
rect -2620 8370 -2600 8450
rect -2520 8370 -2430 8450
rect -2350 8370 -2330 8450
rect -2620 8050 -2330 8370
rect -2620 7980 -2590 8050
rect -2500 7980 -2450 8050
rect -2360 7980 -2330 8050
rect -2620 7910 -2330 7980
rect -2620 7830 -2600 7910
rect -2520 7830 -2430 7910
rect -2350 7830 -2330 7910
rect -2620 7820 -2330 7830
rect -1920 8860 -1770 8920
rect -1920 8790 -1910 8860
rect -1780 8790 -1770 8860
rect -1920 8320 -1770 8790
rect -1920 8250 -1910 8320
rect -1780 8250 -1770 8320
rect -3890 7590 -3870 7670
rect -3790 7590 -3700 7670
rect -3620 7590 -3600 7670
rect -3480 7740 -3400 7750
rect -3480 7650 -3400 7660
rect -3330 7740 -3250 7750
rect -3330 7650 -3250 7660
rect -3160 7710 -3150 7780
rect -3020 7710 -3010 7780
rect -3890 7570 -3600 7590
rect -3160 7240 -3010 7710
rect -1920 7780 -1770 8250
rect -1920 7710 -1910 7780
rect -1780 7710 -1770 7780
rect -2590 7520 -2510 7530
rect -2590 7430 -2510 7440
rect -2420 7520 -2340 7530
rect -2420 7430 -2340 7440
rect -3160 7170 -3150 7240
rect -3020 7170 -3010 7240
rect -3890 7130 -3600 7160
rect -3890 7050 -3870 7130
rect -3790 7050 -3700 7130
rect -3620 7050 -3600 7130
rect -3890 6550 -3600 7050
rect -3890 6470 -3870 6550
rect -3790 6470 -3700 6550
rect -3620 6470 -3600 6550
rect -9940 6270 -9810 6280
rect -9940 6120 -9810 6130
rect -9690 6270 -9560 6280
rect -9690 6120 -9560 6130
rect -3890 5940 -3600 6470
rect -3160 6660 -3010 7170
rect -3160 6590 -3150 6660
rect -3020 6590 -3010 6660
rect -3160 6080 -3010 6590
rect -2610 7390 -2320 7430
rect -2610 7310 -2590 7390
rect -2510 7310 -2420 7390
rect -2340 7310 -2320 7390
rect -2610 6810 -2320 7310
rect -1920 7240 -1770 7710
rect -1370 8750 -1080 8950
rect -130 8910 -110 8990
rect -30 8910 60 8990
rect 140 8910 160 8990
rect 2330 9110 2620 9150
rect 2330 9030 2350 9110
rect 2430 9030 2520 9110
rect 2600 9030 2620 9110
rect 2330 8980 2620 9030
rect -690 8860 -540 8910
rect -1370 8670 -1350 8750
rect -1270 8670 -1180 8750
rect -1100 8670 -1080 8750
rect -990 8820 -910 8830
rect -990 8730 -910 8740
rect -840 8820 -760 8830
rect -840 8730 -760 8740
rect -690 8790 -680 8860
rect -550 8790 -540 8860
rect -1370 8210 -1080 8670
rect -690 8320 -540 8790
rect -1370 8130 -1350 8210
rect -1270 8130 -1180 8210
rect -1100 8130 -1080 8210
rect -990 8280 -910 8290
rect -990 8190 -910 8200
rect -840 8280 -760 8290
rect -840 8190 -760 8200
rect -690 8250 -680 8320
rect -550 8250 -540 8320
rect -1370 7670 -1080 8130
rect -690 7780 -540 8250
rect -130 8450 160 8910
rect -130 8370 -110 8450
rect -30 8370 60 8450
rect 140 8370 160 8450
rect -130 8060 160 8370
rect -130 8050 50 8060
rect -130 7980 -110 8050
rect -20 7990 50 8050
rect 140 7990 160 8060
rect -20 7980 160 7990
rect -130 7920 160 7980
rect -130 7840 -110 7920
rect -30 7840 60 7920
rect 140 7840 160 7920
rect -130 7820 160 7840
rect 550 8860 700 8910
rect 550 8790 560 8860
rect 690 8790 700 8860
rect 550 8320 700 8790
rect 550 8250 560 8320
rect 690 8250 700 8320
rect -1370 7590 -1350 7670
rect -1270 7590 -1180 7670
rect -1100 7590 -1080 7670
rect -990 7740 -910 7750
rect -990 7650 -910 7660
rect -840 7740 -760 7750
rect -840 7650 -760 7660
rect -690 7710 -680 7780
rect -550 7710 -540 7780
rect -1370 7560 -1080 7590
rect -1920 7170 -1910 7240
rect -1780 7170 -1770 7240
rect -690 7240 -540 7710
rect 550 7780 700 8250
rect 550 7710 560 7780
rect 690 7710 700 7780
rect -110 7520 -30 7530
rect 60 7520 140 7530
rect -2190 7140 -2110 7150
rect -2190 7050 -2110 7060
rect -2080 7140 -2000 7150
rect -2080 7050 -2000 7060
rect -2610 6730 -2590 6810
rect -2510 6730 -2420 6810
rect -2340 6730 -2320 6810
rect -2610 6360 -2320 6730
rect -1920 6660 -1770 7170
rect -1920 6590 -1910 6660
rect -1780 6590 -1770 6660
rect -2190 6530 -2110 6540
rect -2190 6440 -2110 6450
rect -2080 6530 -2000 6540
rect -2080 6440 -2000 6450
rect -2610 6280 -2590 6360
rect -2500 6280 -2430 6360
rect -2340 6280 -2320 6360
rect -2610 6230 -2320 6280
rect -2610 6150 -2590 6230
rect -2510 6150 -2420 6230
rect -2340 6150 -2320 6230
rect -2610 6130 -2320 6150
rect -3160 6010 -3150 6080
rect -3020 6010 -3010 6080
rect -3160 5970 -3010 6010
rect -1920 6080 -1770 6590
rect -1920 6010 -1910 6080
rect -1780 6010 -1770 6080
rect -5720 5790 -5430 5870
rect -3810 5860 -3680 5940
rect -2210 5890 -1980 5980
rect -1920 5930 -1770 6010
rect -1388 7130 -1056 7180
rect -1388 7050 -1360 7130
rect -1280 7050 -1190 7130
rect -1110 7050 -1056 7130
rect -1388 6550 -1056 7050
rect -1388 6470 -1360 6550
rect -1280 6470 -1190 6550
rect -1110 6470 -1056 6550
rect -1388 5970 -1056 6470
rect -690 7170 -680 7240
rect -550 7170 -540 7240
rect -690 6660 -540 7170
rect -690 6590 -670 6660
rect -690 6080 -540 6590
rect -130 7400 160 7440
rect -130 7320 -110 7400
rect -30 7320 60 7400
rect 140 7320 160 7400
rect -130 6820 160 7320
rect 550 7240 700 7710
rect 1120 8750 1410 8950
rect 2330 8900 2350 8980
rect 2430 8900 2520 8980
rect 2600 8900 2620 8980
rect 1790 8860 1940 8900
rect 1120 8670 1140 8750
rect 1220 8670 1310 8750
rect 1390 8670 1410 8750
rect 1490 8820 1570 8830
rect 1490 8730 1570 8740
rect 1640 8820 1720 8830
rect 1640 8730 1720 8740
rect 1790 8790 1800 8860
rect 1930 8790 1940 8860
rect 1120 8210 1410 8670
rect 1790 8570 1940 8790
rect 1780 8320 1940 8570
rect 1120 8130 1140 8210
rect 1220 8130 1310 8210
rect 1390 8130 1410 8210
rect 1490 8280 1570 8290
rect 1490 8190 1570 8200
rect 1640 8280 1720 8290
rect 1640 8190 1720 8200
rect 1780 8250 1800 8320
rect 1930 8250 1940 8320
rect 1120 7660 1410 8130
rect 1780 7780 1940 8250
rect 1120 7580 1140 7660
rect 1220 7580 1310 7660
rect 1390 7580 1410 7660
rect 1500 7740 1580 7750
rect 1500 7650 1580 7660
rect 1640 7740 1720 7750
rect 1640 7650 1720 7660
rect 1780 7710 1800 7780
rect 1930 7710 1940 7780
rect 1780 7670 1940 7710
rect 2330 8440 2620 8900
rect 2330 8360 2350 8440
rect 2430 8360 2520 8440
rect 2600 8360 2620 8440
rect 2330 8060 2620 8360
rect 2330 7990 2350 8060
rect 2430 7990 2520 8060
rect 2600 7990 2620 8060
rect 2330 7900 2620 7990
rect 2330 7820 2350 7900
rect 2430 7820 2520 7900
rect 2600 7820 2620 7900
rect 1120 7560 1410 7580
rect 550 7170 560 7240
rect 690 7170 700 7240
rect 1780 7240 1930 7670
rect 2330 7570 2620 7820
rect 3020 8860 3170 8890
rect 3020 8790 3030 8860
rect 3160 8790 3170 8860
rect 3020 8320 3170 8790
rect 3020 8250 3030 8320
rect 3160 8250 3170 8320
rect 3020 7780 3170 8250
rect 3020 7710 3030 7780
rect 3160 7710 3170 7780
rect 2350 7520 2430 7530
rect 2520 7520 2600 7530
rect 1780 7170 1790 7240
rect 1920 7170 1930 7240
rect 220 7140 300 7150
rect 220 7050 300 7060
rect 330 7140 410 7150
rect 330 7050 410 7060
rect -130 6740 -110 6820
rect -30 6740 60 6820
rect 140 6740 160 6820
rect -130 6350 160 6740
rect 550 6660 700 7170
rect 550 6590 560 6660
rect 690 6590 700 6660
rect 220 6550 300 6560
rect 220 6460 300 6470
rect 330 6550 410 6560
rect 330 6460 410 6470
rect -130 6280 -110 6350
rect -30 6280 60 6350
rect 140 6280 160 6350
rect -130 6240 160 6280
rect -130 6160 -110 6240
rect -30 6160 60 6240
rect 140 6160 160 6240
rect -130 6140 160 6160
rect -690 6010 -680 6080
rect -550 6010 -540 6080
rect -690 5980 -540 6010
rect 550 6080 700 6590
rect 550 6010 560 6080
rect 690 6010 700 6080
rect 550 5980 700 6010
rect 1110 7130 1400 7170
rect 1110 7050 1130 7130
rect 1210 7050 1300 7130
rect 1380 7050 1400 7130
rect 1110 6540 1400 7050
rect 1110 6460 1130 6540
rect 1210 6460 1300 6540
rect 1380 6460 1400 6540
rect -1388 5890 -1360 5970
rect -1280 5890 -1190 5970
rect -1110 5890 -1056 5970
rect -3890 5850 -3810 5860
rect -3680 5850 -3600 5860
rect -1388 5832 -1056 5890
rect 220 5970 300 5980
rect 220 5880 300 5890
rect 330 5970 410 5980
rect 330 5880 410 5890
rect 1110 5970 1400 6460
rect 1780 6660 1930 7170
rect 1780 6590 1790 6660
rect 1920 6590 1930 6660
rect 1780 6080 1930 6590
rect 2330 7390 2620 7440
rect 2330 7310 2350 7390
rect 2430 7310 2520 7390
rect 2600 7310 2620 7390
rect 2330 6810 2620 7310
rect 3020 7240 3170 7710
rect 3570 8750 3860 9020
rect 3570 8670 3590 8750
rect 3670 8670 3760 8750
rect 3840 8670 3860 8750
rect 3570 8200 3860 8670
rect 3570 8120 3590 8200
rect 3670 8120 3760 8200
rect 3840 8120 3860 8200
rect 3570 7670 3860 8120
rect 3570 7590 3590 7670
rect 3670 7590 3760 7670
rect 3840 7590 3860 7670
rect 3570 7580 3860 7590
rect 3020 7170 3030 7240
rect 3160 7170 3170 7240
rect 2680 7130 2760 7140
rect 2680 7040 2760 7050
rect 2790 7130 2870 7140
rect 2790 7040 2870 7050
rect 2330 6730 2350 6810
rect 2430 6730 2520 6810
rect 2600 6730 2620 6810
rect 2330 6350 2620 6730
rect 3020 6660 3170 7170
rect 3020 6590 3030 6660
rect 3160 6590 3170 6660
rect 2680 6550 2760 6560
rect 2680 6460 2760 6470
rect 2790 6550 2870 6560
rect 2790 6460 2870 6470
rect 2330 6280 2350 6350
rect 2430 6280 2520 6350
rect 2600 6280 2620 6350
rect 2330 6230 2620 6280
rect 2330 6150 2350 6230
rect 2430 6150 2520 6230
rect 2600 6150 2620 6230
rect 2330 6140 2620 6150
rect 1780 6010 1790 6080
rect 1920 6010 1930 6080
rect 1780 5970 1930 6010
rect 3020 6080 3170 6590
rect 3020 6010 3030 6080
rect 3160 6010 3170 6080
rect 3020 5980 3170 6010
rect 3600 7130 3890 7220
rect 3600 7050 3620 7130
rect 3700 7050 3790 7130
rect 3870 7050 3890 7130
rect 3600 6550 3890 7050
rect 3600 6470 3620 6550
rect 3700 6470 3790 6550
rect 3870 6470 3890 6550
rect 2680 5970 2760 5980
rect 1110 5890 1130 5970
rect 1210 5890 1300 5970
rect 1380 5890 1400 5970
rect 1110 5870 1400 5890
rect 2680 5880 2760 5890
rect 2790 5970 2870 5980
rect 2790 5880 2870 5890
rect 3600 5970 3890 6470
rect 9560 6440 9690 6450
rect 9560 6290 9690 6300
rect 9820 6440 9950 6450
rect 9820 6290 9950 6300
rect 3600 5890 3620 5970
rect 3700 5890 3790 5970
rect 3870 5890 3890 5970
rect 3600 5870 3890 5890
rect -5720 5680 -5700 5790
rect -5610 5680 -5540 5790
rect -5450 5680 -5430 5790
rect 4210 5740 4500 5780
rect -5720 5420 -5430 5680
rect -4470 5700 -4160 5720
rect -4390 5620 -4240 5700
rect -5640 5340 -5510 5420
rect -5720 4880 -5430 5340
rect -5640 4800 -5510 4880
rect -5720 4340 -5430 4800
rect -5640 4260 -5510 4340
rect -5720 3800 -5430 4260
rect -5000 5540 -4850 5570
rect -5000 5470 -4990 5540
rect -4860 5470 -4850 5540
rect -5000 5010 -4850 5470
rect -5000 4940 -4990 5010
rect -4860 4940 -4850 5010
rect -5000 4460 -4850 4940
rect -5000 4390 -4990 4460
rect -4860 4390 -4850 4460
rect -5000 3920 -4850 4390
rect -4470 5280 -4160 5620
rect -1940 5690 -1650 5720
rect -1940 5610 -1920 5690
rect -1840 5610 -1750 5690
rect -1670 5610 -1650 5690
rect -4470 5200 -4450 5280
rect -4360 5200 -4270 5280
rect -4180 5200 -4160 5280
rect -4470 5160 -4160 5200
rect -4390 5080 -4240 5160
rect -4470 4620 -4160 5080
rect -4390 4540 -4240 4620
rect -4470 4210 -4160 4540
rect -4470 4200 -4270 4210
rect -4470 4120 -4450 4200
rect -4360 4130 -4270 4200
rect -4180 4130 -4160 4210
rect -4360 4120 -4160 4130
rect -4470 4070 -4160 4120
rect -4390 3990 -4240 4070
rect -4470 3980 -4160 3990
rect -3760 5540 -3610 5580
rect -3760 5470 -3750 5540
rect -3620 5470 -3610 5540
rect -3760 5000 -3610 5470
rect -2530 5540 -2380 5570
rect -2530 5470 -2520 5540
rect -2390 5470 -2380 5540
rect -3760 4930 -3750 5000
rect -3620 4930 -3610 5000
rect -3760 4460 -3610 4930
rect -3760 4390 -3750 4460
rect -3620 4390 -3610 4460
rect -5000 3850 -4990 3920
rect -4860 3850 -4850 3920
rect -5000 3810 -4850 3850
rect -3760 3920 -3610 4390
rect -3760 3850 -3750 3920
rect -3620 3850 -3610 3920
rect -5640 3720 -5510 3800
rect -5720 3710 -5430 3720
rect -8810 3390 -8720 3400
rect -8810 3250 -8720 3260
rect -8600 3390 -8510 3400
rect -8600 3250 -8510 3260
rect -3760 3270 -3610 3850
rect -3250 5420 -2930 5450
rect -3250 5340 -3240 5420
rect -3160 5340 -3020 5420
rect -2940 5340 -2930 5420
rect -3250 4880 -2930 5340
rect -3250 4800 -3240 4880
rect -3160 4800 -3020 4880
rect -2940 4800 -2930 4880
rect -3250 4340 -2930 4800
rect -3170 4260 -3010 4340
rect -3250 3870 -2930 4260
rect -2530 5000 -2380 5470
rect -2530 4930 -2520 5000
rect -2390 4930 -2380 5000
rect -2530 4460 -2380 4930
rect -2530 4390 -2520 4460
rect -2390 4390 -2380 4460
rect -2530 3920 -2380 4390
rect -1940 5280 -1650 5610
rect 530 5690 820 5730
rect 530 5610 540 5690
rect 620 5610 730 5690
rect 810 5610 820 5690
rect -1940 5200 -1920 5280
rect -1830 5200 -1760 5280
rect -1670 5200 -1650 5280
rect -1940 5160 -1650 5200
rect -1940 5150 -1750 5160
rect -1940 5070 -1920 5150
rect -1840 5080 -1750 5150
rect -1670 5080 -1650 5160
rect -1840 5070 -1650 5080
rect -1940 4610 -1650 5070
rect -1940 4530 -1930 4610
rect -1850 4530 -1760 4610
rect -1680 4530 -1650 4610
rect -1940 4200 -1650 4530
rect -1940 4120 -1920 4200
rect -1830 4120 -1760 4200
rect -1670 4120 -1650 4200
rect -1940 4080 -1650 4120
rect -1860 4000 -1750 4080
rect -1670 4000 -1650 4080
rect -1940 3970 -1650 4000
rect -1290 5540 -1140 5570
rect -1290 5470 -1280 5540
rect -1150 5470 -1140 5540
rect -50 5540 100 5560
rect -1290 5000 -1140 5470
rect -1290 4930 -1280 5000
rect -1150 4930 -1140 5000
rect -1290 4460 -1140 4930
rect -1290 4390 -1280 4460
rect -1150 4390 -1140 4460
rect -3250 3790 -2840 3870
rect -3170 3710 -3010 3790
rect -2930 3710 -2840 3790
rect -3250 3610 -2840 3710
rect -3760 3200 -3750 3270
rect -3620 3200 -3610 3270
rect -3760 3190 -3610 3200
rect -3810 3000 -3720 3010
rect -3670 3000 -3580 3010
rect -3720 2920 -3670 2990
rect -3810 2770 -3580 2920
rect -3720 2690 -3670 2770
rect -3810 720 -3580 2690
rect -3500 2510 -3230 2520
rect -3500 2430 -3480 2510
rect -3400 2430 -3330 2510
rect -3250 2430 -3230 2510
rect -3480 2420 -3400 2430
rect -3330 2420 -3250 2430
rect -3030 2310 -2840 3610
rect -2530 3850 -2520 3920
rect -2390 3850 -2380 3920
rect -2530 3260 -2380 3850
rect -1290 3920 -1140 4390
rect -1290 3850 -1280 3920
rect -1150 3850 -1140 3920
rect -2530 3190 -2520 3260
rect -2390 3190 -2380 3260
rect -2530 3140 -2380 3190
rect -2190 3270 -2110 3280
rect -2190 3180 -2110 3190
rect -2080 3270 -2000 3280
rect -2080 3180 -2000 3190
rect -1290 3260 -1140 3850
rect -1290 3190 -1280 3260
rect -1150 3190 -1140 3260
rect -1290 3100 -1140 3190
rect -720 5420 -430 5510
rect -720 5340 -710 5420
rect -630 5340 -530 5420
rect -450 5340 -430 5420
rect -720 4880 -430 5340
rect -720 4800 -710 4880
rect -630 4800 -520 4880
rect -440 4800 -430 4880
rect -720 4340 -430 4800
rect -720 4260 -710 4340
rect -630 4260 -530 4340
rect -450 4260 -430 4340
rect -720 3800 -430 4260
rect -720 3720 -710 3800
rect -630 3720 -520 3800
rect -440 3720 -430 3800
rect -2290 2910 -2180 2920
rect -2290 2790 -2180 2800
rect -1430 2910 -1320 2920
rect -1430 2790 -1320 2800
rect -990 2530 -910 2540
rect -990 2440 -910 2450
rect -840 2530 -760 2540
rect -840 2440 -760 2450
rect -3120 2280 -2810 2310
rect -3120 2200 -3030 2280
rect -2950 2200 -2920 2280
rect -2840 2200 -2810 2280
rect -720 2250 -430 3720
rect -50 5470 -40 5540
rect 90 5470 100 5540
rect -50 5000 100 5470
rect -50 4930 -40 5000
rect 90 4930 100 5000
rect -50 4460 100 4930
rect -50 4390 -40 4460
rect 90 4390 100 4460
rect -50 3920 100 4390
rect 530 5280 820 5610
rect 2980 5690 3270 5720
rect 2980 5610 2990 5690
rect 3070 5610 3180 5690
rect 3260 5610 3270 5690
rect 530 5200 550 5280
rect 640 5200 710 5280
rect 800 5200 820 5280
rect 530 5160 820 5200
rect 530 5080 540 5160
rect 620 5080 730 5160
rect 810 5080 820 5160
rect 530 4610 820 5080
rect 530 4530 540 4610
rect 620 4530 720 4610
rect 800 4530 820 4610
rect 530 4200 820 4530
rect 530 4120 550 4200
rect 640 4120 710 4200
rect 800 4120 820 4200
rect 530 4070 820 4120
rect 530 3990 540 4070
rect 620 3990 730 4070
rect 810 3990 820 4070
rect 530 3980 820 3990
rect 1180 5540 1330 5570
rect 1180 5470 1190 5540
rect 1320 5470 1330 5540
rect 2420 5540 2570 5590
rect 1180 5000 1330 5470
rect 1180 4930 1190 5000
rect 1320 4930 1330 5000
rect 1180 4460 1330 4930
rect 1180 4390 1190 4460
rect 1320 4390 1330 4460
rect -50 3850 -40 3920
rect 90 3850 100 3920
rect -50 3260 100 3850
rect 1180 3920 1330 4390
rect 1180 3850 1190 3920
rect 1320 3850 1330 3920
rect -50 3190 -40 3260
rect 90 3190 100 3260
rect -50 3120 100 3190
rect 220 3270 300 3280
rect 220 3180 300 3190
rect 330 3270 410 3280
rect 330 3180 410 3190
rect 1180 3260 1330 3850
rect 1740 5410 2030 5510
rect 1740 5330 1750 5410
rect 1830 5330 1930 5410
rect 2010 5330 2030 5410
rect 1740 4870 2030 5330
rect 1740 4790 1750 4870
rect 1830 4790 1930 4870
rect 2010 4790 2030 4870
rect 1740 4330 2030 4790
rect 1740 4250 1760 4330
rect 1840 4250 1930 4330
rect 2010 4250 2030 4330
rect 1740 3890 2030 4250
rect 2420 5470 2430 5540
rect 2560 5470 2570 5540
rect 2420 5000 2570 5470
rect 2420 4930 2430 5000
rect 2560 4930 2570 5000
rect 2420 4460 2570 4930
rect 2420 4390 2430 4460
rect 2560 4390 2570 4460
rect 2420 3920 2570 4390
rect 1740 3790 2040 3890
rect 1740 3710 1750 3790
rect 1830 3710 1940 3790
rect 2020 3710 2040 3790
rect 1740 3690 2040 3710
rect 1180 3190 1190 3260
rect 1320 3190 1330 3260
rect 1180 3180 1330 3190
rect 1200 3020 1290 3030
rect 1340 3020 1430 3030
rect 1290 2940 1340 3020
rect -220 2910 -110 2920
rect -220 2790 -110 2800
rect 630 2910 740 2920
rect 630 2790 740 2800
rect -720 2200 -620 2250
rect -3120 2180 -2810 2200
rect -540 2200 -430 2250
rect 1200 2760 1430 2940
rect 1290 2680 1340 2760
rect -1850 2100 -1770 2130
rect -3110 1920 -3030 1950
rect -3110 1830 -3030 1840
rect -3110 1790 -2850 1830
rect -3110 1700 -3000 1790
rect -2890 1700 -2850 1790
rect -3110 1660 -2850 1700
rect -3110 1300 -3030 1660
rect -3110 1210 -3030 1220
rect -2460 1480 -2250 1500
rect -2370 1400 -2340 1480
rect -3720 640 -3670 720
rect -3810 100 -3580 640
rect -2460 880 -2250 1400
rect -1850 1480 -1770 2020
rect -620 1630 -540 2170
rect -620 1540 -540 1550
rect 560 2100 640 2130
rect -1850 1390 -1770 1400
rect -10 1480 200 1500
rect 80 1400 110 1480
rect -2370 800 -2340 880
rect -3060 590 -2940 600
rect -3060 480 -2940 490
rect -2460 280 -2250 800
rect -1230 1050 -1140 1080
rect -1840 590 -1720 600
rect -1840 480 -1720 490
rect -1230 450 -1140 970
rect -10 880 200 1400
rect 560 1480 640 2020
rect 560 1390 640 1400
rect 80 800 110 880
rect -630 590 -510 600
rect -630 480 -510 490
rect -1230 360 -1140 370
rect -2370 200 -2340 280
rect -2460 190 -2250 200
rect -10 280 200 800
rect 1200 720 1430 2680
rect 1490 2530 1570 2540
rect 1490 2440 1570 2450
rect 1630 2530 1710 2540
rect 1630 2440 1710 2450
rect 1820 2270 2040 3690
rect 2420 3850 2430 3920
rect 2560 3850 2570 3920
rect 2420 3280 2570 3850
rect 2980 5280 3270 5610
rect 4210 5660 4230 5740
rect 4310 5660 4400 5740
rect 4480 5660 4500 5740
rect 2980 5200 3000 5280
rect 3090 5200 3160 5280
rect 3250 5200 3270 5280
rect 2980 5150 3270 5200
rect 2980 5070 2990 5150
rect 3070 5070 3180 5150
rect 3260 5070 3270 5150
rect 2980 4610 3270 5070
rect 2980 4530 2990 4610
rect 3070 4530 3180 4610
rect 3260 4530 3270 4610
rect 2980 4200 3270 4530
rect 2980 4120 3000 4200
rect 3090 4120 3160 4200
rect 3250 4120 3270 4200
rect 2980 4070 3270 4120
rect 2980 3990 2990 4070
rect 3070 3990 3180 4070
rect 3260 3990 3270 4070
rect 2980 3740 3270 3990
rect 3650 5540 3800 5580
rect 3650 5470 3660 5540
rect 3790 5470 3800 5540
rect 3650 5000 3800 5470
rect 3650 4930 3660 5000
rect 3790 4930 3800 5000
rect 3650 4460 3800 4930
rect 3650 4390 3660 4460
rect 3790 4390 3800 4460
rect 3650 3920 3800 4390
rect 3650 3850 3660 3920
rect 3790 3850 3800 3920
rect 2420 3210 2430 3280
rect 2560 3210 2570 3280
rect 2420 3150 2570 3210
rect 2680 3280 2760 3290
rect 2680 3190 2760 3200
rect 2790 3280 2870 3290
rect 2790 3190 2870 3200
rect 3650 3260 3800 3850
rect 4210 5410 4500 5660
rect 5480 5690 5770 5710
rect 5480 5610 5500 5690
rect 5580 5610 5670 5690
rect 5750 5610 5770 5690
rect 4210 5330 4230 5410
rect 4310 5330 4400 5410
rect 4480 5330 4500 5410
rect 4210 4870 4500 5330
rect 4210 4790 4230 4870
rect 4310 4790 4400 4870
rect 4480 4790 4500 4870
rect 4210 4330 4500 4790
rect 4210 4250 4230 4330
rect 4310 4250 4400 4330
rect 4480 4250 4500 4330
rect 4210 3780 4500 4250
rect 4890 5540 5040 5580
rect 4890 5470 4900 5540
rect 5030 5470 5040 5540
rect 4890 5000 5040 5470
rect 4890 4930 4900 5000
rect 5030 4930 5040 5000
rect 4890 4460 5040 4930
rect 4890 4390 4900 4460
rect 5030 4390 5040 4460
rect 4890 3920 5040 4390
rect 5480 5280 5770 5610
rect 5480 5200 5500 5280
rect 5590 5200 5660 5280
rect 5750 5200 5770 5280
rect 5480 5150 5770 5200
rect 5480 5070 5500 5150
rect 5580 5070 5670 5150
rect 5750 5070 5770 5150
rect 5480 4610 5770 5070
rect 5480 4530 5500 4610
rect 5580 4530 5670 4610
rect 5750 4530 5770 4610
rect 5480 4200 5770 4530
rect 5480 4120 5500 4200
rect 5590 4120 5660 4200
rect 5750 4120 5770 4200
rect 5480 4060 5770 4120
rect 5480 3980 5500 4060
rect 5580 3980 5670 4060
rect 5750 3980 5770 4060
rect 5480 3960 5770 3980
rect 4890 3850 4900 3920
rect 5030 3850 5040 3920
rect 4890 3820 5040 3850
rect 4210 3700 4230 3780
rect 4310 3700 4400 3780
rect 4480 3700 4500 3780
rect 4210 3690 4500 3700
rect 8500 3380 8570 3390
rect 8500 3280 8570 3290
rect 8660 3380 8730 3390
rect 8660 3280 8730 3290
rect 3650 3190 3660 3260
rect 3790 3190 3800 3260
rect 3650 3150 3800 3190
rect 2200 2910 2310 2920
rect 2200 2790 2310 2800
rect 3080 2910 3190 2920
rect 3080 2790 3190 2800
rect 1820 2190 1830 2270
rect 1910 2190 1950 2270
rect 2030 2190 2040 2270
rect 2980 2260 3270 2270
rect 2980 2220 3030 2260
rect 1820 2180 2040 2190
rect 3110 2220 3270 2260
rect 1780 1920 1860 1950
rect 1780 1830 1860 1840
rect 1780 1790 2050 1830
rect 1780 1700 1910 1790
rect 2020 1700 2050 1790
rect 1780 1660 2050 1700
rect 1780 1300 1860 1660
rect 3030 1640 3110 2180
rect 3030 1550 3110 1560
rect 1780 1210 1860 1220
rect 2420 1480 2630 1500
rect 2510 1400 2540 1480
rect 1290 640 1340 720
rect 590 590 710 600
rect 590 480 710 490
rect 80 200 110 280
rect -10 190 200 200
rect -3720 20 -3670 100
rect 1200 120 1430 640
rect 2420 880 2630 1400
rect 2510 800 2540 880
rect 1820 580 1940 590
rect 1820 470 1940 480
rect 2420 280 2630 800
rect 3650 1070 3740 1100
rect 3030 590 3150 600
rect 3030 480 3150 490
rect 3650 470 3740 990
rect 3650 380 3740 390
rect 2510 200 2540 280
rect 2420 190 2630 200
rect 1290 40 1340 120
rect 1200 30 1430 40
rect -3810 10 -3580 20
<< via2 >>
rect -2600 9030 -2510 9100
rect -2430 9030 -2340 9100
rect -110 9030 -20 9100
rect 60 9030 150 9100
rect -3480 8740 -3400 8820
rect -3330 8740 -3250 8820
rect -3480 8200 -3400 8280
rect -3330 8200 -3250 8280
rect -2590 7980 -2500 8050
rect -2450 7980 -2360 8050
rect -3480 7660 -3400 7740
rect -3330 7660 -3250 7740
rect -2590 7440 -2510 7520
rect -2420 7440 -2340 7520
rect -9940 6130 -9810 6270
rect -9690 6130 -9560 6270
rect 2350 9030 2430 9110
rect 2520 9030 2600 9110
rect -990 8740 -910 8820
rect -840 8740 -760 8820
rect -990 8200 -910 8280
rect -840 8200 -760 8280
rect -110 7980 -20 8050
rect 50 7990 140 8060
rect -990 7660 -910 7740
rect -840 7660 -760 7740
rect -110 7440 -30 7520
rect 60 7440 140 7520
rect -2190 7060 -2110 7140
rect -2080 7060 -2000 7140
rect -2190 6450 -2110 6530
rect -2080 6450 -2000 6530
rect -2590 6280 -2500 6360
rect -2430 6280 -2340 6360
rect 1490 8740 1570 8820
rect 1640 8740 1720 8820
rect 1490 8200 1570 8280
rect 1640 8200 1720 8280
rect 1500 7660 1580 7740
rect 1640 7660 1720 7740
rect 2350 7990 2430 8060
rect 2520 7990 2600 8060
rect 2350 7440 2430 7520
rect 2520 7440 2600 7520
rect 220 7060 300 7140
rect 330 7060 410 7140
rect 220 6470 300 6550
rect 330 6470 410 6550
rect -110 6280 -30 6350
rect 60 6280 140 6350
rect 220 5890 300 5970
rect 330 5890 410 5970
rect 2680 7050 2760 7130
rect 2790 7050 2870 7130
rect 2680 6470 2760 6550
rect 2790 6470 2870 6550
rect 2350 6280 2430 6350
rect 2520 6280 2600 6350
rect 2680 5890 2760 5970
rect 2790 5890 2870 5970
rect 9560 6300 9690 6440
rect 9820 6300 9950 6440
rect -5700 5680 -5610 5790
rect -5540 5680 -5450 5790
rect -4450 5200 -4360 5280
rect -4270 5200 -4180 5280
rect -4450 4120 -4360 4200
rect -4270 4130 -4180 4210
rect -8810 3260 -8720 3390
rect -8600 3260 -8510 3390
rect -1920 5200 -1830 5280
rect -1760 5200 -1670 5280
rect -1920 4120 -1830 4200
rect -1760 4120 -1670 4200
rect -3480 2430 -3400 2510
rect -3330 2430 -3250 2510
rect -2190 3190 -2110 3270
rect -2080 3190 -2000 3270
rect -2290 2800 -2180 2910
rect -1430 2800 -1320 2910
rect -990 2450 -910 2530
rect -840 2450 -760 2530
rect 550 5200 640 5280
rect 710 5200 800 5280
rect 550 4120 640 4200
rect 710 4120 800 4200
rect 220 3190 300 3270
rect 330 3190 410 3270
rect -220 2800 -110 2910
rect 630 2800 740 2910
rect -3000 1700 -2890 1790
rect -3060 490 -2940 590
rect -1840 490 -1720 590
rect -630 490 -510 590
rect 1490 2450 1570 2530
rect 1630 2450 1710 2530
rect 4230 5660 4310 5740
rect 4400 5660 4480 5740
rect 3000 5200 3090 5280
rect 3160 5200 3250 5280
rect 3000 4120 3090 4200
rect 3160 4120 3250 4200
rect 2680 3200 2760 3280
rect 2790 3200 2870 3280
rect 5500 5200 5590 5280
rect 5660 5200 5750 5280
rect 5500 4120 5590 4200
rect 5660 4120 5750 4200
rect 8500 3290 8570 3380
rect 8660 3290 8730 3380
rect 2200 2800 2310 2910
rect 3080 2800 3190 2910
rect 1910 1700 2020 1790
rect 590 490 710 590
rect 3030 490 3150 590
<< metal3 >>
rect -9960 13130 -9520 13180
rect -9960 13000 -9930 13130
rect -9830 13000 -9670 13130
rect -9570 13000 -9520 13130
rect -9960 6270 -9520 13000
rect 9540 13130 9970 13190
rect 9540 13000 9560 13130
rect 9670 13000 9820 13130
rect 9930 13000 9970 13130
rect -4650 9110 6930 9350
rect -4650 9100 2350 9110
rect -4650 9030 -2600 9100
rect -2510 9030 -2430 9100
rect -2340 9030 -110 9100
rect -20 9030 60 9100
rect 150 9030 2350 9100
rect 2430 9030 2520 9110
rect 2600 9030 6930 9110
rect -4650 8990 6930 9030
rect -3500 8820 -3230 8840
rect -3500 8740 -3480 8820
rect -3400 8740 -3330 8820
rect -3250 8740 -3230 8820
rect -3500 8720 -3230 8740
rect -1010 8820 -740 8830
rect -1010 8740 -990 8820
rect -910 8740 -840 8820
rect -760 8740 -740 8820
rect -1010 8720 -740 8740
rect 1470 8820 1740 8840
rect 1470 8740 1490 8820
rect 1570 8740 1640 8820
rect 1720 8740 1740 8820
rect 1470 8720 1740 8740
rect -3500 8280 -3230 8300
rect -3500 8200 -3480 8280
rect -3400 8200 -3330 8280
rect -3250 8200 -3230 8280
rect -3500 8180 -3230 8200
rect -1010 8280 -740 8290
rect -1010 8200 -990 8280
rect -910 8200 -840 8280
rect -760 8200 -740 8280
rect -1010 8180 -740 8200
rect 1470 8280 1740 8300
rect 1470 8200 1490 8280
rect 1570 8200 1640 8280
rect 1720 8200 1740 8280
rect 1470 8180 1740 8200
rect 6520 8120 6930 8990
rect -4890 8060 6930 8120
rect -4890 8050 50 8060
rect -4890 7980 -2590 8050
rect -2500 7980 -2450 8050
rect -2360 7980 -110 8050
rect -20 7990 50 8050
rect 140 7990 2350 8060
rect 2430 7990 2520 8060
rect 2600 7990 6930 8060
rect -20 7980 6930 7990
rect -4890 7890 6930 7980
rect -3500 7740 -3230 7770
rect -3500 7660 -3480 7740
rect -3400 7660 -3330 7740
rect -3250 7660 -3230 7740
rect -3500 7640 -3230 7660
rect -1010 7740 -740 7750
rect -1010 7660 -990 7740
rect -910 7660 -840 7740
rect -760 7660 -740 7740
rect -1010 7640 -740 7660
rect 1470 7740 1740 7770
rect 1470 7660 1500 7740
rect 1580 7660 1640 7740
rect 1720 7660 1740 7740
rect 1470 7640 1740 7660
rect 6520 7530 6930 7890
rect -4500 7520 6930 7530
rect -4500 7440 -2590 7520
rect -2510 7440 -2420 7520
rect -2340 7440 -110 7520
rect -30 7440 60 7520
rect 140 7440 2350 7520
rect 2430 7440 2520 7520
rect 2600 7440 6930 7520
rect -4500 7310 6930 7440
rect -2210 7140 -1980 7160
rect -2210 7060 -2190 7140
rect -2110 7060 -2080 7140
rect -2000 7060 -1980 7140
rect -2210 7030 -1980 7060
rect 200 7140 430 7160
rect 200 7060 220 7140
rect 300 7060 330 7140
rect 410 7060 430 7140
rect 200 7050 430 7060
rect 2660 7130 2890 7140
rect 2660 7050 2680 7130
rect 2760 7050 2790 7130
rect 2870 7050 2890 7130
rect 2660 7030 2890 7050
rect 200 6550 430 6560
rect -2210 6530 -1980 6540
rect -2210 6450 -2190 6530
rect -2110 6450 -2080 6530
rect -2000 6450 -1980 6530
rect 200 6470 220 6550
rect 300 6470 330 6550
rect 410 6470 430 6550
rect 200 6450 430 6470
rect 2660 6550 2890 6560
rect 2660 6470 2680 6550
rect 2760 6470 2790 6550
rect 2870 6470 2890 6550
rect 2660 6450 2890 6470
rect -2210 6440 -1980 6450
rect 6520 6370 6930 7310
rect -9960 6130 -9940 6270
rect -9810 6130 -9690 6270
rect -9560 6130 -9520 6270
rect -4580 6360 6930 6370
rect -4580 6280 -2590 6360
rect -2500 6280 -2430 6360
rect -2340 6350 6930 6360
rect -2340 6280 -110 6350
rect -30 6280 60 6350
rect 140 6280 2350 6350
rect 2430 6280 2520 6350
rect 2600 6280 6930 6350
rect 9540 6440 9970 13000
rect 9540 6300 9560 6440
rect 9690 6300 9820 6440
rect 9950 6300 9970 6440
rect 9540 6290 9970 6300
rect -4580 6190 6930 6280
rect -9960 6110 -9520 6130
rect -2210 5970 -1980 5990
rect -2210 5890 -2190 5970
rect -2110 5890 -2080 5970
rect -2000 5890 -1980 5970
rect -2210 5870 -1980 5890
rect 200 5970 430 5980
rect 200 5890 220 5970
rect 300 5890 330 5970
rect 410 5890 430 5970
rect 200 5870 430 5890
rect 2660 5970 2890 5980
rect 2660 5890 2680 5970
rect 2760 5890 2790 5970
rect 2870 5890 2890 5970
rect 2660 5870 2890 5890
rect -5720 5790 -5430 5810
rect -5720 5680 -5700 5790
rect -5610 5680 -5540 5790
rect -5450 5680 -5430 5790
rect -5720 5670 -5430 5680
rect 4210 5740 4502 5750
rect 4210 5660 4230 5740
rect 4310 5660 4400 5740
rect 4480 5660 4502 5740
rect 4210 5652 4502 5660
rect 6520 5460 6930 6190
rect -6730 5280 6930 5460
rect -6730 5200 -4450 5280
rect -4360 5200 -4270 5280
rect -4180 5200 -1920 5280
rect -1830 5200 -1760 5280
rect -1670 5200 550 5280
rect 640 5200 710 5280
rect 800 5200 3000 5280
rect 3090 5200 3160 5280
rect 3250 5200 5500 5280
rect 5590 5200 5660 5280
rect 5750 5200 6930 5280
rect -6730 5100 6930 5200
rect 6520 4330 6930 5100
rect -6360 4210 6930 4330
rect -6360 4200 -4270 4210
rect -6360 4120 -4450 4200
rect -4360 4130 -4270 4200
rect -4180 4200 6930 4210
rect -4180 4130 -1920 4200
rect -4360 4120 -1920 4130
rect -1830 4120 -1760 4200
rect -1670 4120 550 4200
rect 640 4120 710 4200
rect 800 4120 3000 4200
rect 3090 4120 3160 4200
rect 3250 4120 5500 4200
rect 5590 4120 5660 4200
rect 5750 4120 6930 4200
rect -6360 3990 6930 4120
rect -8830 3390 -8480 3400
rect -8830 3260 -8810 3390
rect -8720 3260 -8600 3390
rect -8510 3260 -8480 3390
rect 8490 3380 8750 3390
rect 8490 3290 8500 3380
rect 8570 3290 8660 3380
rect 8730 3290 8750 3380
rect -8830 3060 -8480 3260
rect -2210 3270 -1980 3280
rect -2210 3190 -2190 3270
rect -2110 3190 -2080 3270
rect -2000 3190 -1980 3270
rect -2210 3180 -1980 3190
rect 200 3270 430 3290
rect 200 3190 220 3270
rect 300 3190 330 3270
rect 410 3190 430 3270
rect 2660 3280 2890 3290
rect 2660 3200 2680 3280
rect 2760 3200 2790 3280
rect 2870 3200 2890 3280
rect 2660 3190 2890 3200
rect 200 3180 430 3190
rect -9330 3050 -4660 3060
rect 8490 3050 8750 3290
rect -9330 2910 9880 3050
rect -9330 2830 -2290 2910
rect -4940 2800 -2290 2830
rect -2180 2800 -1430 2910
rect -1320 2800 -220 2910
rect -110 2800 630 2910
rect 740 2800 2200 2910
rect 2310 2800 3080 2910
rect 3190 2800 9880 2910
rect -4940 2690 9880 2800
rect -4940 1990 -4660 2690
rect 4830 2680 9880 2690
rect -1010 2530 -740 2540
rect -3500 2510 -3230 2530
rect -3500 2430 -3480 2510
rect -3400 2430 -3330 2510
rect -3250 2430 -3230 2510
rect -1010 2450 -990 2530
rect -910 2450 -840 2530
rect -760 2450 -740 2530
rect -1010 2430 -740 2450
rect 1470 2530 1740 2540
rect 1470 2450 1490 2530
rect 1570 2450 1630 2530
rect 1710 2450 1740 2530
rect 1470 2430 1740 2450
rect -3500 2400 -3230 2430
rect 4900 1990 5120 2680
rect -4940 1790 5120 1990
rect -4940 1700 -3000 1790
rect -2890 1700 1910 1790
rect 2020 1700 5120 1790
rect -4940 1530 5120 1700
rect -4940 810 -4660 1530
rect 4900 810 5120 1530
rect -4940 590 5120 810
rect -4940 490 -3060 590
rect -2940 490 -1840 590
rect -1720 490 -630 590
rect -510 490 590 590
rect 710 580 3030 590
rect 710 490 1820 580
rect -4940 480 1820 490
rect 1940 490 3030 580
rect 3150 490 5120 590
rect 1940 480 5120 490
rect -4940 350 5120 480
<< via3 >>
rect -9930 13000 -9830 13130
rect -9670 13000 -9570 13130
rect 9560 13000 9670 13130
rect 9820 13000 9930 13130
rect -3480 8740 -3400 8820
rect -3330 8740 -3250 8820
rect -990 8740 -910 8820
rect -840 8740 -760 8820
rect 1490 8740 1570 8820
rect 1640 8740 1720 8820
rect -3480 8200 -3400 8280
rect -3330 8200 -3250 8280
rect -990 8200 -910 8280
rect -840 8200 -760 8280
rect 1490 8200 1570 8280
rect 1640 8200 1720 8280
rect -3480 7660 -3400 7740
rect -3330 7660 -3250 7740
rect -990 7660 -910 7740
rect -840 7660 -760 7740
rect 1500 7660 1580 7740
rect 1640 7660 1720 7740
rect -2190 7060 -2110 7140
rect -2080 7060 -2000 7140
rect 220 7060 300 7140
rect 330 7060 410 7140
rect 2680 7050 2760 7130
rect 2790 7050 2870 7130
rect -2190 6450 -2110 6530
rect -2080 6450 -2000 6530
rect 220 6470 300 6550
rect 330 6470 410 6550
rect 2680 6470 2760 6550
rect 2790 6470 2870 6550
rect -2190 5890 -2110 5970
rect -2080 5890 -2000 5970
rect 220 5890 300 5970
rect 330 5890 410 5970
rect 2680 5890 2760 5970
rect 2790 5890 2870 5970
rect -5700 5680 -5610 5790
rect -5540 5680 -5450 5790
rect 4230 5660 4310 5740
rect 4400 5660 4480 5740
rect -2190 3190 -2110 3270
rect -2080 3190 -2000 3270
rect 220 3190 300 3270
rect 330 3190 410 3270
rect 2680 3200 2760 3280
rect 2790 3200 2870 3280
rect -3480 2430 -3400 2510
rect -3330 2430 -3250 2510
rect -990 2450 -910 2530
rect -840 2450 -760 2530
rect 1490 2450 1570 2530
rect 1630 2450 1710 2530
rect 1820 480 1940 580
<< metal4 >>
rect -9970 13130 9970 13190
rect -9970 13000 -9930 13130
rect -9830 13000 -9670 13130
rect -9570 13000 9560 13130
rect 9670 13000 9820 13130
rect 9930 13000 9970 13130
rect -9970 12950 9970 13000
rect -4230 11330 4250 11690
rect -3920 9510 -3750 11330
rect -5720 9320 -3750 9510
rect 3720 9530 3880 11330
rect 3720 9400 4500 9530
rect -5720 5790 -5430 9320
rect -5720 5680 -5700 5790
rect -5610 5680 -5540 5790
rect -5450 5680 -5430 5790
rect -5720 5460 -5430 5680
rect -3500 8820 -3230 8950
rect -3500 8740 -3480 8820
rect -3400 8740 -3330 8820
rect -3250 8740 -3230 8820
rect -3500 8280 -3230 8740
rect -3500 8200 -3480 8280
rect -3400 8200 -3330 8280
rect -3250 8200 -3230 8280
rect -3500 7740 -3230 8200
rect -3500 7660 -3480 7740
rect -3400 7660 -3330 7740
rect -3250 7660 -3230 7740
rect -3500 2510 -3230 7660
rect -1010 8820 -740 9000
rect -1010 8740 -990 8820
rect -910 8740 -840 8820
rect -760 8740 -740 8820
rect -1010 8280 -740 8740
rect -1010 8200 -990 8280
rect -910 8200 -840 8280
rect -760 8200 -740 8280
rect -1010 7740 -740 8200
rect -1010 7660 -990 7740
rect -910 7660 -840 7740
rect -760 7660 -740 7740
rect -2210 7140 -1980 7160
rect -2210 7060 -2190 7140
rect -2110 7060 -2080 7140
rect -2000 7060 -1980 7140
rect -2210 6530 -1980 7060
rect -2210 6450 -2190 6530
rect -2110 6450 -2080 6530
rect -2000 6450 -1980 6530
rect -2210 5970 -1980 6450
rect -2210 5890 -2190 5970
rect -2110 5890 -2080 5970
rect -2000 5890 -1980 5970
rect -2210 3270 -1980 5890
rect -2210 3190 -2190 3270
rect -2110 3190 -2080 3270
rect -2000 3190 -1980 3270
rect -2210 3170 -1980 3190
rect -3500 2430 -3480 2510
rect -3400 2430 -3330 2510
rect -3250 2430 -3230 2510
rect -1010 2530 -740 7660
rect 1470 8820 1740 9010
rect 1470 8740 1490 8820
rect 1570 8740 1640 8820
rect 1720 8740 1740 8820
rect 1470 8280 1740 8740
rect 1470 8200 1490 8280
rect 1570 8200 1640 8280
rect 1720 8200 1740 8280
rect 1470 7740 1740 8200
rect 1470 7660 1500 7740
rect 1580 7660 1640 7740
rect 1720 7660 1740 7740
rect 200 7140 430 7160
rect 200 7060 220 7140
rect 300 7060 330 7140
rect 410 7060 430 7140
rect 200 6550 430 7060
rect 200 6470 220 6550
rect 300 6470 330 6550
rect 410 6470 430 6550
rect 200 5970 430 6470
rect 200 5890 220 5970
rect 300 5890 330 5970
rect 410 5890 430 5970
rect 200 3270 430 5890
rect 200 3190 220 3270
rect 300 3190 330 3270
rect 410 3190 430 3270
rect 200 3170 430 3190
rect -1010 2450 -990 2530
rect -910 2450 -840 2530
rect -760 2450 -740 2530
rect -1010 2430 -740 2450
rect 1470 2530 1740 7660
rect 2660 7130 2890 7170
rect 2660 7050 2680 7130
rect 2760 7050 2790 7130
rect 2870 7050 2890 7130
rect 2660 6550 2890 7050
rect 2660 6470 2680 6550
rect 2760 6470 2790 6550
rect 2870 6470 2890 6550
rect 2660 5970 2890 6470
rect 2660 5890 2680 5970
rect 2760 5890 2790 5970
rect 2870 5890 2890 5970
rect 2660 3280 2890 5890
rect 4210 5740 4500 9400
rect 4210 5660 4230 5740
rect 4310 5660 4400 5740
rect 4480 5660 4500 5740
rect 4210 5250 4500 5660
rect 2660 3200 2680 3280
rect 2760 3200 2790 3280
rect 2870 3200 2890 3280
rect 2660 3180 2890 3200
rect 1470 2450 1490 2530
rect 1570 2450 1630 2530
rect 1710 2450 1740 2530
rect 1470 2430 1740 2450
rect -3500 2400 -3230 2430
rect 1819 580 1941 581
rect 1819 480 1820 580
rect 1940 480 1941 580
rect 1819 479 1941 480
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_0
timestamp 1683391037
transform 0 -1 5700 1 0 11330
box -1750 -1700 1749 1700
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_1
timestamp 1683391037
transform 0 -1 -1900 1 0 11330
box -1750 -1700 1749 1700
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_2
timestamp 1683391037
transform 0 -1 1900 1 0 11330
box -1750 -1700 1749 1700
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_3
timestamp 1683391037
transform 0 -1 -5700 1 0 11330
box -1750 -1700 1749 1700
use sky130_fd_pr__nfet_01v8_GG6QWW  sky130_fd_pr__nfet_01v8_GG6QWW_0
timestamp 1683391037
transform 0 1 -5 -1 0 1436
box -296 -3755 296 3755
use sky130_fd_pr__nfet_01v8_GG6QWW  sky130_fd_pr__nfet_01v8_GG6QWW_1
timestamp 1683391037
transform 0 1 -5 -1 0 2056
box -296 -3755 296 3755
use sky130_fd_pr__nfet_01v8_K6FQWW  sky130_fd_pr__nfet_01v8_K6FQWW_0
timestamp 1683391037
transform 0 1 44 -1 0 2606
box -246 -4364 246 4364
use sky130_fd_pr__nfet_01v8_KG6QWW  sky130_fd_pr__nfet_01v8_KG6QWW_0
timestamp 1683391037
transform 0 1 44 -1 0 236
box -296 -4364 296 4364
use sky130_fd_pr__nfet_01v8_KG6QWW  sky130_fd_pr__nfet_01v8_KG6QWW_1
timestamp 1683391037
transform 0 1 44 -1 0 836
box -296 -4364 296 4364
use sky130_fd_pr__nfet_01v8_R8BLL7  sky130_fd_pr__nfet_01v8_R8BLL7_0
timestamp 1683391037
transform 0 1 44 -1 0 3106
box -246 -4364 246 4364
use sky130_fd_pr__pfet_01v8_SDAUVS  sky130_fd_pr__pfet_01v8_SDAUVS_0
timestamp 1683391037
transform 0 1 21 -1 0 3886
box -246 -6281 246 6281
use sky130_fd_pr__pfet_01v8_SDAUVS  sky130_fd_pr__pfet_01v8_SDAUVS_1
timestamp 1683391037
transform 0 1 21 -1 0 4426
box -246 -6281 246 6281
use sky130_fd_pr__pfet_01v8_SDAUVS  sky130_fd_pr__pfet_01v8_SDAUVS_2
timestamp 1683391037
transform 0 1 21 -1 0 5506
box -246 -6281 246 6281
use sky130_fd_pr__pfet_01v8_SDAUVS  sky130_fd_pr__pfet_01v8_SDAUVS_3
timestamp 1683391037
transform 0 1 21 -1 0 4966
box -246 -6281 246 6281
use sky130_fd_pr__pfet_01v8_T9YF2H  sky130_fd_pr__pfet_01v8_T9YF2H_0
timestamp 1683391037
transform 0 1 7 -1 0 6046
box -246 -4427 246 4427
use sky130_fd_pr__pfet_01v8_T9YF2H  sky130_fd_pr__pfet_01v8_T9YF2H_1
timestamp 1683391037
transform 0 1 7 -1 0 7746
box -246 -4427 246 4427
use sky130_fd_pr__pfet_01v8_T9YF2H  sky130_fd_pr__pfet_01v8_T9YF2H_2
timestamp 1683391037
transform 0 1 7 -1 0 6626
box -246 -4427 246 4427
use sky130_fd_pr__pfet_01v8_T9YF2H  sky130_fd_pr__pfet_01v8_T9YF2H_3
timestamp 1683391037
transform 0 1 7 -1 0 8286
box -246 -4427 246 4427
use sky130_fd_pr__pfet_01v8_T9YF2H  sky130_fd_pr__pfet_01v8_T9YF2H_4
timestamp 1683391037
transform 0 1 7 -1 0 8826
box -246 -4427 246 4427
use sky130_fd_pr__pfet_01v8_T9YF2H  sky130_fd_pr__pfet_01v8_T9YF2H_5
timestamp 1683391037
transform 0 1 7 -1 0 7206
box -246 -4427 246 4427
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_0
timestamp 1683391037
transform 0 1 8645 -1 0 4066
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_1
timestamp 1683391037
transform 0 1 8645 -1 0 5536
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_2
timestamp 1683391037
transform 0 1 -8415 -1 0 4066
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_3
timestamp 1683391037
transform 0 1 -8415 -1 0 5536
box -739 -1598 739 1598
<< end >>
