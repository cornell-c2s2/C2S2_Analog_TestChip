magic
tech sky130A
magscale 1 2
timestamp 1676504078
<< nwell >>
rect -7685 1941 7570 5876
<< pwell >>
rect -835 1575 240 1625
<< metal1 >>
rect -4160 7050 4160 7060
rect -4160 6990 -3820 7050
rect -3750 6990 -3660 7050
rect -3590 6990 -190 7050
rect -120 6990 -30 7050
rect 40 6990 3590 7050
rect 3660 6990 3750 7050
rect 3820 6990 4160 7050
rect -4250 6890 4260 6920
rect -4250 6860 2220 6890
rect -4250 6790 -2580 6860
rect -2510 6790 -2440 6860
rect -2370 6820 2220 6860
rect 2290 6820 2380 6890
rect 2450 6820 4260 6890
rect -2370 6790 4260 6820
rect -4250 6750 4260 6790
rect -4250 6680 -1380 6750
rect -1310 6680 -1220 6750
rect -1150 6740 4260 6750
rect -1150 6680 1050 6740
rect -4250 6670 1050 6680
rect 1120 6670 1210 6740
rect 1280 6670 4260 6740
rect -4250 6660 4260 6670
rect -4160 6450 4160 6465
rect -4160 6385 -3820 6450
rect -3750 6385 -3660 6450
rect -3590 6385 -190 6450
rect -120 6385 -30 6450
rect 40 6385 3590 6450
rect 3660 6385 3750 6450
rect 3820 6385 4160 6450
rect -4460 6300 4250 6310
rect -4460 6260 2220 6300
rect -4460 6190 -2570 6260
rect -2500 6190 -2440 6260
rect -2370 6230 2220 6260
rect 2290 6230 2380 6300
rect 2450 6230 4250 6300
rect -2370 6190 4250 6230
rect -4460 6120 -4440 6190
rect -4370 6120 -4300 6190
rect -4230 6160 4250 6190
rect -4230 6140 -770 6160
rect -4230 6120 -1380 6140
rect -4460 6070 -1380 6120
rect -1310 6070 -1220 6140
rect -1150 6090 -770 6140
rect -700 6090 -630 6160
rect -560 6140 4250 6160
rect -560 6130 2970 6140
rect -560 6090 1050 6130
rect -1150 6070 1050 6090
rect -4460 6060 1050 6070
rect 1120 6060 1210 6130
rect 1280 6070 2970 6130
rect 3040 6070 3110 6140
rect 3180 6070 4250 6140
rect 1280 6060 4250 6070
rect -4460 6050 4250 6060
rect -6060 5770 6970 5780
rect -6060 5750 6710 5770
rect -6060 5690 -4440 5750
rect -4370 5690 -4300 5750
rect -4230 5690 -770 5750
rect -700 5690 -630 5750
rect -560 5740 6710 5750
rect -560 5690 2970 5740
rect 3040 5690 3110 5740
rect 3180 5700 6710 5740
rect 6780 5700 6850 5770
rect 6920 5700 6970 5770
rect 3180 5690 6970 5700
rect -6150 5540 -5680 5610
rect -5610 5540 -5540 5610
rect -5470 5540 -2000 5610
rect -1930 5540 -1860 5610
rect -1790 5600 6150 5610
rect -1790 5540 1640 5600
rect -6150 5530 1640 5540
rect 1710 5530 1780 5600
rect 1850 5530 5470 5600
rect 5540 5530 5610 5600
rect 5680 5530 6150 5600
rect -6990 5430 -6710 5480
rect -6990 5360 -6950 5430
rect -6880 5360 -6810 5430
rect -6740 5370 -3260 5430
rect -3190 5370 -3120 5430
rect -3050 5370 500 5430
rect 570 5370 640 5430
rect 710 5380 4210 5430
rect 4280 5380 4350 5430
rect 4420 5380 6070 5430
rect 710 5370 6070 5380
rect -6740 5360 6070 5370
rect -6990 5330 -6710 5360
rect -7290 5060 7330 5070
rect -7290 4990 -4440 5060
rect -4370 4990 -4300 5060
rect -4230 4990 -770 5060
rect -700 4990 -630 5060
rect -560 5040 6710 5060
rect -560 4990 2970 5040
rect 3040 4990 3110 5040
rect 3180 4990 6710 5040
rect 6780 4990 6850 5060
rect 6920 4990 7330 5060
rect 6680 4970 6760 4990
rect 6810 4970 6890 4990
rect -7390 4820 -5680 4890
rect -5610 4820 -5540 4890
rect -5470 4820 -2000 4890
rect -1930 4820 -1860 4890
rect -1790 4880 7400 4890
rect -1790 4820 1640 4880
rect -7390 4810 1640 4820
rect 1710 4810 1780 4880
rect 1850 4810 5470 4880
rect 5540 4810 5610 4880
rect 5680 4810 7400 4880
rect -7300 4670 -6950 4730
rect -6880 4670 -6810 4730
rect -6740 4670 -3260 4730
rect -7300 4660 -3260 4670
rect -3190 4660 -3120 4730
rect -3050 4670 500 4730
rect 570 4670 640 4730
rect 710 4680 4210 4730
rect 4280 4680 4350 4730
rect 4420 4680 7320 4730
rect 710 4670 7320 4680
rect -3050 4660 7320 4670
rect -7300 4650 7320 4660
rect -7300 4360 7320 4370
rect -7300 4290 -4440 4360
rect -4370 4290 -4300 4360
rect -4230 4290 -770 4360
rect -700 4290 -630 4360
rect -560 4350 7320 4360
rect -560 4340 6710 4350
rect -560 4290 2970 4340
rect 3040 4290 3110 4340
rect 3180 4290 6710 4340
rect 6680 4280 6710 4290
rect 6780 4290 6850 4350
rect 6830 4280 6850 4290
rect 6920 4290 7320 4350
rect 6680 4270 6760 4280
rect 6830 4270 6910 4280
rect -7380 4140 -5680 4210
rect -5610 4140 -5540 4210
rect -5470 4140 -2000 4210
rect -1930 4140 -1860 4210
rect -1790 4200 7410 4210
rect -1790 4140 1640 4200
rect -7380 4130 1640 4140
rect 1710 4130 1780 4200
rect 1850 4130 5470 4200
rect 5540 4130 5610 4200
rect 5680 4130 7410 4200
rect -7300 3970 -6950 4030
rect -6880 3970 -6810 4030
rect -6740 3970 -3260 4030
rect -7300 3960 -3260 3970
rect -3190 3960 -3120 4030
rect -3050 3970 500 4030
rect 570 3970 640 4030
rect 710 3980 4210 4030
rect 4280 3980 4350 4030
rect 4420 3980 7320 4030
rect 710 3970 7320 3980
rect -3050 3960 7320 3970
rect -7300 3950 7320 3960
rect -7300 3620 7320 3640
rect -7300 3560 -4440 3620
rect -4370 3560 -4300 3620
rect -4230 3560 -770 3620
rect -700 3560 -630 3620
rect -560 3610 6710 3620
rect -560 3560 2970 3610
rect 3040 3560 3110 3610
rect 3180 3560 6710 3610
rect 6780 3560 6850 3620
rect 6920 3560 7320 3620
rect -7400 3460 7390 3470
rect -7400 3390 -5680 3460
rect -5610 3390 -5540 3460
rect -5470 3390 -2000 3460
rect -1930 3390 -1860 3460
rect -1790 3390 1640 3460
rect 1710 3390 1770 3460
rect 1840 3390 5470 3460
rect 5540 3390 5610 3460
rect 5680 3390 7390 3460
rect -7400 3380 7390 3390
rect -7310 3240 -6950 3300
rect -6880 3240 -6810 3300
rect -6740 3240 -3260 3300
rect -7310 3230 -3260 3240
rect -3190 3230 -3120 3300
rect -3050 3240 500 3300
rect 570 3240 640 3300
rect 710 3250 4210 3300
rect 4280 3250 4350 3300
rect 4420 3250 7310 3300
rect 710 3240 7310 3250
rect -3050 3230 7310 3240
rect -7310 3220 7310 3230
rect -3590 2960 3600 3030
rect -3690 2860 3670 2870
rect -3690 2790 -1720 2860
rect -1650 2790 -1500 2860
rect -1430 2790 1460 2860
rect 1530 2790 1700 2860
rect 1770 2790 3670 2860
rect -3690 2782 3670 2790
rect -3696 2634 3688 2782
rect -3600 2630 3590 2634
rect -3590 2370 3580 2450
rect -3680 2270 3676 2280
rect -3680 2200 -1720 2270
rect -1650 2200 -1500 2270
rect -1430 2200 1460 2270
rect 1530 2200 1700 2270
rect 1770 2200 3676 2270
rect -3680 2190 3676 2200
rect -3600 2040 -560 2110
rect -490 2040 -450 2110
rect -380 2040 380 2110
rect 450 2040 490 2110
rect 560 2040 3570 2110
rect -3600 2030 3570 2040
rect -920 1550 900 1620
rect -920 1540 380 1550
rect -920 1470 -560 1540
rect -490 1470 -450 1540
rect -380 1480 380 1540
rect 450 1480 490 1550
rect 560 1480 900 1550
rect -380 1470 900 1480
rect -900 1390 900 1470
rect -550 1350 -390 1390
rect -80 1350 75 1390
rect 390 1350 545 1390
rect -840 1265 830 1320
rect 1440 1030 1790 1050
rect -1740 1010 1460 1030
rect -1740 940 -1720 1010
rect -1650 940 -1510 1010
rect -1440 960 1460 1010
rect 1530 960 1700 1030
rect 1770 960 1790 1030
rect -1440 940 1790 960
rect -1740 920 1460 940
rect -1740 850 -1720 920
rect -1650 850 -1510 920
rect -1440 870 1460 920
rect 1530 870 1700 940
rect 1770 870 1790 940
rect -1440 850 1790 870
rect -1740 820 -1410 850
rect -615 790 620 795
rect -615 780 -560 790
rect -620 720 -560 780
rect -490 720 -450 790
rect -380 720 380 790
rect 450 720 490 790
rect 560 780 620 790
rect 560 720 630 780
rect -620 710 630 720
rect -3550 490 3540 495
rect -3550 420 -1720 490
rect -1650 420 -1500 490
rect -1430 420 1460 490
rect 1530 420 1700 490
rect 1770 420 3540 490
rect -3620 340 3615 345
rect -3620 270 -560 340
rect -490 270 -450 340
rect -380 270 380 340
rect 450 270 490 340
rect 560 270 3615 340
rect -3620 260 3615 270
rect -3550 95 3540 170
rect -2060 -290 -1830 95
rect -750 -290 -520 95
rect 530 -290 760 95
rect 1790 -290 2020 95
rect -2500 -720 2540 -290
rect -2500 -11670 2540 -11240
<< via1 >>
rect -3820 6980 -3750 7050
rect -3660 6980 -3590 7050
rect -190 6980 -120 7050
rect -30 6980 40 7050
rect 3590 6980 3660 7050
rect 3750 6980 3820 7050
rect -2580 6790 -2510 6860
rect -2440 6790 -2370 6860
rect 2220 6820 2290 6890
rect 2380 6820 2450 6890
rect -1380 6680 -1310 6750
rect -1220 6680 -1150 6750
rect 1050 6670 1120 6740
rect 1210 6670 1280 6740
rect -3820 6380 -3750 6450
rect -3660 6380 -3590 6450
rect -190 6380 -120 6450
rect -30 6380 40 6450
rect 3590 6380 3660 6450
rect 3750 6380 3820 6450
rect -2570 6190 -2500 6260
rect -2440 6190 -2370 6260
rect 2220 6230 2290 6300
rect 2380 6230 2450 6300
rect -4440 6120 -4370 6190
rect -4300 6120 -4230 6190
rect -1380 6070 -1310 6140
rect -1220 6070 -1150 6140
rect -770 6090 -700 6160
rect -630 6090 -560 6160
rect 1050 6060 1120 6130
rect 1210 6060 1280 6130
rect 2970 6070 3040 6140
rect 3110 6070 3180 6140
rect -4440 5680 -4370 5750
rect -4300 5680 -4230 5750
rect -770 5680 -700 5750
rect -630 5680 -560 5750
rect 2970 5670 3040 5740
rect 3110 5670 3180 5740
rect 6710 5700 6780 5770
rect 6850 5700 6920 5770
rect -5680 5540 -5610 5610
rect -5540 5540 -5470 5610
rect -2000 5540 -1930 5610
rect -1860 5540 -1790 5610
rect 1640 5530 1710 5600
rect 1780 5530 1850 5600
rect 5470 5530 5540 5600
rect 5610 5530 5680 5600
rect -6950 5360 -6880 5430
rect -6810 5360 -6740 5430
rect -3260 5370 -3190 5440
rect -3120 5370 -3050 5440
rect 500 5370 570 5440
rect 640 5370 710 5440
rect 4210 5380 4280 5450
rect 4350 5380 4420 5450
rect -4440 4990 -4370 5060
rect -4300 4990 -4230 5060
rect -770 4990 -700 5060
rect -630 4990 -560 5060
rect 2970 4970 3040 5040
rect 3110 4970 3180 5040
rect 6710 4990 6780 5060
rect 6850 4990 6920 5060
rect -5680 4820 -5610 4890
rect -5540 4820 -5470 4890
rect -2000 4820 -1930 4890
rect -1860 4820 -1790 4890
rect 1640 4810 1710 4880
rect 1780 4810 1850 4880
rect 5470 4810 5540 4880
rect 5610 4810 5680 4880
rect -6950 4670 -6880 4740
rect -6810 4670 -6740 4740
rect -3260 4660 -3190 4730
rect -3120 4660 -3050 4730
rect 500 4670 570 4740
rect 640 4670 710 4740
rect 4210 4680 4280 4750
rect 4350 4680 4420 4750
rect -4440 4290 -4370 4360
rect -4300 4290 -4230 4360
rect -770 4290 -700 4360
rect -630 4290 -560 4360
rect 2970 4270 3040 4340
rect 3110 4270 3180 4340
rect 6710 4280 6780 4350
rect 6850 4280 6920 4350
rect -5680 4140 -5610 4210
rect -5540 4140 -5470 4210
rect -2000 4140 -1930 4210
rect -1860 4140 -1790 4210
rect 1640 4130 1710 4200
rect 1780 4130 1850 4200
rect 5470 4130 5540 4200
rect 5610 4130 5680 4200
rect -6950 3970 -6880 4040
rect -6810 3970 -6740 4040
rect -3260 3960 -3190 4030
rect -3120 3960 -3050 4030
rect 500 3970 570 4040
rect 640 3970 710 4040
rect 4210 3980 4280 4050
rect 4350 3980 4420 4050
rect -4440 3550 -4370 3620
rect -4300 3550 -4230 3620
rect -770 3550 -700 3620
rect -630 3550 -560 3620
rect 2970 3540 3040 3610
rect 3110 3540 3180 3610
rect 6710 3550 6780 3620
rect 6850 3550 6920 3620
rect -5680 3390 -5610 3460
rect -5540 3390 -5470 3460
rect -2000 3390 -1930 3460
rect -1860 3390 -1790 3460
rect 1640 3390 1710 3460
rect 1770 3390 1840 3460
rect 5470 3390 5540 3460
rect 5610 3390 5680 3460
rect -6950 3240 -6880 3310
rect -6810 3240 -6740 3310
rect -3260 3230 -3190 3300
rect -3120 3230 -3050 3300
rect 500 3240 570 3310
rect 640 3240 710 3310
rect 4210 3250 4280 3320
rect 4350 3250 4420 3320
rect -1720 2790 -1650 2860
rect -1500 2790 -1430 2860
rect 1460 2790 1530 2860
rect 1700 2790 1770 2860
rect -1720 2200 -1650 2270
rect -1500 2200 -1430 2270
rect 1460 2200 1530 2270
rect 1700 2200 1770 2270
rect -560 2040 -490 2110
rect -450 2040 -380 2110
rect 380 2040 450 2110
rect 490 2040 560 2110
rect -560 1470 -490 1540
rect -450 1470 -380 1540
rect 380 1480 450 1550
rect 490 1480 560 1550
rect -1720 940 -1650 1010
rect -1510 940 -1440 1010
rect 1460 960 1530 1030
rect 1700 960 1770 1030
rect -1720 850 -1650 920
rect -1510 850 -1440 920
rect 1460 870 1530 940
rect 1700 870 1770 940
rect -560 720 -490 790
rect -450 720 -380 790
rect 380 720 450 790
rect 490 720 560 790
rect -1720 420 -1650 490
rect -1500 420 -1430 490
rect 1460 420 1530 490
rect 1700 420 1770 490
rect -560 270 -490 340
rect -450 270 -380 340
rect 380 270 450 340
rect 490 270 560 340
<< metal2 >>
rect -3840 7050 -3570 7060
rect -3840 6980 -3820 7050
rect -3750 6980 -3660 7050
rect -3590 6980 -3570 7050
rect -3840 6450 -3570 6980
rect -3840 6380 -3820 6450
rect -3750 6380 -3660 6450
rect -3590 6380 -3570 6450
rect -4460 6190 -4210 6310
rect -4460 6120 -4440 6190
rect -4370 6120 -4300 6190
rect -4230 6120 -4210 6190
rect -5700 5610 -5450 5780
rect -5700 5540 -5680 5610
rect -5610 5540 -5540 5610
rect -5470 5540 -5450 5610
rect -6970 5430 -6720 5480
rect -6970 5360 -6950 5430
rect -6880 5360 -6810 5430
rect -6740 5360 -6720 5430
rect -6970 4740 -6720 5360
rect -6970 4670 -6950 4740
rect -6880 4670 -6810 4740
rect -6740 4670 -6720 4740
rect -6970 4040 -6720 4670
rect -6970 3970 -6950 4040
rect -6880 3970 -6810 4040
rect -6740 3970 -6720 4040
rect -6970 3310 -6720 3970
rect -6970 3240 -6950 3310
rect -6880 3240 -6810 3310
rect -6740 3240 -6720 3310
rect -6970 3220 -6720 3240
rect -5700 4890 -5450 5540
rect -5700 4820 -5680 4890
rect -5610 4820 -5540 4890
rect -5470 4820 -5450 4890
rect -5700 4210 -5450 4820
rect -5700 4140 -5680 4210
rect -5610 4140 -5540 4210
rect -5470 4140 -5450 4210
rect -5700 3460 -5450 4140
rect -5700 3390 -5680 3460
rect -5610 3390 -5540 3460
rect -5470 3390 -5450 3460
rect -5700 3220 -5450 3390
rect -4460 5750 -4210 6120
rect -3840 6050 -3570 6380
rect -2610 6860 -2340 7060
rect -2610 6790 -2580 6860
rect -2510 6790 -2440 6860
rect -2370 6790 -2340 6860
rect -2610 6260 -2340 6790
rect -2610 6190 -2570 6260
rect -2500 6190 -2440 6260
rect -2370 6190 -2340 6260
rect -2610 6050 -2340 6190
rect -1400 6750 -1130 7060
rect -1400 6680 -1380 6750
rect -1310 6680 -1220 6750
rect -1150 6680 -1130 6750
rect -1400 6140 -1130 6680
rect -210 7050 60 7070
rect -210 6980 -190 7050
rect -120 6980 -30 7050
rect 40 6980 60 7050
rect -210 6450 60 6980
rect -210 6380 -190 6450
rect -120 6380 -30 6450
rect 40 6380 60 6450
rect -1400 6070 -1380 6140
rect -1310 6070 -1220 6140
rect -1150 6070 -1130 6140
rect -1400 6050 -1130 6070
rect -790 6160 -540 6300
rect -790 6090 -770 6160
rect -700 6090 -630 6160
rect -560 6090 -540 6160
rect -4460 5680 -4440 5750
rect -4370 5680 -4300 5750
rect -4230 5680 -4210 5750
rect -4460 5060 -4210 5680
rect -4460 4990 -4440 5060
rect -4370 4990 -4300 5060
rect -4230 4990 -4210 5060
rect -4460 4360 -4210 4990
rect -4460 4290 -4440 4360
rect -4370 4290 -4300 4360
rect -4230 4290 -4210 4360
rect -4460 3620 -4210 4290
rect -4460 3550 -4440 3620
rect -4370 3550 -4300 3620
rect -4230 3550 -4210 3620
rect -4460 3230 -4210 3550
rect -3280 5440 -3030 5780
rect -3280 5370 -3260 5440
rect -3190 5370 -3120 5440
rect -3050 5370 -3030 5440
rect -3280 4730 -3030 5370
rect -3280 4660 -3260 4730
rect -3190 4660 -3120 4730
rect -3050 4660 -3030 4730
rect -3280 4030 -3030 4660
rect -3280 3960 -3260 4030
rect -3190 3960 -3120 4030
rect -3050 3960 -3030 4030
rect -3280 3300 -3030 3960
rect -3280 3230 -3260 3300
rect -3190 3230 -3120 3300
rect -3050 3230 -3030 3300
rect -3280 3220 -3030 3230
rect -2020 5610 -1770 5780
rect -2020 5540 -2000 5610
rect -1930 5540 -1860 5610
rect -1790 5540 -1770 5610
rect -2020 4890 -1770 5540
rect -2020 4820 -2000 4890
rect -1930 4820 -1860 4890
rect -1790 4820 -1770 4890
rect -2020 4210 -1770 4820
rect -2020 4140 -2000 4210
rect -1930 4140 -1860 4210
rect -1790 4140 -1770 4210
rect -2020 3460 -1770 4140
rect -2020 3390 -2000 3460
rect -1930 3390 -1860 3460
rect -1790 3390 -1770 3460
rect -2020 2860 -1770 3390
rect -790 5750 -540 6090
rect -210 6060 60 6380
rect 1030 6740 1300 7060
rect 3570 7050 3840 7060
rect 1030 6670 1050 6740
rect 1120 6670 1210 6740
rect 1280 6670 1300 6740
rect 1030 6130 1300 6670
rect 1030 6060 1050 6130
rect 1120 6060 1210 6130
rect 1280 6060 1300 6130
rect 1030 6050 1300 6060
rect 2200 6890 2470 7050
rect 2200 6820 2220 6890
rect 2290 6820 2380 6890
rect 2450 6820 2470 6890
rect 2200 6300 2470 6820
rect 2200 6230 2220 6300
rect 2290 6230 2380 6300
rect 2450 6230 2470 6300
rect 2200 6040 2470 6230
rect 3570 6980 3590 7050
rect 3660 6980 3750 7050
rect 3820 6980 3840 7050
rect 3570 6450 3840 6980
rect 3570 6380 3590 6450
rect 3660 6380 3750 6450
rect 3820 6380 3840 6450
rect 2950 6140 3200 6220
rect 2950 6070 2970 6140
rect 3040 6070 3110 6140
rect 3180 6070 3200 6140
rect -790 5680 -770 5750
rect -700 5680 -630 5750
rect -560 5680 -540 5750
rect -790 5060 -540 5680
rect -790 4990 -770 5060
rect -700 4990 -630 5060
rect -560 4990 -540 5060
rect -790 4360 -540 4990
rect -790 4290 -770 4360
rect -700 4290 -630 4360
rect -560 4290 -540 4360
rect -790 3620 -540 4290
rect -790 3550 -770 3620
rect -700 3550 -630 3620
rect -560 3550 -540 3620
rect -790 3210 -540 3550
rect 480 5440 730 5790
rect 480 5370 500 5440
rect 570 5370 640 5440
rect 710 5370 730 5440
rect 480 4740 730 5370
rect 480 4670 500 4740
rect 570 4670 640 4740
rect 710 4670 730 4740
rect 480 4040 730 4670
rect 480 3970 500 4040
rect 570 3970 640 4040
rect 710 3970 730 4040
rect 480 3310 730 3970
rect 480 3240 500 3310
rect 570 3240 640 3310
rect 710 3240 730 3310
rect 480 3220 730 3240
rect 1620 5600 1870 5790
rect 1620 5530 1640 5600
rect 1710 5530 1780 5600
rect 1850 5530 1870 5600
rect 1620 4880 1870 5530
rect 1620 4810 1640 4880
rect 1710 4810 1780 4880
rect 1850 4810 1870 4880
rect 1620 4200 1870 4810
rect 1620 4130 1640 4200
rect 1710 4130 1780 4200
rect 1850 4130 1870 4200
rect 1620 3460 1870 4130
rect 1620 3390 1640 3460
rect 1710 3390 1770 3460
rect 1840 3390 1870 3460
rect 1620 2870 1870 3390
rect 2950 5740 3200 6070
rect 3570 6050 3840 6380
rect 2950 5670 2970 5740
rect 3040 5670 3110 5740
rect 3180 5670 3200 5740
rect 2950 5040 3200 5670
rect 2950 4970 2970 5040
rect 3040 4970 3110 5040
rect 3180 4970 3200 5040
rect 2950 4340 3200 4970
rect 2950 4270 2970 4340
rect 3040 4270 3110 4340
rect 3180 4270 3200 4340
rect 2950 3610 3200 4270
rect 2950 3540 2970 3610
rect 3040 3540 3110 3610
rect 3180 3540 3200 3610
rect 2950 3260 3200 3540
rect 4190 5450 4440 5790
rect 4190 5380 4210 5450
rect 4280 5380 4350 5450
rect 4420 5380 4440 5450
rect 4190 4750 4440 5380
rect 4190 4680 4210 4750
rect 4280 4680 4350 4750
rect 4420 4680 4440 4750
rect 4190 4050 4440 4680
rect 4190 3980 4210 4050
rect 4280 3980 4350 4050
rect 4420 3980 4440 4050
rect 4190 3320 4440 3980
rect 4190 3250 4210 3320
rect 4280 3250 4350 3320
rect 4420 3250 4440 3320
rect 4190 3230 4440 3250
rect 5450 5600 5700 5780
rect 5450 5530 5470 5600
rect 5540 5530 5610 5600
rect 5680 5530 5700 5600
rect 5450 4880 5700 5530
rect 5450 4810 5470 4880
rect 5540 4810 5610 4880
rect 5680 4810 5700 4880
rect 5450 4200 5700 4810
rect 5450 4130 5470 4200
rect 5540 4130 5610 4200
rect 5680 4130 5700 4200
rect 5450 3460 5700 4130
rect 5450 3390 5470 3460
rect 5540 3390 5610 3460
rect 5680 3390 5700 3460
rect 5450 3220 5700 3390
rect 6690 5770 6940 5780
rect 6690 5700 6710 5770
rect 6780 5700 6850 5770
rect 6920 5700 6940 5770
rect 6690 5060 6940 5700
rect 6690 4990 6710 5060
rect 6780 4990 6850 5060
rect 6920 4990 6940 5060
rect 6690 4350 6940 4990
rect 6690 4280 6710 4350
rect 6780 4280 6850 4350
rect 6920 4280 6940 4350
rect 6690 3620 6940 4280
rect 6690 3550 6710 3620
rect 6780 3550 6850 3620
rect 6920 3550 6940 3620
rect 6690 3220 6940 3550
rect 1440 2860 1870 2870
rect -2020 2790 -1720 2860
rect -1650 2790 -1500 2860
rect -1430 2790 -1410 2860
rect -2020 2780 -1410 2790
rect -1740 2270 -1410 2780
rect -1740 2200 -1720 2270
rect -1650 2200 -1500 2270
rect -1430 2200 -1410 2270
rect -1740 1010 -1410 2200
rect 1440 2790 1460 2860
rect 1530 2790 1700 2860
rect 1770 2790 1870 2860
rect 1440 2780 1870 2790
rect 1440 2270 1790 2780
rect 1440 2200 1460 2270
rect 1530 2200 1700 2270
rect 1770 2200 1790 2270
rect -1740 940 -1720 1010
rect -1650 940 -1510 1010
rect -1440 940 -1410 1010
rect -1740 920 -1410 940
rect -1740 850 -1720 920
rect -1650 850 -1510 920
rect -1440 850 -1410 920
rect -1740 490 -1410 850
rect -1740 420 -1720 490
rect -1650 420 -1500 490
rect -1430 420 -1410 490
rect -1740 410 -1410 420
rect -580 2110 -360 2120
rect -580 2040 -560 2110
rect -490 2040 -450 2110
rect -380 2040 -360 2110
rect -580 1540 -360 2040
rect -580 1470 -560 1540
rect -490 1470 -450 1540
rect -380 1470 -360 1540
rect -580 790 -360 1470
rect -580 720 -560 790
rect -490 720 -450 790
rect -380 720 -360 790
rect -580 340 -360 720
rect -580 270 -560 340
rect -490 270 -450 340
rect -380 270 -360 340
rect -580 200 -360 270
rect 360 2110 580 2130
rect 360 2040 380 2110
rect 450 2040 490 2110
rect 560 2040 580 2110
rect 360 1550 580 2040
rect 360 1480 380 1550
rect 450 1480 490 1550
rect 560 1480 580 1550
rect 360 790 580 1480
rect 360 720 380 790
rect 450 720 490 790
rect 560 720 580 790
rect 360 340 580 720
rect 1440 1030 1790 2200
rect 1440 960 1460 1030
rect 1530 960 1700 1030
rect 1770 960 1790 1030
rect 1440 940 1790 960
rect 1440 870 1460 940
rect 1530 870 1700 940
rect 1770 870 1790 940
rect 1440 490 1790 870
rect 1440 420 1460 490
rect 1530 420 1700 490
rect 1770 420 1790 490
rect 1440 390 1790 420
rect 360 270 380 340
rect 450 270 490 340
rect 560 270 580 340
rect 360 210 580 270
use sky130_fd_pr__nfet_01v8_GG6QWW  sky130_fd_pr__nfet_01v8_GG6QWW_0
timestamp 1676503286
transform 0 1 0 -1 0 296
box -296 -3755 296 3755
use sky130_fd_pr__nfet_01v8_JTC45A  sky130_fd_pr__nfet_01v8_JTC45A_0
timestamp 1676503286
transform 0 1 -3 -1 0 1446
box -296 -1037 296 1037
use sky130_fd_pr__nfet_01v8_KG6QWW  sky130_fd_pr__nfet_01v8_KG6QWW_0
timestamp 1676134575
transform 0 1 1 -1 0 6258
box -296 -4364 296 4364
use sky130_fd_pr__nfet_01v8_KG6QWW  sky130_fd_pr__nfet_01v8_KG6QWW_1
timestamp 1676134575
transform 0 1 -1 -1 0 6861
box -296 -4364 296 4364
use sky130_fd_pr__nfet_01v8_N53VJN  sky130_fd_pr__nfet_01v8_N53VJN_0
timestamp 1676503286
transform 0 1 -1 -1 0 871
box -246 -819 246 819
use sky130_fd_pr__pfet_01v8_A3L74C  sky130_fd_pr__pfet_01v8_A3L74C_0
timestamp 1676503286
transform 0 1 -1 -1 0 3428
box -296 -7517 296 7517
use sky130_fd_pr__pfet_01v8_A3L74C  sky130_fd_pr__pfet_01v8_A3L74C_1
timestamp 1676503286
transform 0 1 2 -1 0 4161
box -296 -7517 296 7517
use sky130_fd_pr__pfet_01v8_A3L74C  sky130_fd_pr__pfet_01v8_A3L74C_2
timestamp 1676503286
transform 0 1 2 -1 0 4861
box -296 -7517 296 7517
use sky130_fd_pr__pfet_01v8_MKLXZC  sky130_fd_pr__pfet_01v8_MKLXZC_0
timestamp 1676503286
transform 0 1 -1 -1 0 2236
box -296 -3809 296 3809
use sky130_fd_pr__pfet_01v8_MKLXZC  sky130_fd_pr__pfet_01v8_MKLXZC_1
timestamp 1676503286
transform 0 1 -1 -1 0 2826
box -296 -3809 296 3809
use sky130_fd_pr__pfet_01v8_PKLTV8  sky130_fd_pr__pfet_01v8_PKLTV8_0
timestamp 1676133442
transform 0 1 3 -1 0 5558
box -296 -6281 296 6281
use sky130_fd_pr__res_xhigh_po_5p73_9YMCJE  sky130_fd_pr__res_xhigh_po_5p73_9YMCJE_0
timestamp 1676143463
transform -1 0 1970 0 -1 -5972
box -575 -5682 575 5682
use sky130_fd_pr__res_xhigh_po_5p73_9YMCJE  sky130_fd_pr__res_xhigh_po_5p73_9YMCJE_1
timestamp 1676143463
transform -1 0 660 0 -1 -5972
box -575 -5682 575 5682
use sky130_fd_pr__res_xhigh_po_5p73_9YMCJE  sky130_fd_pr__res_xhigh_po_5p73_9YMCJE_2
timestamp 1676143463
transform -1 0 -650 0 -1 -5978
box -575 -5682 575 5682
use sky130_fd_pr__res_xhigh_po_5p73_9YMCJE  sky130_fd_pr__res_xhigh_po_5p73_9YMCJE_3
timestamp 1676143463
transform -1 0 -1920 0 -1 -5978
box -575 -5682 575 5682
<< end >>
