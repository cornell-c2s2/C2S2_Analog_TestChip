magic
tech sky130A
magscale 1 2
timestamp 1676503286
<< pwell >>
rect -296 -3755 296 3755
<< nmos >>
rect -100 2545 100 3545
rect -100 1327 100 2327
rect -100 109 100 1109
rect -100 -1109 100 -109
rect -100 -2327 100 -1327
rect -100 -3545 100 -2545
<< ndiff >>
rect -158 3533 -100 3545
rect -158 2557 -146 3533
rect -112 2557 -100 3533
rect -158 2545 -100 2557
rect 100 3533 158 3545
rect 100 2557 112 3533
rect 146 2557 158 3533
rect 100 2545 158 2557
rect -158 2315 -100 2327
rect -158 1339 -146 2315
rect -112 1339 -100 2315
rect -158 1327 -100 1339
rect 100 2315 158 2327
rect 100 1339 112 2315
rect 146 1339 158 2315
rect 100 1327 158 1339
rect -158 1097 -100 1109
rect -158 121 -146 1097
rect -112 121 -100 1097
rect -158 109 -100 121
rect 100 1097 158 1109
rect 100 121 112 1097
rect 146 121 158 1097
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -1097 -146 -121
rect -112 -1097 -100 -121
rect -158 -1109 -100 -1097
rect 100 -121 158 -109
rect 100 -1097 112 -121
rect 146 -1097 158 -121
rect 100 -1109 158 -1097
rect -158 -1339 -100 -1327
rect -158 -2315 -146 -1339
rect -112 -2315 -100 -1339
rect -158 -2327 -100 -2315
rect 100 -1339 158 -1327
rect 100 -2315 112 -1339
rect 146 -2315 158 -1339
rect 100 -2327 158 -2315
rect -158 -2557 -100 -2545
rect -158 -3533 -146 -2557
rect -112 -3533 -100 -2557
rect -158 -3545 -100 -3533
rect 100 -2557 158 -2545
rect 100 -3533 112 -2557
rect 146 -3533 158 -2557
rect 100 -3545 158 -3533
<< ndiffc >>
rect -146 2557 -112 3533
rect 112 2557 146 3533
rect -146 1339 -112 2315
rect 112 1339 146 2315
rect -146 121 -112 1097
rect 112 121 146 1097
rect -146 -1097 -112 -121
rect 112 -1097 146 -121
rect -146 -2315 -112 -1339
rect 112 -2315 146 -1339
rect -146 -3533 -112 -2557
rect 112 -3533 146 -2557
<< psubdiff >>
rect -260 3685 -164 3719
rect 164 3685 260 3719
rect -260 3623 -226 3685
rect 226 3623 260 3685
rect -260 -3685 -226 -3623
rect 226 -3685 260 -3623
rect -260 -3719 -164 -3685
rect 164 -3719 260 -3685
<< psubdiffcont >>
rect -164 3685 164 3719
rect -260 -3623 -226 3623
rect 226 -3623 260 3623
rect -164 -3719 164 -3685
<< poly >>
rect -100 3617 100 3633
rect -100 3583 -84 3617
rect 84 3583 100 3617
rect -100 3545 100 3583
rect -100 2507 100 2545
rect -100 2473 -84 2507
rect 84 2473 100 2507
rect -100 2457 100 2473
rect -100 2399 100 2415
rect -100 2365 -84 2399
rect 84 2365 100 2399
rect -100 2327 100 2365
rect -100 1289 100 1327
rect -100 1255 -84 1289
rect 84 1255 100 1289
rect -100 1239 100 1255
rect -100 1181 100 1197
rect -100 1147 -84 1181
rect 84 1147 100 1181
rect -100 1109 100 1147
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -1147 100 -1109
rect -100 -1181 -84 -1147
rect 84 -1181 100 -1147
rect -100 -1197 100 -1181
rect -100 -1255 100 -1239
rect -100 -1289 -84 -1255
rect 84 -1289 100 -1255
rect -100 -1327 100 -1289
rect -100 -2365 100 -2327
rect -100 -2399 -84 -2365
rect 84 -2399 100 -2365
rect -100 -2415 100 -2399
rect -100 -2473 100 -2457
rect -100 -2507 -84 -2473
rect 84 -2507 100 -2473
rect -100 -2545 100 -2507
rect -100 -3583 100 -3545
rect -100 -3617 -84 -3583
rect 84 -3617 100 -3583
rect -100 -3633 100 -3617
<< polycont >>
rect -84 3583 84 3617
rect -84 2473 84 2507
rect -84 2365 84 2399
rect -84 1255 84 1289
rect -84 1147 84 1181
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1181 84 -1147
rect -84 -1289 84 -1255
rect -84 -2399 84 -2365
rect -84 -2507 84 -2473
rect -84 -3617 84 -3583
<< locali >>
rect -260 3685 -164 3719
rect 164 3685 260 3719
rect -260 3623 -226 3685
rect 226 3623 260 3685
rect -100 3583 -84 3617
rect 84 3583 100 3617
rect -146 3533 -112 3549
rect -146 2541 -112 2557
rect 112 3533 146 3549
rect 112 2541 146 2557
rect -100 2473 -84 2507
rect 84 2473 100 2507
rect -100 2365 -84 2399
rect 84 2365 100 2399
rect -146 2315 -112 2331
rect -146 1323 -112 1339
rect 112 2315 146 2331
rect 112 1323 146 1339
rect -100 1255 -84 1289
rect 84 1255 100 1289
rect -100 1147 -84 1181
rect 84 1147 100 1181
rect -146 1097 -112 1113
rect -146 105 -112 121
rect 112 1097 146 1113
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -1113 -112 -1097
rect 112 -121 146 -105
rect 112 -1113 146 -1097
rect -100 -1181 -84 -1147
rect 84 -1181 100 -1147
rect -100 -1289 -84 -1255
rect 84 -1289 100 -1255
rect -146 -1339 -112 -1323
rect -146 -2331 -112 -2315
rect 112 -1339 146 -1323
rect 112 -2331 146 -2315
rect -100 -2399 -84 -2365
rect 84 -2399 100 -2365
rect -100 -2507 -84 -2473
rect 84 -2507 100 -2473
rect -146 -2557 -112 -2541
rect -146 -3549 -112 -3533
rect 112 -2557 146 -2541
rect 112 -3549 146 -3533
rect -100 -3617 -84 -3583
rect 84 -3617 100 -3583
rect -260 -3685 -226 -3623
rect 226 -3685 260 -3623
rect -260 -3719 -164 -3685
rect 164 -3719 260 -3685
<< viali >>
rect -84 3583 84 3617
rect -146 2557 -112 3533
rect 112 2557 146 3533
rect -84 2473 84 2507
rect -84 2365 84 2399
rect -146 1339 -112 2315
rect 112 1339 146 2315
rect -84 1255 84 1289
rect -84 1147 84 1181
rect -146 121 -112 1097
rect 112 121 146 1097
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1097 -112 -121
rect 112 -1097 146 -121
rect -84 -1181 84 -1147
rect -84 -1289 84 -1255
rect -146 -2315 -112 -1339
rect 112 -2315 146 -1339
rect -84 -2399 84 -2365
rect -84 -2507 84 -2473
rect -146 -3533 -112 -2557
rect 112 -3533 146 -2557
rect -84 -3617 84 -3583
<< metal1 >>
rect -96 3617 96 3623
rect -96 3583 -84 3617
rect 84 3583 96 3617
rect -96 3577 96 3583
rect -152 3533 -106 3545
rect -152 2557 -146 3533
rect -112 2557 -106 3533
rect -152 2545 -106 2557
rect 106 3533 152 3545
rect 106 2557 112 3533
rect 146 2557 152 3533
rect 106 2545 152 2557
rect -96 2507 96 2513
rect -96 2473 -84 2507
rect 84 2473 96 2507
rect -96 2467 96 2473
rect -96 2399 96 2405
rect -96 2365 -84 2399
rect 84 2365 96 2399
rect -96 2359 96 2365
rect -152 2315 -106 2327
rect -152 1339 -146 2315
rect -112 1339 -106 2315
rect -152 1327 -106 1339
rect 106 2315 152 2327
rect 106 1339 112 2315
rect 146 1339 152 2315
rect 106 1327 152 1339
rect -96 1289 96 1295
rect -96 1255 -84 1289
rect 84 1255 96 1289
rect -96 1249 96 1255
rect -96 1181 96 1187
rect -96 1147 -84 1181
rect 84 1147 96 1181
rect -96 1141 96 1147
rect -152 1097 -106 1109
rect -152 121 -146 1097
rect -112 121 -106 1097
rect -152 109 -106 121
rect 106 1097 152 1109
rect 106 121 112 1097
rect 146 121 152 1097
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -1097 -146 -121
rect -112 -1097 -106 -121
rect -152 -1109 -106 -1097
rect 106 -121 152 -109
rect 106 -1097 112 -121
rect 146 -1097 152 -121
rect 106 -1109 152 -1097
rect -96 -1147 96 -1141
rect -96 -1181 -84 -1147
rect 84 -1181 96 -1147
rect -96 -1187 96 -1181
rect -96 -1255 96 -1249
rect -96 -1289 -84 -1255
rect 84 -1289 96 -1255
rect -96 -1295 96 -1289
rect -152 -1339 -106 -1327
rect -152 -2315 -146 -1339
rect -112 -2315 -106 -1339
rect -152 -2327 -106 -2315
rect 106 -1339 152 -1327
rect 106 -2315 112 -1339
rect 146 -2315 152 -1339
rect 106 -2327 152 -2315
rect -96 -2365 96 -2359
rect -96 -2399 -84 -2365
rect 84 -2399 96 -2365
rect -96 -2405 96 -2399
rect -96 -2473 96 -2467
rect -96 -2507 -84 -2473
rect 84 -2507 96 -2473
rect -96 -2513 96 -2507
rect -152 -2557 -106 -2545
rect -152 -3533 -146 -2557
rect -112 -3533 -106 -2557
rect -152 -3545 -106 -3533
rect 106 -2557 152 -2545
rect 106 -3533 112 -2557
rect 146 -3533 152 -2557
rect 106 -3545 152 -3533
rect -96 -3583 96 -3577
rect -96 -3617 -84 -3583
rect 84 -3617 96 -3583
rect -96 -3623 96 -3617
<< properties >>
string FIXED_BBOX -243 -3702 243 3702
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 1 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
