magic
tech sky130A
magscale 1 2
timestamp 1676503286
<< pwell >>
rect -246 -819 246 819
<< nmos >>
rect -50 109 50 609
rect -50 -609 50 -109
<< ndiff >>
rect -108 597 -50 609
rect -108 121 -96 597
rect -62 121 -50 597
rect -108 109 -50 121
rect 50 597 108 609
rect 50 121 62 597
rect 96 121 108 597
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -597 -96 -121
rect -62 -597 -50 -121
rect -108 -609 -50 -597
rect 50 -121 108 -109
rect 50 -597 62 -121
rect 96 -597 108 -121
rect 50 -609 108 -597
<< ndiffc >>
rect -96 121 -62 597
rect 62 121 96 597
rect -96 -597 -62 -121
rect 62 -597 96 -121
<< psubdiff >>
rect -210 749 -114 783
rect 114 749 210 783
rect -210 687 -176 749
rect 176 687 210 749
rect -210 -749 -176 -687
rect 176 -749 210 -687
rect -210 -783 -114 -749
rect 114 -783 210 -749
<< psubdiffcont >>
rect -114 749 114 783
rect -210 -687 -176 687
rect 176 -687 210 687
rect -114 -783 114 -749
<< poly >>
rect -50 681 50 697
rect -50 647 -34 681
rect 34 647 50 681
rect -50 609 50 647
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -647 50 -609
rect -50 -681 -34 -647
rect 34 -681 50 -647
rect -50 -697 50 -681
<< polycont >>
rect -34 647 34 681
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -681 34 -647
<< locali >>
rect -210 749 -114 783
rect 114 749 210 783
rect -210 687 -176 749
rect 176 687 210 749
rect -50 647 -34 681
rect 34 647 50 681
rect -96 597 -62 613
rect -96 105 -62 121
rect 62 597 96 613
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -613 -62 -597
rect 62 -121 96 -105
rect 62 -613 96 -597
rect -50 -681 -34 -647
rect 34 -681 50 -647
rect -210 -749 -176 -687
rect 176 -749 210 -687
rect -210 -783 -114 -749
rect 114 -783 210 -749
<< viali >>
rect -34 647 34 681
rect -96 121 -62 597
rect 62 121 96 597
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -597 -62 -121
rect 62 -597 96 -121
rect -34 -681 34 -647
<< metal1 >>
rect -46 681 46 687
rect -46 647 -34 681
rect 34 647 46 681
rect -46 641 46 647
rect -102 597 -56 609
rect -102 121 -96 597
rect -62 121 -56 597
rect -102 109 -56 121
rect 56 597 102 609
rect 56 121 62 597
rect 96 121 102 597
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -597 -96 -121
rect -62 -597 -56 -121
rect -102 -609 -56 -597
rect 56 -121 102 -109
rect 56 -597 62 -121
rect 96 -597 102 -121
rect 56 -609 102 -597
rect -46 -647 46 -641
rect -46 -681 -34 -647
rect 34 -681 46 -647
rect -46 -687 46 -681
<< properties >>
string FIXED_BBOX -193 -766 193 766
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l .5 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
