magic
tech sky130A
magscale 1 2
timestamp 1679679663
<< nwell >>
rect -3322 26510 3338 31260
rect -3840 18401 3830 19642
rect -3810 18400 3808 18401
<< pwell >>
rect -7300 30630 -4104 32108
rect 4118 31982 7294 32068
rect -7300 29130 -4104 30608
rect 4118 30696 4204 31982
rect 7208 30696 7294 31982
rect 4118 30610 7294 30696
rect 4118 30502 7294 30588
rect 4118 29216 4204 30502
rect 7208 29216 7294 30502
rect 4118 29130 7294 29216
rect -711 23340 709 26381
rect -1702 21820 1708 23340
rect -1962 20420 1964 21820
rect -1040 17610 1034 18202
rect -820 17085 818 17577
rect -3755 16460 3755 17052
rect -3290 10140 3290 15452
rect -3290 2638 3280 10140
<< nmos >>
rect -525 25181 -425 26181
rect -367 25181 -267 26181
rect -209 25181 -109 26181
rect -51 25181 49 26181
rect 107 25181 207 26181
rect 265 25181 365 26181
rect 423 25181 523 26181
rect -525 23661 -425 24661
rect -367 23661 -267 24661
rect -209 23661 -109 24661
rect -51 23661 49 24661
rect 107 23661 207 24661
rect 265 23661 365 24661
rect 423 23661 523 24661
rect -1516 22140 -1316 23140
rect -1258 22140 -1058 23140
rect -1000 22140 -800 23140
rect -742 22140 -542 23140
rect -484 22140 -284 23140
rect -226 22140 -26 23140
rect 32 22140 232 23140
rect 290 22140 490 23140
rect 548 22140 748 23140
rect 806 22140 1006 23140
rect 1064 22140 1264 23140
rect 1322 22140 1522 23140
rect -1776 20620 -1576 21620
rect -1518 20620 -1318 21620
rect -1260 20620 -1060 21620
rect -1002 20620 -802 21620
rect -744 20620 -544 21620
rect -486 20620 -286 21620
rect -228 20620 -28 21620
rect 30 20620 230 21620
rect 288 20620 488 21620
rect 546 20620 746 21620
rect 804 20620 1004 21620
rect 1062 20620 1262 21620
rect 1320 20620 1520 21620
rect 1578 20620 1778 21620
rect -830 17806 -580 18006
rect -362 17806 -112 18006
rect 106 17806 356 18006
rect 574 17806 824 18006
rect -610 17281 -110 17381
rect 108 17281 608 17381
rect -3545 16656 -2545 16856
rect -2327 16656 -1327 16856
rect -1109 16656 -109 16856
rect 109 16656 1109 16856
rect 1327 16656 2327 16856
rect 2545 16656 3545 16856
<< pmos >>
rect -3126 29959 -3026 30959
rect -2968 29959 -2868 30959
rect -2810 29959 -2710 30959
rect -2652 29959 -2552 30959
rect -2494 29959 -2394 30959
rect -2336 29959 -2236 30959
rect -2178 29959 -2078 30959
rect -2020 29959 -1920 30959
rect -1862 29959 -1762 30959
rect -1704 29959 -1604 30959
rect -1546 29959 -1446 30959
rect -1388 29959 -1288 30959
rect -1230 29959 -1130 30959
rect -1072 29959 -972 30959
rect -914 29959 -814 30959
rect -756 29959 -656 30959
rect -598 29959 -498 30959
rect -440 29959 -340 30959
rect -282 29959 -182 30959
rect -124 29959 -24 30959
rect 34 29959 134 30959
rect 192 29959 292 30959
rect 350 29959 450 30959
rect 508 29959 608 30959
rect 666 29959 766 30959
rect 824 29959 924 30959
rect 982 29959 1082 30959
rect 1140 29959 1240 30959
rect 1298 29959 1398 30959
rect 1456 29959 1556 30959
rect 1614 29959 1714 30959
rect 1772 29959 1872 30959
rect 1930 29959 2030 30959
rect 2088 29959 2188 30959
rect 2246 29959 2346 30959
rect 2404 29959 2504 30959
rect 2562 29959 2662 30959
rect 2720 29959 2820 30959
rect 2878 29959 2978 30959
rect 3036 29959 3136 30959
rect -1626 28289 -1526 29289
rect -1468 28289 -1368 29289
rect -1310 28289 -1210 29289
rect -1152 28289 -1052 29289
rect -994 28289 -894 29289
rect -836 28289 -736 29289
rect -678 28289 -578 29289
rect -520 28289 -420 29289
rect -362 28289 -262 29289
rect -204 28289 -104 29289
rect -46 28289 54 29289
rect 112 28289 212 29289
rect 270 28289 370 29289
rect 428 28289 528 29289
rect 586 28289 686 29289
rect 744 28289 844 29289
rect 902 28289 1002 29289
rect 1060 28289 1160 29289
rect 1218 28289 1318 29289
rect 1376 28289 1476 29289
rect 1534 28289 1634 29289
rect -1626 26749 -1526 27749
rect -1468 26749 -1368 27749
rect -1310 26749 -1210 27749
rect -1152 26749 -1052 27749
rect -994 26749 -894 27749
rect -836 26749 -736 27749
rect -678 26749 -578 27749
rect -520 26749 -420 27749
rect -362 26749 -262 27749
rect -204 26749 -104 27749
rect -46 26749 54 27749
rect 112 26749 212 27749
rect 270 26749 370 27749
rect 428 26749 528 27749
rect 586 26749 686 27749
rect 744 26749 844 27749
rect 902 26749 1002 27749
rect 1060 26749 1160 27749
rect 1218 26749 1318 27749
rect 1376 26749 1476 27749
rect 1534 26749 1634 27749
rect -3591 19186 -2591 19386
rect -2355 19186 -1355 19386
rect -1119 19186 -119 19386
rect 117 19186 1117 19386
rect 1353 19186 2353 19386
rect 2589 19186 3589 19386
rect -3591 18596 -2591 18796
rect -2355 18596 -1355 18796
rect -1119 18596 -119 18796
rect 117 18596 1117 18796
rect 1353 18596 2353 18796
rect 2589 18596 3589 18796
<< ndiff >>
rect -583 26140 -525 26181
rect -583 26106 -571 26140
rect -537 26106 -525 26140
rect -583 26072 -525 26106
rect -583 26038 -571 26072
rect -537 26038 -525 26072
rect -583 26004 -525 26038
rect -583 25970 -571 26004
rect -537 25970 -525 26004
rect -583 25936 -525 25970
rect -583 25902 -571 25936
rect -537 25902 -525 25936
rect -583 25868 -525 25902
rect -583 25834 -571 25868
rect -537 25834 -525 25868
rect -583 25800 -525 25834
rect -583 25766 -571 25800
rect -537 25766 -525 25800
rect -583 25732 -525 25766
rect -583 25698 -571 25732
rect -537 25698 -525 25732
rect -583 25664 -525 25698
rect -583 25630 -571 25664
rect -537 25630 -525 25664
rect -583 25596 -525 25630
rect -583 25562 -571 25596
rect -537 25562 -525 25596
rect -583 25528 -525 25562
rect -583 25494 -571 25528
rect -537 25494 -525 25528
rect -583 25460 -525 25494
rect -583 25426 -571 25460
rect -537 25426 -525 25460
rect -583 25392 -525 25426
rect -583 25358 -571 25392
rect -537 25358 -525 25392
rect -583 25324 -525 25358
rect -583 25290 -571 25324
rect -537 25290 -525 25324
rect -583 25256 -525 25290
rect -583 25222 -571 25256
rect -537 25222 -525 25256
rect -583 25181 -525 25222
rect -425 26140 -367 26181
rect -425 26106 -413 26140
rect -379 26106 -367 26140
rect -425 26072 -367 26106
rect -425 26038 -413 26072
rect -379 26038 -367 26072
rect -425 26004 -367 26038
rect -425 25970 -413 26004
rect -379 25970 -367 26004
rect -425 25936 -367 25970
rect -425 25902 -413 25936
rect -379 25902 -367 25936
rect -425 25868 -367 25902
rect -425 25834 -413 25868
rect -379 25834 -367 25868
rect -425 25800 -367 25834
rect -425 25766 -413 25800
rect -379 25766 -367 25800
rect -425 25732 -367 25766
rect -425 25698 -413 25732
rect -379 25698 -367 25732
rect -425 25664 -367 25698
rect -425 25630 -413 25664
rect -379 25630 -367 25664
rect -425 25596 -367 25630
rect -425 25562 -413 25596
rect -379 25562 -367 25596
rect -425 25528 -367 25562
rect -425 25494 -413 25528
rect -379 25494 -367 25528
rect -425 25460 -367 25494
rect -425 25426 -413 25460
rect -379 25426 -367 25460
rect -425 25392 -367 25426
rect -425 25358 -413 25392
rect -379 25358 -367 25392
rect -425 25324 -367 25358
rect -425 25290 -413 25324
rect -379 25290 -367 25324
rect -425 25256 -367 25290
rect -425 25222 -413 25256
rect -379 25222 -367 25256
rect -425 25181 -367 25222
rect -267 26140 -209 26181
rect -267 26106 -255 26140
rect -221 26106 -209 26140
rect -267 26072 -209 26106
rect -267 26038 -255 26072
rect -221 26038 -209 26072
rect -267 26004 -209 26038
rect -267 25970 -255 26004
rect -221 25970 -209 26004
rect -267 25936 -209 25970
rect -267 25902 -255 25936
rect -221 25902 -209 25936
rect -267 25868 -209 25902
rect -267 25834 -255 25868
rect -221 25834 -209 25868
rect -267 25800 -209 25834
rect -267 25766 -255 25800
rect -221 25766 -209 25800
rect -267 25732 -209 25766
rect -267 25698 -255 25732
rect -221 25698 -209 25732
rect -267 25664 -209 25698
rect -267 25630 -255 25664
rect -221 25630 -209 25664
rect -267 25596 -209 25630
rect -267 25562 -255 25596
rect -221 25562 -209 25596
rect -267 25528 -209 25562
rect -267 25494 -255 25528
rect -221 25494 -209 25528
rect -267 25460 -209 25494
rect -267 25426 -255 25460
rect -221 25426 -209 25460
rect -267 25392 -209 25426
rect -267 25358 -255 25392
rect -221 25358 -209 25392
rect -267 25324 -209 25358
rect -267 25290 -255 25324
rect -221 25290 -209 25324
rect -267 25256 -209 25290
rect -267 25222 -255 25256
rect -221 25222 -209 25256
rect -267 25181 -209 25222
rect -109 26140 -51 26181
rect -109 26106 -97 26140
rect -63 26106 -51 26140
rect -109 26072 -51 26106
rect -109 26038 -97 26072
rect -63 26038 -51 26072
rect -109 26004 -51 26038
rect -109 25970 -97 26004
rect -63 25970 -51 26004
rect -109 25936 -51 25970
rect -109 25902 -97 25936
rect -63 25902 -51 25936
rect -109 25868 -51 25902
rect -109 25834 -97 25868
rect -63 25834 -51 25868
rect -109 25800 -51 25834
rect -109 25766 -97 25800
rect -63 25766 -51 25800
rect -109 25732 -51 25766
rect -109 25698 -97 25732
rect -63 25698 -51 25732
rect -109 25664 -51 25698
rect -109 25630 -97 25664
rect -63 25630 -51 25664
rect -109 25596 -51 25630
rect -109 25562 -97 25596
rect -63 25562 -51 25596
rect -109 25528 -51 25562
rect -109 25494 -97 25528
rect -63 25494 -51 25528
rect -109 25460 -51 25494
rect -109 25426 -97 25460
rect -63 25426 -51 25460
rect -109 25392 -51 25426
rect -109 25358 -97 25392
rect -63 25358 -51 25392
rect -109 25324 -51 25358
rect -109 25290 -97 25324
rect -63 25290 -51 25324
rect -109 25256 -51 25290
rect -109 25222 -97 25256
rect -63 25222 -51 25256
rect -109 25181 -51 25222
rect 49 26140 107 26181
rect 49 26106 61 26140
rect 95 26106 107 26140
rect 49 26072 107 26106
rect 49 26038 61 26072
rect 95 26038 107 26072
rect 49 26004 107 26038
rect 49 25970 61 26004
rect 95 25970 107 26004
rect 49 25936 107 25970
rect 49 25902 61 25936
rect 95 25902 107 25936
rect 49 25868 107 25902
rect 49 25834 61 25868
rect 95 25834 107 25868
rect 49 25800 107 25834
rect 49 25766 61 25800
rect 95 25766 107 25800
rect 49 25732 107 25766
rect 49 25698 61 25732
rect 95 25698 107 25732
rect 49 25664 107 25698
rect 49 25630 61 25664
rect 95 25630 107 25664
rect 49 25596 107 25630
rect 49 25562 61 25596
rect 95 25562 107 25596
rect 49 25528 107 25562
rect 49 25494 61 25528
rect 95 25494 107 25528
rect 49 25460 107 25494
rect 49 25426 61 25460
rect 95 25426 107 25460
rect 49 25392 107 25426
rect 49 25358 61 25392
rect 95 25358 107 25392
rect 49 25324 107 25358
rect 49 25290 61 25324
rect 95 25290 107 25324
rect 49 25256 107 25290
rect 49 25222 61 25256
rect 95 25222 107 25256
rect 49 25181 107 25222
rect 207 26140 265 26181
rect 207 26106 219 26140
rect 253 26106 265 26140
rect 207 26072 265 26106
rect 207 26038 219 26072
rect 253 26038 265 26072
rect 207 26004 265 26038
rect 207 25970 219 26004
rect 253 25970 265 26004
rect 207 25936 265 25970
rect 207 25902 219 25936
rect 253 25902 265 25936
rect 207 25868 265 25902
rect 207 25834 219 25868
rect 253 25834 265 25868
rect 207 25800 265 25834
rect 207 25766 219 25800
rect 253 25766 265 25800
rect 207 25732 265 25766
rect 207 25698 219 25732
rect 253 25698 265 25732
rect 207 25664 265 25698
rect 207 25630 219 25664
rect 253 25630 265 25664
rect 207 25596 265 25630
rect 207 25562 219 25596
rect 253 25562 265 25596
rect 207 25528 265 25562
rect 207 25494 219 25528
rect 253 25494 265 25528
rect 207 25460 265 25494
rect 207 25426 219 25460
rect 253 25426 265 25460
rect 207 25392 265 25426
rect 207 25358 219 25392
rect 253 25358 265 25392
rect 207 25324 265 25358
rect 207 25290 219 25324
rect 253 25290 265 25324
rect 207 25256 265 25290
rect 207 25222 219 25256
rect 253 25222 265 25256
rect 207 25181 265 25222
rect 365 26140 423 26181
rect 365 26106 377 26140
rect 411 26106 423 26140
rect 365 26072 423 26106
rect 365 26038 377 26072
rect 411 26038 423 26072
rect 365 26004 423 26038
rect 365 25970 377 26004
rect 411 25970 423 26004
rect 365 25936 423 25970
rect 365 25902 377 25936
rect 411 25902 423 25936
rect 365 25868 423 25902
rect 365 25834 377 25868
rect 411 25834 423 25868
rect 365 25800 423 25834
rect 365 25766 377 25800
rect 411 25766 423 25800
rect 365 25732 423 25766
rect 365 25698 377 25732
rect 411 25698 423 25732
rect 365 25664 423 25698
rect 365 25630 377 25664
rect 411 25630 423 25664
rect 365 25596 423 25630
rect 365 25562 377 25596
rect 411 25562 423 25596
rect 365 25528 423 25562
rect 365 25494 377 25528
rect 411 25494 423 25528
rect 365 25460 423 25494
rect 365 25426 377 25460
rect 411 25426 423 25460
rect 365 25392 423 25426
rect 365 25358 377 25392
rect 411 25358 423 25392
rect 365 25324 423 25358
rect 365 25290 377 25324
rect 411 25290 423 25324
rect 365 25256 423 25290
rect 365 25222 377 25256
rect 411 25222 423 25256
rect 365 25181 423 25222
rect 523 26140 581 26181
rect 523 26106 535 26140
rect 569 26106 581 26140
rect 523 26072 581 26106
rect 523 26038 535 26072
rect 569 26038 581 26072
rect 523 26004 581 26038
rect 523 25970 535 26004
rect 569 25970 581 26004
rect 523 25936 581 25970
rect 523 25902 535 25936
rect 569 25902 581 25936
rect 523 25868 581 25902
rect 523 25834 535 25868
rect 569 25834 581 25868
rect 523 25800 581 25834
rect 523 25766 535 25800
rect 569 25766 581 25800
rect 523 25732 581 25766
rect 523 25698 535 25732
rect 569 25698 581 25732
rect 523 25664 581 25698
rect 523 25630 535 25664
rect 569 25630 581 25664
rect 523 25596 581 25630
rect 523 25562 535 25596
rect 569 25562 581 25596
rect 523 25528 581 25562
rect 523 25494 535 25528
rect 569 25494 581 25528
rect 523 25460 581 25494
rect 523 25426 535 25460
rect 569 25426 581 25460
rect 523 25392 581 25426
rect 523 25358 535 25392
rect 569 25358 581 25392
rect 523 25324 581 25358
rect 523 25290 535 25324
rect 569 25290 581 25324
rect 523 25256 581 25290
rect 523 25222 535 25256
rect 569 25222 581 25256
rect 523 25181 581 25222
rect -583 24620 -525 24661
rect -583 24586 -571 24620
rect -537 24586 -525 24620
rect -583 24552 -525 24586
rect -583 24518 -571 24552
rect -537 24518 -525 24552
rect -583 24484 -525 24518
rect -583 24450 -571 24484
rect -537 24450 -525 24484
rect -583 24416 -525 24450
rect -583 24382 -571 24416
rect -537 24382 -525 24416
rect -583 24348 -525 24382
rect -583 24314 -571 24348
rect -537 24314 -525 24348
rect -583 24280 -525 24314
rect -583 24246 -571 24280
rect -537 24246 -525 24280
rect -583 24212 -525 24246
rect -583 24178 -571 24212
rect -537 24178 -525 24212
rect -583 24144 -525 24178
rect -583 24110 -571 24144
rect -537 24110 -525 24144
rect -583 24076 -525 24110
rect -583 24042 -571 24076
rect -537 24042 -525 24076
rect -583 24008 -525 24042
rect -583 23974 -571 24008
rect -537 23974 -525 24008
rect -583 23940 -525 23974
rect -583 23906 -571 23940
rect -537 23906 -525 23940
rect -583 23872 -525 23906
rect -583 23838 -571 23872
rect -537 23838 -525 23872
rect -583 23804 -525 23838
rect -583 23770 -571 23804
rect -537 23770 -525 23804
rect -583 23736 -525 23770
rect -583 23702 -571 23736
rect -537 23702 -525 23736
rect -583 23661 -525 23702
rect -425 24620 -367 24661
rect -425 24586 -413 24620
rect -379 24586 -367 24620
rect -425 24552 -367 24586
rect -425 24518 -413 24552
rect -379 24518 -367 24552
rect -425 24484 -367 24518
rect -425 24450 -413 24484
rect -379 24450 -367 24484
rect -425 24416 -367 24450
rect -425 24382 -413 24416
rect -379 24382 -367 24416
rect -425 24348 -367 24382
rect -425 24314 -413 24348
rect -379 24314 -367 24348
rect -425 24280 -367 24314
rect -425 24246 -413 24280
rect -379 24246 -367 24280
rect -425 24212 -367 24246
rect -425 24178 -413 24212
rect -379 24178 -367 24212
rect -425 24144 -367 24178
rect -425 24110 -413 24144
rect -379 24110 -367 24144
rect -425 24076 -367 24110
rect -425 24042 -413 24076
rect -379 24042 -367 24076
rect -425 24008 -367 24042
rect -425 23974 -413 24008
rect -379 23974 -367 24008
rect -425 23940 -367 23974
rect -425 23906 -413 23940
rect -379 23906 -367 23940
rect -425 23872 -367 23906
rect -425 23838 -413 23872
rect -379 23838 -367 23872
rect -425 23804 -367 23838
rect -425 23770 -413 23804
rect -379 23770 -367 23804
rect -425 23736 -367 23770
rect -425 23702 -413 23736
rect -379 23702 -367 23736
rect -425 23661 -367 23702
rect -267 24620 -209 24661
rect -267 24586 -255 24620
rect -221 24586 -209 24620
rect -267 24552 -209 24586
rect -267 24518 -255 24552
rect -221 24518 -209 24552
rect -267 24484 -209 24518
rect -267 24450 -255 24484
rect -221 24450 -209 24484
rect -267 24416 -209 24450
rect -267 24382 -255 24416
rect -221 24382 -209 24416
rect -267 24348 -209 24382
rect -267 24314 -255 24348
rect -221 24314 -209 24348
rect -267 24280 -209 24314
rect -267 24246 -255 24280
rect -221 24246 -209 24280
rect -267 24212 -209 24246
rect -267 24178 -255 24212
rect -221 24178 -209 24212
rect -267 24144 -209 24178
rect -267 24110 -255 24144
rect -221 24110 -209 24144
rect -267 24076 -209 24110
rect -267 24042 -255 24076
rect -221 24042 -209 24076
rect -267 24008 -209 24042
rect -267 23974 -255 24008
rect -221 23974 -209 24008
rect -267 23940 -209 23974
rect -267 23906 -255 23940
rect -221 23906 -209 23940
rect -267 23872 -209 23906
rect -267 23838 -255 23872
rect -221 23838 -209 23872
rect -267 23804 -209 23838
rect -267 23770 -255 23804
rect -221 23770 -209 23804
rect -267 23736 -209 23770
rect -267 23702 -255 23736
rect -221 23702 -209 23736
rect -267 23661 -209 23702
rect -109 24620 -51 24661
rect -109 24586 -97 24620
rect -63 24586 -51 24620
rect -109 24552 -51 24586
rect -109 24518 -97 24552
rect -63 24518 -51 24552
rect -109 24484 -51 24518
rect -109 24450 -97 24484
rect -63 24450 -51 24484
rect -109 24416 -51 24450
rect -109 24382 -97 24416
rect -63 24382 -51 24416
rect -109 24348 -51 24382
rect -109 24314 -97 24348
rect -63 24314 -51 24348
rect -109 24280 -51 24314
rect -109 24246 -97 24280
rect -63 24246 -51 24280
rect -109 24212 -51 24246
rect -109 24178 -97 24212
rect -63 24178 -51 24212
rect -109 24144 -51 24178
rect -109 24110 -97 24144
rect -63 24110 -51 24144
rect -109 24076 -51 24110
rect -109 24042 -97 24076
rect -63 24042 -51 24076
rect -109 24008 -51 24042
rect -109 23974 -97 24008
rect -63 23974 -51 24008
rect -109 23940 -51 23974
rect -109 23906 -97 23940
rect -63 23906 -51 23940
rect -109 23872 -51 23906
rect -109 23838 -97 23872
rect -63 23838 -51 23872
rect -109 23804 -51 23838
rect -109 23770 -97 23804
rect -63 23770 -51 23804
rect -109 23736 -51 23770
rect -109 23702 -97 23736
rect -63 23702 -51 23736
rect -109 23661 -51 23702
rect 49 24620 107 24661
rect 49 24586 61 24620
rect 95 24586 107 24620
rect 49 24552 107 24586
rect 49 24518 61 24552
rect 95 24518 107 24552
rect 49 24484 107 24518
rect 49 24450 61 24484
rect 95 24450 107 24484
rect 49 24416 107 24450
rect 49 24382 61 24416
rect 95 24382 107 24416
rect 49 24348 107 24382
rect 49 24314 61 24348
rect 95 24314 107 24348
rect 49 24280 107 24314
rect 49 24246 61 24280
rect 95 24246 107 24280
rect 49 24212 107 24246
rect 49 24178 61 24212
rect 95 24178 107 24212
rect 49 24144 107 24178
rect 49 24110 61 24144
rect 95 24110 107 24144
rect 49 24076 107 24110
rect 49 24042 61 24076
rect 95 24042 107 24076
rect 49 24008 107 24042
rect 49 23974 61 24008
rect 95 23974 107 24008
rect 49 23940 107 23974
rect 49 23906 61 23940
rect 95 23906 107 23940
rect 49 23872 107 23906
rect 49 23838 61 23872
rect 95 23838 107 23872
rect 49 23804 107 23838
rect 49 23770 61 23804
rect 95 23770 107 23804
rect 49 23736 107 23770
rect 49 23702 61 23736
rect 95 23702 107 23736
rect 49 23661 107 23702
rect 207 24620 265 24661
rect 207 24586 219 24620
rect 253 24586 265 24620
rect 207 24552 265 24586
rect 207 24518 219 24552
rect 253 24518 265 24552
rect 207 24484 265 24518
rect 207 24450 219 24484
rect 253 24450 265 24484
rect 207 24416 265 24450
rect 207 24382 219 24416
rect 253 24382 265 24416
rect 207 24348 265 24382
rect 207 24314 219 24348
rect 253 24314 265 24348
rect 207 24280 265 24314
rect 207 24246 219 24280
rect 253 24246 265 24280
rect 207 24212 265 24246
rect 207 24178 219 24212
rect 253 24178 265 24212
rect 207 24144 265 24178
rect 207 24110 219 24144
rect 253 24110 265 24144
rect 207 24076 265 24110
rect 207 24042 219 24076
rect 253 24042 265 24076
rect 207 24008 265 24042
rect 207 23974 219 24008
rect 253 23974 265 24008
rect 207 23940 265 23974
rect 207 23906 219 23940
rect 253 23906 265 23940
rect 207 23872 265 23906
rect 207 23838 219 23872
rect 253 23838 265 23872
rect 207 23804 265 23838
rect 207 23770 219 23804
rect 253 23770 265 23804
rect 207 23736 265 23770
rect 207 23702 219 23736
rect 253 23702 265 23736
rect 207 23661 265 23702
rect 365 24620 423 24661
rect 365 24586 377 24620
rect 411 24586 423 24620
rect 365 24552 423 24586
rect 365 24518 377 24552
rect 411 24518 423 24552
rect 365 24484 423 24518
rect 365 24450 377 24484
rect 411 24450 423 24484
rect 365 24416 423 24450
rect 365 24382 377 24416
rect 411 24382 423 24416
rect 365 24348 423 24382
rect 365 24314 377 24348
rect 411 24314 423 24348
rect 365 24280 423 24314
rect 365 24246 377 24280
rect 411 24246 423 24280
rect 365 24212 423 24246
rect 365 24178 377 24212
rect 411 24178 423 24212
rect 365 24144 423 24178
rect 365 24110 377 24144
rect 411 24110 423 24144
rect 365 24076 423 24110
rect 365 24042 377 24076
rect 411 24042 423 24076
rect 365 24008 423 24042
rect 365 23974 377 24008
rect 411 23974 423 24008
rect 365 23940 423 23974
rect 365 23906 377 23940
rect 411 23906 423 23940
rect 365 23872 423 23906
rect 365 23838 377 23872
rect 411 23838 423 23872
rect 365 23804 423 23838
rect 365 23770 377 23804
rect 411 23770 423 23804
rect 365 23736 423 23770
rect 365 23702 377 23736
rect 411 23702 423 23736
rect 365 23661 423 23702
rect 523 24620 581 24661
rect 523 24586 535 24620
rect 569 24586 581 24620
rect 523 24552 581 24586
rect 523 24518 535 24552
rect 569 24518 581 24552
rect 523 24484 581 24518
rect 523 24450 535 24484
rect 569 24450 581 24484
rect 523 24416 581 24450
rect 523 24382 535 24416
rect 569 24382 581 24416
rect 523 24348 581 24382
rect 523 24314 535 24348
rect 569 24314 581 24348
rect 523 24280 581 24314
rect 523 24246 535 24280
rect 569 24246 581 24280
rect 523 24212 581 24246
rect 523 24178 535 24212
rect 569 24178 581 24212
rect 523 24144 581 24178
rect 523 24110 535 24144
rect 569 24110 581 24144
rect 523 24076 581 24110
rect 523 24042 535 24076
rect 569 24042 581 24076
rect 523 24008 581 24042
rect 523 23974 535 24008
rect 569 23974 581 24008
rect 523 23940 581 23974
rect 523 23906 535 23940
rect 569 23906 581 23940
rect 523 23872 581 23906
rect 523 23838 535 23872
rect 569 23838 581 23872
rect 523 23804 581 23838
rect 523 23770 535 23804
rect 569 23770 581 23804
rect 523 23736 581 23770
rect 523 23702 535 23736
rect 569 23702 581 23736
rect 523 23661 581 23702
rect -1574 23099 -1516 23140
rect -1574 23065 -1562 23099
rect -1528 23065 -1516 23099
rect -1574 23031 -1516 23065
rect -1574 22997 -1562 23031
rect -1528 22997 -1516 23031
rect -1574 22963 -1516 22997
rect -1574 22929 -1562 22963
rect -1528 22929 -1516 22963
rect -1574 22895 -1516 22929
rect -1574 22861 -1562 22895
rect -1528 22861 -1516 22895
rect -1574 22827 -1516 22861
rect -1574 22793 -1562 22827
rect -1528 22793 -1516 22827
rect -1574 22759 -1516 22793
rect -1574 22725 -1562 22759
rect -1528 22725 -1516 22759
rect -1574 22691 -1516 22725
rect -1574 22657 -1562 22691
rect -1528 22657 -1516 22691
rect -1574 22623 -1516 22657
rect -1574 22589 -1562 22623
rect -1528 22589 -1516 22623
rect -1574 22555 -1516 22589
rect -1574 22521 -1562 22555
rect -1528 22521 -1516 22555
rect -1574 22487 -1516 22521
rect -1574 22453 -1562 22487
rect -1528 22453 -1516 22487
rect -1574 22419 -1516 22453
rect -1574 22385 -1562 22419
rect -1528 22385 -1516 22419
rect -1574 22351 -1516 22385
rect -1574 22317 -1562 22351
rect -1528 22317 -1516 22351
rect -1574 22283 -1516 22317
rect -1574 22249 -1562 22283
rect -1528 22249 -1516 22283
rect -1574 22215 -1516 22249
rect -1574 22181 -1562 22215
rect -1528 22181 -1516 22215
rect -1574 22140 -1516 22181
rect -1316 23099 -1258 23140
rect -1316 23065 -1304 23099
rect -1270 23065 -1258 23099
rect -1316 23031 -1258 23065
rect -1316 22997 -1304 23031
rect -1270 22997 -1258 23031
rect -1316 22963 -1258 22997
rect -1316 22929 -1304 22963
rect -1270 22929 -1258 22963
rect -1316 22895 -1258 22929
rect -1316 22861 -1304 22895
rect -1270 22861 -1258 22895
rect -1316 22827 -1258 22861
rect -1316 22793 -1304 22827
rect -1270 22793 -1258 22827
rect -1316 22759 -1258 22793
rect -1316 22725 -1304 22759
rect -1270 22725 -1258 22759
rect -1316 22691 -1258 22725
rect -1316 22657 -1304 22691
rect -1270 22657 -1258 22691
rect -1316 22623 -1258 22657
rect -1316 22589 -1304 22623
rect -1270 22589 -1258 22623
rect -1316 22555 -1258 22589
rect -1316 22521 -1304 22555
rect -1270 22521 -1258 22555
rect -1316 22487 -1258 22521
rect -1316 22453 -1304 22487
rect -1270 22453 -1258 22487
rect -1316 22419 -1258 22453
rect -1316 22385 -1304 22419
rect -1270 22385 -1258 22419
rect -1316 22351 -1258 22385
rect -1316 22317 -1304 22351
rect -1270 22317 -1258 22351
rect -1316 22283 -1258 22317
rect -1316 22249 -1304 22283
rect -1270 22249 -1258 22283
rect -1316 22215 -1258 22249
rect -1316 22181 -1304 22215
rect -1270 22181 -1258 22215
rect -1316 22140 -1258 22181
rect -1058 23099 -1000 23140
rect -1058 23065 -1046 23099
rect -1012 23065 -1000 23099
rect -1058 23031 -1000 23065
rect -1058 22997 -1046 23031
rect -1012 22997 -1000 23031
rect -1058 22963 -1000 22997
rect -1058 22929 -1046 22963
rect -1012 22929 -1000 22963
rect -1058 22895 -1000 22929
rect -1058 22861 -1046 22895
rect -1012 22861 -1000 22895
rect -1058 22827 -1000 22861
rect -1058 22793 -1046 22827
rect -1012 22793 -1000 22827
rect -1058 22759 -1000 22793
rect -1058 22725 -1046 22759
rect -1012 22725 -1000 22759
rect -1058 22691 -1000 22725
rect -1058 22657 -1046 22691
rect -1012 22657 -1000 22691
rect -1058 22623 -1000 22657
rect -1058 22589 -1046 22623
rect -1012 22589 -1000 22623
rect -1058 22555 -1000 22589
rect -1058 22521 -1046 22555
rect -1012 22521 -1000 22555
rect -1058 22487 -1000 22521
rect -1058 22453 -1046 22487
rect -1012 22453 -1000 22487
rect -1058 22419 -1000 22453
rect -1058 22385 -1046 22419
rect -1012 22385 -1000 22419
rect -1058 22351 -1000 22385
rect -1058 22317 -1046 22351
rect -1012 22317 -1000 22351
rect -1058 22283 -1000 22317
rect -1058 22249 -1046 22283
rect -1012 22249 -1000 22283
rect -1058 22215 -1000 22249
rect -1058 22181 -1046 22215
rect -1012 22181 -1000 22215
rect -1058 22140 -1000 22181
rect -800 23099 -742 23140
rect -800 23065 -788 23099
rect -754 23065 -742 23099
rect -800 23031 -742 23065
rect -800 22997 -788 23031
rect -754 22997 -742 23031
rect -800 22963 -742 22997
rect -800 22929 -788 22963
rect -754 22929 -742 22963
rect -800 22895 -742 22929
rect -800 22861 -788 22895
rect -754 22861 -742 22895
rect -800 22827 -742 22861
rect -800 22793 -788 22827
rect -754 22793 -742 22827
rect -800 22759 -742 22793
rect -800 22725 -788 22759
rect -754 22725 -742 22759
rect -800 22691 -742 22725
rect -800 22657 -788 22691
rect -754 22657 -742 22691
rect -800 22623 -742 22657
rect -800 22589 -788 22623
rect -754 22589 -742 22623
rect -800 22555 -742 22589
rect -800 22521 -788 22555
rect -754 22521 -742 22555
rect -800 22487 -742 22521
rect -800 22453 -788 22487
rect -754 22453 -742 22487
rect -800 22419 -742 22453
rect -800 22385 -788 22419
rect -754 22385 -742 22419
rect -800 22351 -742 22385
rect -800 22317 -788 22351
rect -754 22317 -742 22351
rect -800 22283 -742 22317
rect -800 22249 -788 22283
rect -754 22249 -742 22283
rect -800 22215 -742 22249
rect -800 22181 -788 22215
rect -754 22181 -742 22215
rect -800 22140 -742 22181
rect -542 23099 -484 23140
rect -542 23065 -530 23099
rect -496 23065 -484 23099
rect -542 23031 -484 23065
rect -542 22997 -530 23031
rect -496 22997 -484 23031
rect -542 22963 -484 22997
rect -542 22929 -530 22963
rect -496 22929 -484 22963
rect -542 22895 -484 22929
rect -542 22861 -530 22895
rect -496 22861 -484 22895
rect -542 22827 -484 22861
rect -542 22793 -530 22827
rect -496 22793 -484 22827
rect -542 22759 -484 22793
rect -542 22725 -530 22759
rect -496 22725 -484 22759
rect -542 22691 -484 22725
rect -542 22657 -530 22691
rect -496 22657 -484 22691
rect -542 22623 -484 22657
rect -542 22589 -530 22623
rect -496 22589 -484 22623
rect -542 22555 -484 22589
rect -542 22521 -530 22555
rect -496 22521 -484 22555
rect -542 22487 -484 22521
rect -542 22453 -530 22487
rect -496 22453 -484 22487
rect -542 22419 -484 22453
rect -542 22385 -530 22419
rect -496 22385 -484 22419
rect -542 22351 -484 22385
rect -542 22317 -530 22351
rect -496 22317 -484 22351
rect -542 22283 -484 22317
rect -542 22249 -530 22283
rect -496 22249 -484 22283
rect -542 22215 -484 22249
rect -542 22181 -530 22215
rect -496 22181 -484 22215
rect -542 22140 -484 22181
rect -284 23099 -226 23140
rect -284 23065 -272 23099
rect -238 23065 -226 23099
rect -284 23031 -226 23065
rect -284 22997 -272 23031
rect -238 22997 -226 23031
rect -284 22963 -226 22997
rect -284 22929 -272 22963
rect -238 22929 -226 22963
rect -284 22895 -226 22929
rect -284 22861 -272 22895
rect -238 22861 -226 22895
rect -284 22827 -226 22861
rect -284 22793 -272 22827
rect -238 22793 -226 22827
rect -284 22759 -226 22793
rect -284 22725 -272 22759
rect -238 22725 -226 22759
rect -284 22691 -226 22725
rect -284 22657 -272 22691
rect -238 22657 -226 22691
rect -284 22623 -226 22657
rect -284 22589 -272 22623
rect -238 22589 -226 22623
rect -284 22555 -226 22589
rect -284 22521 -272 22555
rect -238 22521 -226 22555
rect -284 22487 -226 22521
rect -284 22453 -272 22487
rect -238 22453 -226 22487
rect -284 22419 -226 22453
rect -284 22385 -272 22419
rect -238 22385 -226 22419
rect -284 22351 -226 22385
rect -284 22317 -272 22351
rect -238 22317 -226 22351
rect -284 22283 -226 22317
rect -284 22249 -272 22283
rect -238 22249 -226 22283
rect -284 22215 -226 22249
rect -284 22181 -272 22215
rect -238 22181 -226 22215
rect -284 22140 -226 22181
rect -26 23099 32 23140
rect -26 23065 -14 23099
rect 20 23065 32 23099
rect -26 23031 32 23065
rect -26 22997 -14 23031
rect 20 22997 32 23031
rect -26 22963 32 22997
rect -26 22929 -14 22963
rect 20 22929 32 22963
rect -26 22895 32 22929
rect -26 22861 -14 22895
rect 20 22861 32 22895
rect -26 22827 32 22861
rect -26 22793 -14 22827
rect 20 22793 32 22827
rect -26 22759 32 22793
rect -26 22725 -14 22759
rect 20 22725 32 22759
rect -26 22691 32 22725
rect -26 22657 -14 22691
rect 20 22657 32 22691
rect -26 22623 32 22657
rect -26 22589 -14 22623
rect 20 22589 32 22623
rect -26 22555 32 22589
rect -26 22521 -14 22555
rect 20 22521 32 22555
rect -26 22487 32 22521
rect -26 22453 -14 22487
rect 20 22453 32 22487
rect -26 22419 32 22453
rect -26 22385 -14 22419
rect 20 22385 32 22419
rect -26 22351 32 22385
rect -26 22317 -14 22351
rect 20 22317 32 22351
rect -26 22283 32 22317
rect -26 22249 -14 22283
rect 20 22249 32 22283
rect -26 22215 32 22249
rect -26 22181 -14 22215
rect 20 22181 32 22215
rect -26 22140 32 22181
rect 232 23099 290 23140
rect 232 23065 244 23099
rect 278 23065 290 23099
rect 232 23031 290 23065
rect 232 22997 244 23031
rect 278 22997 290 23031
rect 232 22963 290 22997
rect 232 22929 244 22963
rect 278 22929 290 22963
rect 232 22895 290 22929
rect 232 22861 244 22895
rect 278 22861 290 22895
rect 232 22827 290 22861
rect 232 22793 244 22827
rect 278 22793 290 22827
rect 232 22759 290 22793
rect 232 22725 244 22759
rect 278 22725 290 22759
rect 232 22691 290 22725
rect 232 22657 244 22691
rect 278 22657 290 22691
rect 232 22623 290 22657
rect 232 22589 244 22623
rect 278 22589 290 22623
rect 232 22555 290 22589
rect 232 22521 244 22555
rect 278 22521 290 22555
rect 232 22487 290 22521
rect 232 22453 244 22487
rect 278 22453 290 22487
rect 232 22419 290 22453
rect 232 22385 244 22419
rect 278 22385 290 22419
rect 232 22351 290 22385
rect 232 22317 244 22351
rect 278 22317 290 22351
rect 232 22283 290 22317
rect 232 22249 244 22283
rect 278 22249 290 22283
rect 232 22215 290 22249
rect 232 22181 244 22215
rect 278 22181 290 22215
rect 232 22140 290 22181
rect 490 23099 548 23140
rect 490 23065 502 23099
rect 536 23065 548 23099
rect 490 23031 548 23065
rect 490 22997 502 23031
rect 536 22997 548 23031
rect 490 22963 548 22997
rect 490 22929 502 22963
rect 536 22929 548 22963
rect 490 22895 548 22929
rect 490 22861 502 22895
rect 536 22861 548 22895
rect 490 22827 548 22861
rect 490 22793 502 22827
rect 536 22793 548 22827
rect 490 22759 548 22793
rect 490 22725 502 22759
rect 536 22725 548 22759
rect 490 22691 548 22725
rect 490 22657 502 22691
rect 536 22657 548 22691
rect 490 22623 548 22657
rect 490 22589 502 22623
rect 536 22589 548 22623
rect 490 22555 548 22589
rect 490 22521 502 22555
rect 536 22521 548 22555
rect 490 22487 548 22521
rect 490 22453 502 22487
rect 536 22453 548 22487
rect 490 22419 548 22453
rect 490 22385 502 22419
rect 536 22385 548 22419
rect 490 22351 548 22385
rect 490 22317 502 22351
rect 536 22317 548 22351
rect 490 22283 548 22317
rect 490 22249 502 22283
rect 536 22249 548 22283
rect 490 22215 548 22249
rect 490 22181 502 22215
rect 536 22181 548 22215
rect 490 22140 548 22181
rect 748 23099 806 23140
rect 748 23065 760 23099
rect 794 23065 806 23099
rect 748 23031 806 23065
rect 748 22997 760 23031
rect 794 22997 806 23031
rect 748 22963 806 22997
rect 748 22929 760 22963
rect 794 22929 806 22963
rect 748 22895 806 22929
rect 748 22861 760 22895
rect 794 22861 806 22895
rect 748 22827 806 22861
rect 748 22793 760 22827
rect 794 22793 806 22827
rect 748 22759 806 22793
rect 748 22725 760 22759
rect 794 22725 806 22759
rect 748 22691 806 22725
rect 748 22657 760 22691
rect 794 22657 806 22691
rect 748 22623 806 22657
rect 748 22589 760 22623
rect 794 22589 806 22623
rect 748 22555 806 22589
rect 748 22521 760 22555
rect 794 22521 806 22555
rect 748 22487 806 22521
rect 748 22453 760 22487
rect 794 22453 806 22487
rect 748 22419 806 22453
rect 748 22385 760 22419
rect 794 22385 806 22419
rect 748 22351 806 22385
rect 748 22317 760 22351
rect 794 22317 806 22351
rect 748 22283 806 22317
rect 748 22249 760 22283
rect 794 22249 806 22283
rect 748 22215 806 22249
rect 748 22181 760 22215
rect 794 22181 806 22215
rect 748 22140 806 22181
rect 1006 23099 1064 23140
rect 1006 23065 1018 23099
rect 1052 23065 1064 23099
rect 1006 23031 1064 23065
rect 1006 22997 1018 23031
rect 1052 22997 1064 23031
rect 1006 22963 1064 22997
rect 1006 22929 1018 22963
rect 1052 22929 1064 22963
rect 1006 22895 1064 22929
rect 1006 22861 1018 22895
rect 1052 22861 1064 22895
rect 1006 22827 1064 22861
rect 1006 22793 1018 22827
rect 1052 22793 1064 22827
rect 1006 22759 1064 22793
rect 1006 22725 1018 22759
rect 1052 22725 1064 22759
rect 1006 22691 1064 22725
rect 1006 22657 1018 22691
rect 1052 22657 1064 22691
rect 1006 22623 1064 22657
rect 1006 22589 1018 22623
rect 1052 22589 1064 22623
rect 1006 22555 1064 22589
rect 1006 22521 1018 22555
rect 1052 22521 1064 22555
rect 1006 22487 1064 22521
rect 1006 22453 1018 22487
rect 1052 22453 1064 22487
rect 1006 22419 1064 22453
rect 1006 22385 1018 22419
rect 1052 22385 1064 22419
rect 1006 22351 1064 22385
rect 1006 22317 1018 22351
rect 1052 22317 1064 22351
rect 1006 22283 1064 22317
rect 1006 22249 1018 22283
rect 1052 22249 1064 22283
rect 1006 22215 1064 22249
rect 1006 22181 1018 22215
rect 1052 22181 1064 22215
rect 1006 22140 1064 22181
rect 1264 23099 1322 23140
rect 1264 23065 1276 23099
rect 1310 23065 1322 23099
rect 1264 23031 1322 23065
rect 1264 22997 1276 23031
rect 1310 22997 1322 23031
rect 1264 22963 1322 22997
rect 1264 22929 1276 22963
rect 1310 22929 1322 22963
rect 1264 22895 1322 22929
rect 1264 22861 1276 22895
rect 1310 22861 1322 22895
rect 1264 22827 1322 22861
rect 1264 22793 1276 22827
rect 1310 22793 1322 22827
rect 1264 22759 1322 22793
rect 1264 22725 1276 22759
rect 1310 22725 1322 22759
rect 1264 22691 1322 22725
rect 1264 22657 1276 22691
rect 1310 22657 1322 22691
rect 1264 22623 1322 22657
rect 1264 22589 1276 22623
rect 1310 22589 1322 22623
rect 1264 22555 1322 22589
rect 1264 22521 1276 22555
rect 1310 22521 1322 22555
rect 1264 22487 1322 22521
rect 1264 22453 1276 22487
rect 1310 22453 1322 22487
rect 1264 22419 1322 22453
rect 1264 22385 1276 22419
rect 1310 22385 1322 22419
rect 1264 22351 1322 22385
rect 1264 22317 1276 22351
rect 1310 22317 1322 22351
rect 1264 22283 1322 22317
rect 1264 22249 1276 22283
rect 1310 22249 1322 22283
rect 1264 22215 1322 22249
rect 1264 22181 1276 22215
rect 1310 22181 1322 22215
rect 1264 22140 1322 22181
rect 1522 23099 1580 23140
rect 1522 23065 1534 23099
rect 1568 23065 1580 23099
rect 1522 23031 1580 23065
rect 1522 22997 1534 23031
rect 1568 22997 1580 23031
rect 1522 22963 1580 22997
rect 1522 22929 1534 22963
rect 1568 22929 1580 22963
rect 1522 22895 1580 22929
rect 1522 22861 1534 22895
rect 1568 22861 1580 22895
rect 1522 22827 1580 22861
rect 1522 22793 1534 22827
rect 1568 22793 1580 22827
rect 1522 22759 1580 22793
rect 1522 22725 1534 22759
rect 1568 22725 1580 22759
rect 1522 22691 1580 22725
rect 1522 22657 1534 22691
rect 1568 22657 1580 22691
rect 1522 22623 1580 22657
rect 1522 22589 1534 22623
rect 1568 22589 1580 22623
rect 1522 22555 1580 22589
rect 1522 22521 1534 22555
rect 1568 22521 1580 22555
rect 1522 22487 1580 22521
rect 1522 22453 1534 22487
rect 1568 22453 1580 22487
rect 1522 22419 1580 22453
rect 1522 22385 1534 22419
rect 1568 22385 1580 22419
rect 1522 22351 1580 22385
rect 1522 22317 1534 22351
rect 1568 22317 1580 22351
rect 1522 22283 1580 22317
rect 1522 22249 1534 22283
rect 1568 22249 1580 22283
rect 1522 22215 1580 22249
rect 1522 22181 1534 22215
rect 1568 22181 1580 22215
rect 1522 22140 1580 22181
rect -1834 21579 -1776 21620
rect -1834 21545 -1822 21579
rect -1788 21545 -1776 21579
rect -1834 21511 -1776 21545
rect -1834 21477 -1822 21511
rect -1788 21477 -1776 21511
rect -1834 21443 -1776 21477
rect -1834 21409 -1822 21443
rect -1788 21409 -1776 21443
rect -1834 21375 -1776 21409
rect -1834 21341 -1822 21375
rect -1788 21341 -1776 21375
rect -1834 21307 -1776 21341
rect -1834 21273 -1822 21307
rect -1788 21273 -1776 21307
rect -1834 21239 -1776 21273
rect -1834 21205 -1822 21239
rect -1788 21205 -1776 21239
rect -1834 21171 -1776 21205
rect -1834 21137 -1822 21171
rect -1788 21137 -1776 21171
rect -1834 21103 -1776 21137
rect -1834 21069 -1822 21103
rect -1788 21069 -1776 21103
rect -1834 21035 -1776 21069
rect -1834 21001 -1822 21035
rect -1788 21001 -1776 21035
rect -1834 20967 -1776 21001
rect -1834 20933 -1822 20967
rect -1788 20933 -1776 20967
rect -1834 20899 -1776 20933
rect -1834 20865 -1822 20899
rect -1788 20865 -1776 20899
rect -1834 20831 -1776 20865
rect -1834 20797 -1822 20831
rect -1788 20797 -1776 20831
rect -1834 20763 -1776 20797
rect -1834 20729 -1822 20763
rect -1788 20729 -1776 20763
rect -1834 20695 -1776 20729
rect -1834 20661 -1822 20695
rect -1788 20661 -1776 20695
rect -1834 20620 -1776 20661
rect -1576 21579 -1518 21620
rect -1576 21545 -1564 21579
rect -1530 21545 -1518 21579
rect -1576 21511 -1518 21545
rect -1576 21477 -1564 21511
rect -1530 21477 -1518 21511
rect -1576 21443 -1518 21477
rect -1576 21409 -1564 21443
rect -1530 21409 -1518 21443
rect -1576 21375 -1518 21409
rect -1576 21341 -1564 21375
rect -1530 21341 -1518 21375
rect -1576 21307 -1518 21341
rect -1576 21273 -1564 21307
rect -1530 21273 -1518 21307
rect -1576 21239 -1518 21273
rect -1576 21205 -1564 21239
rect -1530 21205 -1518 21239
rect -1576 21171 -1518 21205
rect -1576 21137 -1564 21171
rect -1530 21137 -1518 21171
rect -1576 21103 -1518 21137
rect -1576 21069 -1564 21103
rect -1530 21069 -1518 21103
rect -1576 21035 -1518 21069
rect -1576 21001 -1564 21035
rect -1530 21001 -1518 21035
rect -1576 20967 -1518 21001
rect -1576 20933 -1564 20967
rect -1530 20933 -1518 20967
rect -1576 20899 -1518 20933
rect -1576 20865 -1564 20899
rect -1530 20865 -1518 20899
rect -1576 20831 -1518 20865
rect -1576 20797 -1564 20831
rect -1530 20797 -1518 20831
rect -1576 20763 -1518 20797
rect -1576 20729 -1564 20763
rect -1530 20729 -1518 20763
rect -1576 20695 -1518 20729
rect -1576 20661 -1564 20695
rect -1530 20661 -1518 20695
rect -1576 20620 -1518 20661
rect -1318 21579 -1260 21620
rect -1318 21545 -1306 21579
rect -1272 21545 -1260 21579
rect -1318 21511 -1260 21545
rect -1318 21477 -1306 21511
rect -1272 21477 -1260 21511
rect -1318 21443 -1260 21477
rect -1318 21409 -1306 21443
rect -1272 21409 -1260 21443
rect -1318 21375 -1260 21409
rect -1318 21341 -1306 21375
rect -1272 21341 -1260 21375
rect -1318 21307 -1260 21341
rect -1318 21273 -1306 21307
rect -1272 21273 -1260 21307
rect -1318 21239 -1260 21273
rect -1318 21205 -1306 21239
rect -1272 21205 -1260 21239
rect -1318 21171 -1260 21205
rect -1318 21137 -1306 21171
rect -1272 21137 -1260 21171
rect -1318 21103 -1260 21137
rect -1318 21069 -1306 21103
rect -1272 21069 -1260 21103
rect -1318 21035 -1260 21069
rect -1318 21001 -1306 21035
rect -1272 21001 -1260 21035
rect -1318 20967 -1260 21001
rect -1318 20933 -1306 20967
rect -1272 20933 -1260 20967
rect -1318 20899 -1260 20933
rect -1318 20865 -1306 20899
rect -1272 20865 -1260 20899
rect -1318 20831 -1260 20865
rect -1318 20797 -1306 20831
rect -1272 20797 -1260 20831
rect -1318 20763 -1260 20797
rect -1318 20729 -1306 20763
rect -1272 20729 -1260 20763
rect -1318 20695 -1260 20729
rect -1318 20661 -1306 20695
rect -1272 20661 -1260 20695
rect -1318 20620 -1260 20661
rect -1060 21579 -1002 21620
rect -1060 21545 -1048 21579
rect -1014 21545 -1002 21579
rect -1060 21511 -1002 21545
rect -1060 21477 -1048 21511
rect -1014 21477 -1002 21511
rect -1060 21443 -1002 21477
rect -1060 21409 -1048 21443
rect -1014 21409 -1002 21443
rect -1060 21375 -1002 21409
rect -1060 21341 -1048 21375
rect -1014 21341 -1002 21375
rect -1060 21307 -1002 21341
rect -1060 21273 -1048 21307
rect -1014 21273 -1002 21307
rect -1060 21239 -1002 21273
rect -1060 21205 -1048 21239
rect -1014 21205 -1002 21239
rect -1060 21171 -1002 21205
rect -1060 21137 -1048 21171
rect -1014 21137 -1002 21171
rect -1060 21103 -1002 21137
rect -1060 21069 -1048 21103
rect -1014 21069 -1002 21103
rect -1060 21035 -1002 21069
rect -1060 21001 -1048 21035
rect -1014 21001 -1002 21035
rect -1060 20967 -1002 21001
rect -1060 20933 -1048 20967
rect -1014 20933 -1002 20967
rect -1060 20899 -1002 20933
rect -1060 20865 -1048 20899
rect -1014 20865 -1002 20899
rect -1060 20831 -1002 20865
rect -1060 20797 -1048 20831
rect -1014 20797 -1002 20831
rect -1060 20763 -1002 20797
rect -1060 20729 -1048 20763
rect -1014 20729 -1002 20763
rect -1060 20695 -1002 20729
rect -1060 20661 -1048 20695
rect -1014 20661 -1002 20695
rect -1060 20620 -1002 20661
rect -802 21579 -744 21620
rect -802 21545 -790 21579
rect -756 21545 -744 21579
rect -802 21511 -744 21545
rect -802 21477 -790 21511
rect -756 21477 -744 21511
rect -802 21443 -744 21477
rect -802 21409 -790 21443
rect -756 21409 -744 21443
rect -802 21375 -744 21409
rect -802 21341 -790 21375
rect -756 21341 -744 21375
rect -802 21307 -744 21341
rect -802 21273 -790 21307
rect -756 21273 -744 21307
rect -802 21239 -744 21273
rect -802 21205 -790 21239
rect -756 21205 -744 21239
rect -802 21171 -744 21205
rect -802 21137 -790 21171
rect -756 21137 -744 21171
rect -802 21103 -744 21137
rect -802 21069 -790 21103
rect -756 21069 -744 21103
rect -802 21035 -744 21069
rect -802 21001 -790 21035
rect -756 21001 -744 21035
rect -802 20967 -744 21001
rect -802 20933 -790 20967
rect -756 20933 -744 20967
rect -802 20899 -744 20933
rect -802 20865 -790 20899
rect -756 20865 -744 20899
rect -802 20831 -744 20865
rect -802 20797 -790 20831
rect -756 20797 -744 20831
rect -802 20763 -744 20797
rect -802 20729 -790 20763
rect -756 20729 -744 20763
rect -802 20695 -744 20729
rect -802 20661 -790 20695
rect -756 20661 -744 20695
rect -802 20620 -744 20661
rect -544 21579 -486 21620
rect -544 21545 -532 21579
rect -498 21545 -486 21579
rect -544 21511 -486 21545
rect -544 21477 -532 21511
rect -498 21477 -486 21511
rect -544 21443 -486 21477
rect -544 21409 -532 21443
rect -498 21409 -486 21443
rect -544 21375 -486 21409
rect -544 21341 -532 21375
rect -498 21341 -486 21375
rect -544 21307 -486 21341
rect -544 21273 -532 21307
rect -498 21273 -486 21307
rect -544 21239 -486 21273
rect -544 21205 -532 21239
rect -498 21205 -486 21239
rect -544 21171 -486 21205
rect -544 21137 -532 21171
rect -498 21137 -486 21171
rect -544 21103 -486 21137
rect -544 21069 -532 21103
rect -498 21069 -486 21103
rect -544 21035 -486 21069
rect -544 21001 -532 21035
rect -498 21001 -486 21035
rect -544 20967 -486 21001
rect -544 20933 -532 20967
rect -498 20933 -486 20967
rect -544 20899 -486 20933
rect -544 20865 -532 20899
rect -498 20865 -486 20899
rect -544 20831 -486 20865
rect -544 20797 -532 20831
rect -498 20797 -486 20831
rect -544 20763 -486 20797
rect -544 20729 -532 20763
rect -498 20729 -486 20763
rect -544 20695 -486 20729
rect -544 20661 -532 20695
rect -498 20661 -486 20695
rect -544 20620 -486 20661
rect -286 21579 -228 21620
rect -286 21545 -274 21579
rect -240 21545 -228 21579
rect -286 21511 -228 21545
rect -286 21477 -274 21511
rect -240 21477 -228 21511
rect -286 21443 -228 21477
rect -286 21409 -274 21443
rect -240 21409 -228 21443
rect -286 21375 -228 21409
rect -286 21341 -274 21375
rect -240 21341 -228 21375
rect -286 21307 -228 21341
rect -286 21273 -274 21307
rect -240 21273 -228 21307
rect -286 21239 -228 21273
rect -286 21205 -274 21239
rect -240 21205 -228 21239
rect -286 21171 -228 21205
rect -286 21137 -274 21171
rect -240 21137 -228 21171
rect -286 21103 -228 21137
rect -286 21069 -274 21103
rect -240 21069 -228 21103
rect -286 21035 -228 21069
rect -286 21001 -274 21035
rect -240 21001 -228 21035
rect -286 20967 -228 21001
rect -286 20933 -274 20967
rect -240 20933 -228 20967
rect -286 20899 -228 20933
rect -286 20865 -274 20899
rect -240 20865 -228 20899
rect -286 20831 -228 20865
rect -286 20797 -274 20831
rect -240 20797 -228 20831
rect -286 20763 -228 20797
rect -286 20729 -274 20763
rect -240 20729 -228 20763
rect -286 20695 -228 20729
rect -286 20661 -274 20695
rect -240 20661 -228 20695
rect -286 20620 -228 20661
rect -28 21579 30 21620
rect -28 21545 -16 21579
rect 18 21545 30 21579
rect -28 21511 30 21545
rect -28 21477 -16 21511
rect 18 21477 30 21511
rect -28 21443 30 21477
rect -28 21409 -16 21443
rect 18 21409 30 21443
rect -28 21375 30 21409
rect -28 21341 -16 21375
rect 18 21341 30 21375
rect -28 21307 30 21341
rect -28 21273 -16 21307
rect 18 21273 30 21307
rect -28 21239 30 21273
rect -28 21205 -16 21239
rect 18 21205 30 21239
rect -28 21171 30 21205
rect -28 21137 -16 21171
rect 18 21137 30 21171
rect -28 21103 30 21137
rect -28 21069 -16 21103
rect 18 21069 30 21103
rect -28 21035 30 21069
rect -28 21001 -16 21035
rect 18 21001 30 21035
rect -28 20967 30 21001
rect -28 20933 -16 20967
rect 18 20933 30 20967
rect -28 20899 30 20933
rect -28 20865 -16 20899
rect 18 20865 30 20899
rect -28 20831 30 20865
rect -28 20797 -16 20831
rect 18 20797 30 20831
rect -28 20763 30 20797
rect -28 20729 -16 20763
rect 18 20729 30 20763
rect -28 20695 30 20729
rect -28 20661 -16 20695
rect 18 20661 30 20695
rect -28 20620 30 20661
rect 230 21579 288 21620
rect 230 21545 242 21579
rect 276 21545 288 21579
rect 230 21511 288 21545
rect 230 21477 242 21511
rect 276 21477 288 21511
rect 230 21443 288 21477
rect 230 21409 242 21443
rect 276 21409 288 21443
rect 230 21375 288 21409
rect 230 21341 242 21375
rect 276 21341 288 21375
rect 230 21307 288 21341
rect 230 21273 242 21307
rect 276 21273 288 21307
rect 230 21239 288 21273
rect 230 21205 242 21239
rect 276 21205 288 21239
rect 230 21171 288 21205
rect 230 21137 242 21171
rect 276 21137 288 21171
rect 230 21103 288 21137
rect 230 21069 242 21103
rect 276 21069 288 21103
rect 230 21035 288 21069
rect 230 21001 242 21035
rect 276 21001 288 21035
rect 230 20967 288 21001
rect 230 20933 242 20967
rect 276 20933 288 20967
rect 230 20899 288 20933
rect 230 20865 242 20899
rect 276 20865 288 20899
rect 230 20831 288 20865
rect 230 20797 242 20831
rect 276 20797 288 20831
rect 230 20763 288 20797
rect 230 20729 242 20763
rect 276 20729 288 20763
rect 230 20695 288 20729
rect 230 20661 242 20695
rect 276 20661 288 20695
rect 230 20620 288 20661
rect 488 21579 546 21620
rect 488 21545 500 21579
rect 534 21545 546 21579
rect 488 21511 546 21545
rect 488 21477 500 21511
rect 534 21477 546 21511
rect 488 21443 546 21477
rect 488 21409 500 21443
rect 534 21409 546 21443
rect 488 21375 546 21409
rect 488 21341 500 21375
rect 534 21341 546 21375
rect 488 21307 546 21341
rect 488 21273 500 21307
rect 534 21273 546 21307
rect 488 21239 546 21273
rect 488 21205 500 21239
rect 534 21205 546 21239
rect 488 21171 546 21205
rect 488 21137 500 21171
rect 534 21137 546 21171
rect 488 21103 546 21137
rect 488 21069 500 21103
rect 534 21069 546 21103
rect 488 21035 546 21069
rect 488 21001 500 21035
rect 534 21001 546 21035
rect 488 20967 546 21001
rect 488 20933 500 20967
rect 534 20933 546 20967
rect 488 20899 546 20933
rect 488 20865 500 20899
rect 534 20865 546 20899
rect 488 20831 546 20865
rect 488 20797 500 20831
rect 534 20797 546 20831
rect 488 20763 546 20797
rect 488 20729 500 20763
rect 534 20729 546 20763
rect 488 20695 546 20729
rect 488 20661 500 20695
rect 534 20661 546 20695
rect 488 20620 546 20661
rect 746 21579 804 21620
rect 746 21545 758 21579
rect 792 21545 804 21579
rect 746 21511 804 21545
rect 746 21477 758 21511
rect 792 21477 804 21511
rect 746 21443 804 21477
rect 746 21409 758 21443
rect 792 21409 804 21443
rect 746 21375 804 21409
rect 746 21341 758 21375
rect 792 21341 804 21375
rect 746 21307 804 21341
rect 746 21273 758 21307
rect 792 21273 804 21307
rect 746 21239 804 21273
rect 746 21205 758 21239
rect 792 21205 804 21239
rect 746 21171 804 21205
rect 746 21137 758 21171
rect 792 21137 804 21171
rect 746 21103 804 21137
rect 746 21069 758 21103
rect 792 21069 804 21103
rect 746 21035 804 21069
rect 746 21001 758 21035
rect 792 21001 804 21035
rect 746 20967 804 21001
rect 746 20933 758 20967
rect 792 20933 804 20967
rect 746 20899 804 20933
rect 746 20865 758 20899
rect 792 20865 804 20899
rect 746 20831 804 20865
rect 746 20797 758 20831
rect 792 20797 804 20831
rect 746 20763 804 20797
rect 746 20729 758 20763
rect 792 20729 804 20763
rect 746 20695 804 20729
rect 746 20661 758 20695
rect 792 20661 804 20695
rect 746 20620 804 20661
rect 1004 21579 1062 21620
rect 1004 21545 1016 21579
rect 1050 21545 1062 21579
rect 1004 21511 1062 21545
rect 1004 21477 1016 21511
rect 1050 21477 1062 21511
rect 1004 21443 1062 21477
rect 1004 21409 1016 21443
rect 1050 21409 1062 21443
rect 1004 21375 1062 21409
rect 1004 21341 1016 21375
rect 1050 21341 1062 21375
rect 1004 21307 1062 21341
rect 1004 21273 1016 21307
rect 1050 21273 1062 21307
rect 1004 21239 1062 21273
rect 1004 21205 1016 21239
rect 1050 21205 1062 21239
rect 1004 21171 1062 21205
rect 1004 21137 1016 21171
rect 1050 21137 1062 21171
rect 1004 21103 1062 21137
rect 1004 21069 1016 21103
rect 1050 21069 1062 21103
rect 1004 21035 1062 21069
rect 1004 21001 1016 21035
rect 1050 21001 1062 21035
rect 1004 20967 1062 21001
rect 1004 20933 1016 20967
rect 1050 20933 1062 20967
rect 1004 20899 1062 20933
rect 1004 20865 1016 20899
rect 1050 20865 1062 20899
rect 1004 20831 1062 20865
rect 1004 20797 1016 20831
rect 1050 20797 1062 20831
rect 1004 20763 1062 20797
rect 1004 20729 1016 20763
rect 1050 20729 1062 20763
rect 1004 20695 1062 20729
rect 1004 20661 1016 20695
rect 1050 20661 1062 20695
rect 1004 20620 1062 20661
rect 1262 21579 1320 21620
rect 1262 21545 1274 21579
rect 1308 21545 1320 21579
rect 1262 21511 1320 21545
rect 1262 21477 1274 21511
rect 1308 21477 1320 21511
rect 1262 21443 1320 21477
rect 1262 21409 1274 21443
rect 1308 21409 1320 21443
rect 1262 21375 1320 21409
rect 1262 21341 1274 21375
rect 1308 21341 1320 21375
rect 1262 21307 1320 21341
rect 1262 21273 1274 21307
rect 1308 21273 1320 21307
rect 1262 21239 1320 21273
rect 1262 21205 1274 21239
rect 1308 21205 1320 21239
rect 1262 21171 1320 21205
rect 1262 21137 1274 21171
rect 1308 21137 1320 21171
rect 1262 21103 1320 21137
rect 1262 21069 1274 21103
rect 1308 21069 1320 21103
rect 1262 21035 1320 21069
rect 1262 21001 1274 21035
rect 1308 21001 1320 21035
rect 1262 20967 1320 21001
rect 1262 20933 1274 20967
rect 1308 20933 1320 20967
rect 1262 20899 1320 20933
rect 1262 20865 1274 20899
rect 1308 20865 1320 20899
rect 1262 20831 1320 20865
rect 1262 20797 1274 20831
rect 1308 20797 1320 20831
rect 1262 20763 1320 20797
rect 1262 20729 1274 20763
rect 1308 20729 1320 20763
rect 1262 20695 1320 20729
rect 1262 20661 1274 20695
rect 1308 20661 1320 20695
rect 1262 20620 1320 20661
rect 1520 21579 1578 21620
rect 1520 21545 1532 21579
rect 1566 21545 1578 21579
rect 1520 21511 1578 21545
rect 1520 21477 1532 21511
rect 1566 21477 1578 21511
rect 1520 21443 1578 21477
rect 1520 21409 1532 21443
rect 1566 21409 1578 21443
rect 1520 21375 1578 21409
rect 1520 21341 1532 21375
rect 1566 21341 1578 21375
rect 1520 21307 1578 21341
rect 1520 21273 1532 21307
rect 1566 21273 1578 21307
rect 1520 21239 1578 21273
rect 1520 21205 1532 21239
rect 1566 21205 1578 21239
rect 1520 21171 1578 21205
rect 1520 21137 1532 21171
rect 1566 21137 1578 21171
rect 1520 21103 1578 21137
rect 1520 21069 1532 21103
rect 1566 21069 1578 21103
rect 1520 21035 1578 21069
rect 1520 21001 1532 21035
rect 1566 21001 1578 21035
rect 1520 20967 1578 21001
rect 1520 20933 1532 20967
rect 1566 20933 1578 20967
rect 1520 20899 1578 20933
rect 1520 20865 1532 20899
rect 1566 20865 1578 20899
rect 1520 20831 1578 20865
rect 1520 20797 1532 20831
rect 1566 20797 1578 20831
rect 1520 20763 1578 20797
rect 1520 20729 1532 20763
rect 1566 20729 1578 20763
rect 1520 20695 1578 20729
rect 1520 20661 1532 20695
rect 1566 20661 1578 20695
rect 1520 20620 1578 20661
rect 1778 21579 1836 21620
rect 1778 21545 1790 21579
rect 1824 21545 1836 21579
rect 1778 21511 1836 21545
rect 1778 21477 1790 21511
rect 1824 21477 1836 21511
rect 1778 21443 1836 21477
rect 1778 21409 1790 21443
rect 1824 21409 1836 21443
rect 1778 21375 1836 21409
rect 1778 21341 1790 21375
rect 1824 21341 1836 21375
rect 1778 21307 1836 21341
rect 1778 21273 1790 21307
rect 1824 21273 1836 21307
rect 1778 21239 1836 21273
rect 1778 21205 1790 21239
rect 1824 21205 1836 21239
rect 1778 21171 1836 21205
rect 1778 21137 1790 21171
rect 1824 21137 1836 21171
rect 1778 21103 1836 21137
rect 1778 21069 1790 21103
rect 1824 21069 1836 21103
rect 1778 21035 1836 21069
rect 1778 21001 1790 21035
rect 1824 21001 1836 21035
rect 1778 20967 1836 21001
rect 1778 20933 1790 20967
rect 1824 20933 1836 20967
rect 1778 20899 1836 20933
rect 1778 20865 1790 20899
rect 1824 20865 1836 20899
rect 1778 20831 1836 20865
rect 1778 20797 1790 20831
rect 1824 20797 1836 20831
rect 1778 20763 1836 20797
rect 1778 20729 1790 20763
rect 1824 20729 1836 20763
rect 1778 20695 1836 20729
rect 1778 20661 1790 20695
rect 1824 20661 1836 20695
rect 1778 20620 1836 20661
rect -830 18052 -580 18064
rect -830 18018 -818 18052
rect -592 18018 -580 18052
rect -830 18006 -580 18018
rect -362 18052 -112 18064
rect -362 18018 -350 18052
rect -124 18018 -112 18052
rect -362 18006 -112 18018
rect 106 18052 356 18064
rect 106 18018 118 18052
rect 344 18018 356 18052
rect 106 18006 356 18018
rect 574 18052 824 18064
rect 574 18018 586 18052
rect 812 18018 824 18052
rect 574 18006 824 18018
rect -830 17794 -580 17806
rect -830 17760 -818 17794
rect -592 17760 -580 17794
rect -830 17748 -580 17760
rect -362 17794 -112 17806
rect -362 17760 -350 17794
rect -124 17760 -112 17794
rect -362 17748 -112 17760
rect 106 17794 356 17806
rect 106 17760 118 17794
rect 344 17760 356 17794
rect 106 17748 356 17760
rect 574 17794 824 17806
rect 574 17760 586 17794
rect 812 17760 824 17794
rect 574 17748 824 17760
rect -610 17427 -110 17439
rect -610 17393 -598 17427
rect -122 17393 -110 17427
rect -610 17381 -110 17393
rect 108 17427 608 17439
rect 108 17393 120 17427
rect 596 17393 608 17427
rect 108 17381 608 17393
rect -610 17269 -110 17281
rect -610 17235 -598 17269
rect -122 17235 -110 17269
rect -610 17223 -110 17235
rect 108 17269 608 17281
rect 108 17235 120 17269
rect 596 17235 608 17269
rect 108 17223 608 17235
rect -3545 16902 -2545 16914
rect -3545 16868 -3533 16902
rect -2557 16868 -2545 16902
rect -3545 16856 -2545 16868
rect -2327 16902 -1327 16914
rect -2327 16868 -2315 16902
rect -1339 16868 -1327 16902
rect -2327 16856 -1327 16868
rect -1109 16902 -109 16914
rect -1109 16868 -1097 16902
rect -121 16868 -109 16902
rect -1109 16856 -109 16868
rect 109 16902 1109 16914
rect 109 16868 121 16902
rect 1097 16868 1109 16902
rect 109 16856 1109 16868
rect 1327 16902 2327 16914
rect 1327 16868 1339 16902
rect 2315 16868 2327 16902
rect 1327 16856 2327 16868
rect 2545 16902 3545 16914
rect 2545 16868 2557 16902
rect 3533 16868 3545 16902
rect 2545 16856 3545 16868
rect -3545 16644 -2545 16656
rect -3545 16610 -3533 16644
rect -2557 16610 -2545 16644
rect -3545 16598 -2545 16610
rect -2327 16644 -1327 16656
rect -2327 16610 -2315 16644
rect -1339 16610 -1327 16644
rect -2327 16598 -1327 16610
rect -1109 16644 -109 16656
rect -1109 16610 -1097 16644
rect -121 16610 -109 16644
rect -1109 16598 -109 16610
rect 109 16644 1109 16656
rect 109 16610 121 16644
rect 1097 16610 1109 16644
rect 109 16598 1109 16610
rect 1327 16644 2327 16656
rect 1327 16610 1339 16644
rect 2315 16610 2327 16644
rect 1327 16598 2327 16610
rect 2545 16644 3545 16656
rect 2545 16610 2557 16644
rect 3533 16610 3545 16644
rect 2545 16598 3545 16610
<< pdiff >>
rect -3184 30918 -3126 30959
rect -3184 30884 -3172 30918
rect -3138 30884 -3126 30918
rect -3184 30850 -3126 30884
rect -3184 30816 -3172 30850
rect -3138 30816 -3126 30850
rect -3184 30782 -3126 30816
rect -3184 30748 -3172 30782
rect -3138 30748 -3126 30782
rect -3184 30714 -3126 30748
rect -3184 30680 -3172 30714
rect -3138 30680 -3126 30714
rect -3184 30646 -3126 30680
rect -3184 30612 -3172 30646
rect -3138 30612 -3126 30646
rect -3184 30578 -3126 30612
rect -3184 30544 -3172 30578
rect -3138 30544 -3126 30578
rect -3184 30510 -3126 30544
rect -3184 30476 -3172 30510
rect -3138 30476 -3126 30510
rect -3184 30442 -3126 30476
rect -3184 30408 -3172 30442
rect -3138 30408 -3126 30442
rect -3184 30374 -3126 30408
rect -3184 30340 -3172 30374
rect -3138 30340 -3126 30374
rect -3184 30306 -3126 30340
rect -3184 30272 -3172 30306
rect -3138 30272 -3126 30306
rect -3184 30238 -3126 30272
rect -3184 30204 -3172 30238
rect -3138 30204 -3126 30238
rect -3184 30170 -3126 30204
rect -3184 30136 -3172 30170
rect -3138 30136 -3126 30170
rect -3184 30102 -3126 30136
rect -3184 30068 -3172 30102
rect -3138 30068 -3126 30102
rect -3184 30034 -3126 30068
rect -3184 30000 -3172 30034
rect -3138 30000 -3126 30034
rect -3184 29959 -3126 30000
rect -3026 30918 -2968 30959
rect -3026 30884 -3014 30918
rect -2980 30884 -2968 30918
rect -3026 30850 -2968 30884
rect -3026 30816 -3014 30850
rect -2980 30816 -2968 30850
rect -3026 30782 -2968 30816
rect -3026 30748 -3014 30782
rect -2980 30748 -2968 30782
rect -3026 30714 -2968 30748
rect -3026 30680 -3014 30714
rect -2980 30680 -2968 30714
rect -3026 30646 -2968 30680
rect -3026 30612 -3014 30646
rect -2980 30612 -2968 30646
rect -3026 30578 -2968 30612
rect -3026 30544 -3014 30578
rect -2980 30544 -2968 30578
rect -3026 30510 -2968 30544
rect -3026 30476 -3014 30510
rect -2980 30476 -2968 30510
rect -3026 30442 -2968 30476
rect -3026 30408 -3014 30442
rect -2980 30408 -2968 30442
rect -3026 30374 -2968 30408
rect -3026 30340 -3014 30374
rect -2980 30340 -2968 30374
rect -3026 30306 -2968 30340
rect -3026 30272 -3014 30306
rect -2980 30272 -2968 30306
rect -3026 30238 -2968 30272
rect -3026 30204 -3014 30238
rect -2980 30204 -2968 30238
rect -3026 30170 -2968 30204
rect -3026 30136 -3014 30170
rect -2980 30136 -2968 30170
rect -3026 30102 -2968 30136
rect -3026 30068 -3014 30102
rect -2980 30068 -2968 30102
rect -3026 30034 -2968 30068
rect -3026 30000 -3014 30034
rect -2980 30000 -2968 30034
rect -3026 29959 -2968 30000
rect -2868 30918 -2810 30959
rect -2868 30884 -2856 30918
rect -2822 30884 -2810 30918
rect -2868 30850 -2810 30884
rect -2868 30816 -2856 30850
rect -2822 30816 -2810 30850
rect -2868 30782 -2810 30816
rect -2868 30748 -2856 30782
rect -2822 30748 -2810 30782
rect -2868 30714 -2810 30748
rect -2868 30680 -2856 30714
rect -2822 30680 -2810 30714
rect -2868 30646 -2810 30680
rect -2868 30612 -2856 30646
rect -2822 30612 -2810 30646
rect -2868 30578 -2810 30612
rect -2868 30544 -2856 30578
rect -2822 30544 -2810 30578
rect -2868 30510 -2810 30544
rect -2868 30476 -2856 30510
rect -2822 30476 -2810 30510
rect -2868 30442 -2810 30476
rect -2868 30408 -2856 30442
rect -2822 30408 -2810 30442
rect -2868 30374 -2810 30408
rect -2868 30340 -2856 30374
rect -2822 30340 -2810 30374
rect -2868 30306 -2810 30340
rect -2868 30272 -2856 30306
rect -2822 30272 -2810 30306
rect -2868 30238 -2810 30272
rect -2868 30204 -2856 30238
rect -2822 30204 -2810 30238
rect -2868 30170 -2810 30204
rect -2868 30136 -2856 30170
rect -2822 30136 -2810 30170
rect -2868 30102 -2810 30136
rect -2868 30068 -2856 30102
rect -2822 30068 -2810 30102
rect -2868 30034 -2810 30068
rect -2868 30000 -2856 30034
rect -2822 30000 -2810 30034
rect -2868 29959 -2810 30000
rect -2710 30918 -2652 30959
rect -2710 30884 -2698 30918
rect -2664 30884 -2652 30918
rect -2710 30850 -2652 30884
rect -2710 30816 -2698 30850
rect -2664 30816 -2652 30850
rect -2710 30782 -2652 30816
rect -2710 30748 -2698 30782
rect -2664 30748 -2652 30782
rect -2710 30714 -2652 30748
rect -2710 30680 -2698 30714
rect -2664 30680 -2652 30714
rect -2710 30646 -2652 30680
rect -2710 30612 -2698 30646
rect -2664 30612 -2652 30646
rect -2710 30578 -2652 30612
rect -2710 30544 -2698 30578
rect -2664 30544 -2652 30578
rect -2710 30510 -2652 30544
rect -2710 30476 -2698 30510
rect -2664 30476 -2652 30510
rect -2710 30442 -2652 30476
rect -2710 30408 -2698 30442
rect -2664 30408 -2652 30442
rect -2710 30374 -2652 30408
rect -2710 30340 -2698 30374
rect -2664 30340 -2652 30374
rect -2710 30306 -2652 30340
rect -2710 30272 -2698 30306
rect -2664 30272 -2652 30306
rect -2710 30238 -2652 30272
rect -2710 30204 -2698 30238
rect -2664 30204 -2652 30238
rect -2710 30170 -2652 30204
rect -2710 30136 -2698 30170
rect -2664 30136 -2652 30170
rect -2710 30102 -2652 30136
rect -2710 30068 -2698 30102
rect -2664 30068 -2652 30102
rect -2710 30034 -2652 30068
rect -2710 30000 -2698 30034
rect -2664 30000 -2652 30034
rect -2710 29959 -2652 30000
rect -2552 30918 -2494 30959
rect -2552 30884 -2540 30918
rect -2506 30884 -2494 30918
rect -2552 30850 -2494 30884
rect -2552 30816 -2540 30850
rect -2506 30816 -2494 30850
rect -2552 30782 -2494 30816
rect -2552 30748 -2540 30782
rect -2506 30748 -2494 30782
rect -2552 30714 -2494 30748
rect -2552 30680 -2540 30714
rect -2506 30680 -2494 30714
rect -2552 30646 -2494 30680
rect -2552 30612 -2540 30646
rect -2506 30612 -2494 30646
rect -2552 30578 -2494 30612
rect -2552 30544 -2540 30578
rect -2506 30544 -2494 30578
rect -2552 30510 -2494 30544
rect -2552 30476 -2540 30510
rect -2506 30476 -2494 30510
rect -2552 30442 -2494 30476
rect -2552 30408 -2540 30442
rect -2506 30408 -2494 30442
rect -2552 30374 -2494 30408
rect -2552 30340 -2540 30374
rect -2506 30340 -2494 30374
rect -2552 30306 -2494 30340
rect -2552 30272 -2540 30306
rect -2506 30272 -2494 30306
rect -2552 30238 -2494 30272
rect -2552 30204 -2540 30238
rect -2506 30204 -2494 30238
rect -2552 30170 -2494 30204
rect -2552 30136 -2540 30170
rect -2506 30136 -2494 30170
rect -2552 30102 -2494 30136
rect -2552 30068 -2540 30102
rect -2506 30068 -2494 30102
rect -2552 30034 -2494 30068
rect -2552 30000 -2540 30034
rect -2506 30000 -2494 30034
rect -2552 29959 -2494 30000
rect -2394 30918 -2336 30959
rect -2394 30884 -2382 30918
rect -2348 30884 -2336 30918
rect -2394 30850 -2336 30884
rect -2394 30816 -2382 30850
rect -2348 30816 -2336 30850
rect -2394 30782 -2336 30816
rect -2394 30748 -2382 30782
rect -2348 30748 -2336 30782
rect -2394 30714 -2336 30748
rect -2394 30680 -2382 30714
rect -2348 30680 -2336 30714
rect -2394 30646 -2336 30680
rect -2394 30612 -2382 30646
rect -2348 30612 -2336 30646
rect -2394 30578 -2336 30612
rect -2394 30544 -2382 30578
rect -2348 30544 -2336 30578
rect -2394 30510 -2336 30544
rect -2394 30476 -2382 30510
rect -2348 30476 -2336 30510
rect -2394 30442 -2336 30476
rect -2394 30408 -2382 30442
rect -2348 30408 -2336 30442
rect -2394 30374 -2336 30408
rect -2394 30340 -2382 30374
rect -2348 30340 -2336 30374
rect -2394 30306 -2336 30340
rect -2394 30272 -2382 30306
rect -2348 30272 -2336 30306
rect -2394 30238 -2336 30272
rect -2394 30204 -2382 30238
rect -2348 30204 -2336 30238
rect -2394 30170 -2336 30204
rect -2394 30136 -2382 30170
rect -2348 30136 -2336 30170
rect -2394 30102 -2336 30136
rect -2394 30068 -2382 30102
rect -2348 30068 -2336 30102
rect -2394 30034 -2336 30068
rect -2394 30000 -2382 30034
rect -2348 30000 -2336 30034
rect -2394 29959 -2336 30000
rect -2236 30918 -2178 30959
rect -2236 30884 -2224 30918
rect -2190 30884 -2178 30918
rect -2236 30850 -2178 30884
rect -2236 30816 -2224 30850
rect -2190 30816 -2178 30850
rect -2236 30782 -2178 30816
rect -2236 30748 -2224 30782
rect -2190 30748 -2178 30782
rect -2236 30714 -2178 30748
rect -2236 30680 -2224 30714
rect -2190 30680 -2178 30714
rect -2236 30646 -2178 30680
rect -2236 30612 -2224 30646
rect -2190 30612 -2178 30646
rect -2236 30578 -2178 30612
rect -2236 30544 -2224 30578
rect -2190 30544 -2178 30578
rect -2236 30510 -2178 30544
rect -2236 30476 -2224 30510
rect -2190 30476 -2178 30510
rect -2236 30442 -2178 30476
rect -2236 30408 -2224 30442
rect -2190 30408 -2178 30442
rect -2236 30374 -2178 30408
rect -2236 30340 -2224 30374
rect -2190 30340 -2178 30374
rect -2236 30306 -2178 30340
rect -2236 30272 -2224 30306
rect -2190 30272 -2178 30306
rect -2236 30238 -2178 30272
rect -2236 30204 -2224 30238
rect -2190 30204 -2178 30238
rect -2236 30170 -2178 30204
rect -2236 30136 -2224 30170
rect -2190 30136 -2178 30170
rect -2236 30102 -2178 30136
rect -2236 30068 -2224 30102
rect -2190 30068 -2178 30102
rect -2236 30034 -2178 30068
rect -2236 30000 -2224 30034
rect -2190 30000 -2178 30034
rect -2236 29959 -2178 30000
rect -2078 30918 -2020 30959
rect -2078 30884 -2066 30918
rect -2032 30884 -2020 30918
rect -2078 30850 -2020 30884
rect -2078 30816 -2066 30850
rect -2032 30816 -2020 30850
rect -2078 30782 -2020 30816
rect -2078 30748 -2066 30782
rect -2032 30748 -2020 30782
rect -2078 30714 -2020 30748
rect -2078 30680 -2066 30714
rect -2032 30680 -2020 30714
rect -2078 30646 -2020 30680
rect -2078 30612 -2066 30646
rect -2032 30612 -2020 30646
rect -2078 30578 -2020 30612
rect -2078 30544 -2066 30578
rect -2032 30544 -2020 30578
rect -2078 30510 -2020 30544
rect -2078 30476 -2066 30510
rect -2032 30476 -2020 30510
rect -2078 30442 -2020 30476
rect -2078 30408 -2066 30442
rect -2032 30408 -2020 30442
rect -2078 30374 -2020 30408
rect -2078 30340 -2066 30374
rect -2032 30340 -2020 30374
rect -2078 30306 -2020 30340
rect -2078 30272 -2066 30306
rect -2032 30272 -2020 30306
rect -2078 30238 -2020 30272
rect -2078 30204 -2066 30238
rect -2032 30204 -2020 30238
rect -2078 30170 -2020 30204
rect -2078 30136 -2066 30170
rect -2032 30136 -2020 30170
rect -2078 30102 -2020 30136
rect -2078 30068 -2066 30102
rect -2032 30068 -2020 30102
rect -2078 30034 -2020 30068
rect -2078 30000 -2066 30034
rect -2032 30000 -2020 30034
rect -2078 29959 -2020 30000
rect -1920 30918 -1862 30959
rect -1920 30884 -1908 30918
rect -1874 30884 -1862 30918
rect -1920 30850 -1862 30884
rect -1920 30816 -1908 30850
rect -1874 30816 -1862 30850
rect -1920 30782 -1862 30816
rect -1920 30748 -1908 30782
rect -1874 30748 -1862 30782
rect -1920 30714 -1862 30748
rect -1920 30680 -1908 30714
rect -1874 30680 -1862 30714
rect -1920 30646 -1862 30680
rect -1920 30612 -1908 30646
rect -1874 30612 -1862 30646
rect -1920 30578 -1862 30612
rect -1920 30544 -1908 30578
rect -1874 30544 -1862 30578
rect -1920 30510 -1862 30544
rect -1920 30476 -1908 30510
rect -1874 30476 -1862 30510
rect -1920 30442 -1862 30476
rect -1920 30408 -1908 30442
rect -1874 30408 -1862 30442
rect -1920 30374 -1862 30408
rect -1920 30340 -1908 30374
rect -1874 30340 -1862 30374
rect -1920 30306 -1862 30340
rect -1920 30272 -1908 30306
rect -1874 30272 -1862 30306
rect -1920 30238 -1862 30272
rect -1920 30204 -1908 30238
rect -1874 30204 -1862 30238
rect -1920 30170 -1862 30204
rect -1920 30136 -1908 30170
rect -1874 30136 -1862 30170
rect -1920 30102 -1862 30136
rect -1920 30068 -1908 30102
rect -1874 30068 -1862 30102
rect -1920 30034 -1862 30068
rect -1920 30000 -1908 30034
rect -1874 30000 -1862 30034
rect -1920 29959 -1862 30000
rect -1762 30918 -1704 30959
rect -1762 30884 -1750 30918
rect -1716 30884 -1704 30918
rect -1762 30850 -1704 30884
rect -1762 30816 -1750 30850
rect -1716 30816 -1704 30850
rect -1762 30782 -1704 30816
rect -1762 30748 -1750 30782
rect -1716 30748 -1704 30782
rect -1762 30714 -1704 30748
rect -1762 30680 -1750 30714
rect -1716 30680 -1704 30714
rect -1762 30646 -1704 30680
rect -1762 30612 -1750 30646
rect -1716 30612 -1704 30646
rect -1762 30578 -1704 30612
rect -1762 30544 -1750 30578
rect -1716 30544 -1704 30578
rect -1762 30510 -1704 30544
rect -1762 30476 -1750 30510
rect -1716 30476 -1704 30510
rect -1762 30442 -1704 30476
rect -1762 30408 -1750 30442
rect -1716 30408 -1704 30442
rect -1762 30374 -1704 30408
rect -1762 30340 -1750 30374
rect -1716 30340 -1704 30374
rect -1762 30306 -1704 30340
rect -1762 30272 -1750 30306
rect -1716 30272 -1704 30306
rect -1762 30238 -1704 30272
rect -1762 30204 -1750 30238
rect -1716 30204 -1704 30238
rect -1762 30170 -1704 30204
rect -1762 30136 -1750 30170
rect -1716 30136 -1704 30170
rect -1762 30102 -1704 30136
rect -1762 30068 -1750 30102
rect -1716 30068 -1704 30102
rect -1762 30034 -1704 30068
rect -1762 30000 -1750 30034
rect -1716 30000 -1704 30034
rect -1762 29959 -1704 30000
rect -1604 30918 -1546 30959
rect -1604 30884 -1592 30918
rect -1558 30884 -1546 30918
rect -1604 30850 -1546 30884
rect -1604 30816 -1592 30850
rect -1558 30816 -1546 30850
rect -1604 30782 -1546 30816
rect -1604 30748 -1592 30782
rect -1558 30748 -1546 30782
rect -1604 30714 -1546 30748
rect -1604 30680 -1592 30714
rect -1558 30680 -1546 30714
rect -1604 30646 -1546 30680
rect -1604 30612 -1592 30646
rect -1558 30612 -1546 30646
rect -1604 30578 -1546 30612
rect -1604 30544 -1592 30578
rect -1558 30544 -1546 30578
rect -1604 30510 -1546 30544
rect -1604 30476 -1592 30510
rect -1558 30476 -1546 30510
rect -1604 30442 -1546 30476
rect -1604 30408 -1592 30442
rect -1558 30408 -1546 30442
rect -1604 30374 -1546 30408
rect -1604 30340 -1592 30374
rect -1558 30340 -1546 30374
rect -1604 30306 -1546 30340
rect -1604 30272 -1592 30306
rect -1558 30272 -1546 30306
rect -1604 30238 -1546 30272
rect -1604 30204 -1592 30238
rect -1558 30204 -1546 30238
rect -1604 30170 -1546 30204
rect -1604 30136 -1592 30170
rect -1558 30136 -1546 30170
rect -1604 30102 -1546 30136
rect -1604 30068 -1592 30102
rect -1558 30068 -1546 30102
rect -1604 30034 -1546 30068
rect -1604 30000 -1592 30034
rect -1558 30000 -1546 30034
rect -1604 29959 -1546 30000
rect -1446 30918 -1388 30959
rect -1446 30884 -1434 30918
rect -1400 30884 -1388 30918
rect -1446 30850 -1388 30884
rect -1446 30816 -1434 30850
rect -1400 30816 -1388 30850
rect -1446 30782 -1388 30816
rect -1446 30748 -1434 30782
rect -1400 30748 -1388 30782
rect -1446 30714 -1388 30748
rect -1446 30680 -1434 30714
rect -1400 30680 -1388 30714
rect -1446 30646 -1388 30680
rect -1446 30612 -1434 30646
rect -1400 30612 -1388 30646
rect -1446 30578 -1388 30612
rect -1446 30544 -1434 30578
rect -1400 30544 -1388 30578
rect -1446 30510 -1388 30544
rect -1446 30476 -1434 30510
rect -1400 30476 -1388 30510
rect -1446 30442 -1388 30476
rect -1446 30408 -1434 30442
rect -1400 30408 -1388 30442
rect -1446 30374 -1388 30408
rect -1446 30340 -1434 30374
rect -1400 30340 -1388 30374
rect -1446 30306 -1388 30340
rect -1446 30272 -1434 30306
rect -1400 30272 -1388 30306
rect -1446 30238 -1388 30272
rect -1446 30204 -1434 30238
rect -1400 30204 -1388 30238
rect -1446 30170 -1388 30204
rect -1446 30136 -1434 30170
rect -1400 30136 -1388 30170
rect -1446 30102 -1388 30136
rect -1446 30068 -1434 30102
rect -1400 30068 -1388 30102
rect -1446 30034 -1388 30068
rect -1446 30000 -1434 30034
rect -1400 30000 -1388 30034
rect -1446 29959 -1388 30000
rect -1288 30918 -1230 30959
rect -1288 30884 -1276 30918
rect -1242 30884 -1230 30918
rect -1288 30850 -1230 30884
rect -1288 30816 -1276 30850
rect -1242 30816 -1230 30850
rect -1288 30782 -1230 30816
rect -1288 30748 -1276 30782
rect -1242 30748 -1230 30782
rect -1288 30714 -1230 30748
rect -1288 30680 -1276 30714
rect -1242 30680 -1230 30714
rect -1288 30646 -1230 30680
rect -1288 30612 -1276 30646
rect -1242 30612 -1230 30646
rect -1288 30578 -1230 30612
rect -1288 30544 -1276 30578
rect -1242 30544 -1230 30578
rect -1288 30510 -1230 30544
rect -1288 30476 -1276 30510
rect -1242 30476 -1230 30510
rect -1288 30442 -1230 30476
rect -1288 30408 -1276 30442
rect -1242 30408 -1230 30442
rect -1288 30374 -1230 30408
rect -1288 30340 -1276 30374
rect -1242 30340 -1230 30374
rect -1288 30306 -1230 30340
rect -1288 30272 -1276 30306
rect -1242 30272 -1230 30306
rect -1288 30238 -1230 30272
rect -1288 30204 -1276 30238
rect -1242 30204 -1230 30238
rect -1288 30170 -1230 30204
rect -1288 30136 -1276 30170
rect -1242 30136 -1230 30170
rect -1288 30102 -1230 30136
rect -1288 30068 -1276 30102
rect -1242 30068 -1230 30102
rect -1288 30034 -1230 30068
rect -1288 30000 -1276 30034
rect -1242 30000 -1230 30034
rect -1288 29959 -1230 30000
rect -1130 30918 -1072 30959
rect -1130 30884 -1118 30918
rect -1084 30884 -1072 30918
rect -1130 30850 -1072 30884
rect -1130 30816 -1118 30850
rect -1084 30816 -1072 30850
rect -1130 30782 -1072 30816
rect -1130 30748 -1118 30782
rect -1084 30748 -1072 30782
rect -1130 30714 -1072 30748
rect -1130 30680 -1118 30714
rect -1084 30680 -1072 30714
rect -1130 30646 -1072 30680
rect -1130 30612 -1118 30646
rect -1084 30612 -1072 30646
rect -1130 30578 -1072 30612
rect -1130 30544 -1118 30578
rect -1084 30544 -1072 30578
rect -1130 30510 -1072 30544
rect -1130 30476 -1118 30510
rect -1084 30476 -1072 30510
rect -1130 30442 -1072 30476
rect -1130 30408 -1118 30442
rect -1084 30408 -1072 30442
rect -1130 30374 -1072 30408
rect -1130 30340 -1118 30374
rect -1084 30340 -1072 30374
rect -1130 30306 -1072 30340
rect -1130 30272 -1118 30306
rect -1084 30272 -1072 30306
rect -1130 30238 -1072 30272
rect -1130 30204 -1118 30238
rect -1084 30204 -1072 30238
rect -1130 30170 -1072 30204
rect -1130 30136 -1118 30170
rect -1084 30136 -1072 30170
rect -1130 30102 -1072 30136
rect -1130 30068 -1118 30102
rect -1084 30068 -1072 30102
rect -1130 30034 -1072 30068
rect -1130 30000 -1118 30034
rect -1084 30000 -1072 30034
rect -1130 29959 -1072 30000
rect -972 30918 -914 30959
rect -972 30884 -960 30918
rect -926 30884 -914 30918
rect -972 30850 -914 30884
rect -972 30816 -960 30850
rect -926 30816 -914 30850
rect -972 30782 -914 30816
rect -972 30748 -960 30782
rect -926 30748 -914 30782
rect -972 30714 -914 30748
rect -972 30680 -960 30714
rect -926 30680 -914 30714
rect -972 30646 -914 30680
rect -972 30612 -960 30646
rect -926 30612 -914 30646
rect -972 30578 -914 30612
rect -972 30544 -960 30578
rect -926 30544 -914 30578
rect -972 30510 -914 30544
rect -972 30476 -960 30510
rect -926 30476 -914 30510
rect -972 30442 -914 30476
rect -972 30408 -960 30442
rect -926 30408 -914 30442
rect -972 30374 -914 30408
rect -972 30340 -960 30374
rect -926 30340 -914 30374
rect -972 30306 -914 30340
rect -972 30272 -960 30306
rect -926 30272 -914 30306
rect -972 30238 -914 30272
rect -972 30204 -960 30238
rect -926 30204 -914 30238
rect -972 30170 -914 30204
rect -972 30136 -960 30170
rect -926 30136 -914 30170
rect -972 30102 -914 30136
rect -972 30068 -960 30102
rect -926 30068 -914 30102
rect -972 30034 -914 30068
rect -972 30000 -960 30034
rect -926 30000 -914 30034
rect -972 29959 -914 30000
rect -814 30918 -756 30959
rect -814 30884 -802 30918
rect -768 30884 -756 30918
rect -814 30850 -756 30884
rect -814 30816 -802 30850
rect -768 30816 -756 30850
rect -814 30782 -756 30816
rect -814 30748 -802 30782
rect -768 30748 -756 30782
rect -814 30714 -756 30748
rect -814 30680 -802 30714
rect -768 30680 -756 30714
rect -814 30646 -756 30680
rect -814 30612 -802 30646
rect -768 30612 -756 30646
rect -814 30578 -756 30612
rect -814 30544 -802 30578
rect -768 30544 -756 30578
rect -814 30510 -756 30544
rect -814 30476 -802 30510
rect -768 30476 -756 30510
rect -814 30442 -756 30476
rect -814 30408 -802 30442
rect -768 30408 -756 30442
rect -814 30374 -756 30408
rect -814 30340 -802 30374
rect -768 30340 -756 30374
rect -814 30306 -756 30340
rect -814 30272 -802 30306
rect -768 30272 -756 30306
rect -814 30238 -756 30272
rect -814 30204 -802 30238
rect -768 30204 -756 30238
rect -814 30170 -756 30204
rect -814 30136 -802 30170
rect -768 30136 -756 30170
rect -814 30102 -756 30136
rect -814 30068 -802 30102
rect -768 30068 -756 30102
rect -814 30034 -756 30068
rect -814 30000 -802 30034
rect -768 30000 -756 30034
rect -814 29959 -756 30000
rect -656 30918 -598 30959
rect -656 30884 -644 30918
rect -610 30884 -598 30918
rect -656 30850 -598 30884
rect -656 30816 -644 30850
rect -610 30816 -598 30850
rect -656 30782 -598 30816
rect -656 30748 -644 30782
rect -610 30748 -598 30782
rect -656 30714 -598 30748
rect -656 30680 -644 30714
rect -610 30680 -598 30714
rect -656 30646 -598 30680
rect -656 30612 -644 30646
rect -610 30612 -598 30646
rect -656 30578 -598 30612
rect -656 30544 -644 30578
rect -610 30544 -598 30578
rect -656 30510 -598 30544
rect -656 30476 -644 30510
rect -610 30476 -598 30510
rect -656 30442 -598 30476
rect -656 30408 -644 30442
rect -610 30408 -598 30442
rect -656 30374 -598 30408
rect -656 30340 -644 30374
rect -610 30340 -598 30374
rect -656 30306 -598 30340
rect -656 30272 -644 30306
rect -610 30272 -598 30306
rect -656 30238 -598 30272
rect -656 30204 -644 30238
rect -610 30204 -598 30238
rect -656 30170 -598 30204
rect -656 30136 -644 30170
rect -610 30136 -598 30170
rect -656 30102 -598 30136
rect -656 30068 -644 30102
rect -610 30068 -598 30102
rect -656 30034 -598 30068
rect -656 30000 -644 30034
rect -610 30000 -598 30034
rect -656 29959 -598 30000
rect -498 30918 -440 30959
rect -498 30884 -486 30918
rect -452 30884 -440 30918
rect -498 30850 -440 30884
rect -498 30816 -486 30850
rect -452 30816 -440 30850
rect -498 30782 -440 30816
rect -498 30748 -486 30782
rect -452 30748 -440 30782
rect -498 30714 -440 30748
rect -498 30680 -486 30714
rect -452 30680 -440 30714
rect -498 30646 -440 30680
rect -498 30612 -486 30646
rect -452 30612 -440 30646
rect -498 30578 -440 30612
rect -498 30544 -486 30578
rect -452 30544 -440 30578
rect -498 30510 -440 30544
rect -498 30476 -486 30510
rect -452 30476 -440 30510
rect -498 30442 -440 30476
rect -498 30408 -486 30442
rect -452 30408 -440 30442
rect -498 30374 -440 30408
rect -498 30340 -486 30374
rect -452 30340 -440 30374
rect -498 30306 -440 30340
rect -498 30272 -486 30306
rect -452 30272 -440 30306
rect -498 30238 -440 30272
rect -498 30204 -486 30238
rect -452 30204 -440 30238
rect -498 30170 -440 30204
rect -498 30136 -486 30170
rect -452 30136 -440 30170
rect -498 30102 -440 30136
rect -498 30068 -486 30102
rect -452 30068 -440 30102
rect -498 30034 -440 30068
rect -498 30000 -486 30034
rect -452 30000 -440 30034
rect -498 29959 -440 30000
rect -340 30918 -282 30959
rect -340 30884 -328 30918
rect -294 30884 -282 30918
rect -340 30850 -282 30884
rect -340 30816 -328 30850
rect -294 30816 -282 30850
rect -340 30782 -282 30816
rect -340 30748 -328 30782
rect -294 30748 -282 30782
rect -340 30714 -282 30748
rect -340 30680 -328 30714
rect -294 30680 -282 30714
rect -340 30646 -282 30680
rect -340 30612 -328 30646
rect -294 30612 -282 30646
rect -340 30578 -282 30612
rect -340 30544 -328 30578
rect -294 30544 -282 30578
rect -340 30510 -282 30544
rect -340 30476 -328 30510
rect -294 30476 -282 30510
rect -340 30442 -282 30476
rect -340 30408 -328 30442
rect -294 30408 -282 30442
rect -340 30374 -282 30408
rect -340 30340 -328 30374
rect -294 30340 -282 30374
rect -340 30306 -282 30340
rect -340 30272 -328 30306
rect -294 30272 -282 30306
rect -340 30238 -282 30272
rect -340 30204 -328 30238
rect -294 30204 -282 30238
rect -340 30170 -282 30204
rect -340 30136 -328 30170
rect -294 30136 -282 30170
rect -340 30102 -282 30136
rect -340 30068 -328 30102
rect -294 30068 -282 30102
rect -340 30034 -282 30068
rect -340 30000 -328 30034
rect -294 30000 -282 30034
rect -340 29959 -282 30000
rect -182 30918 -124 30959
rect -182 30884 -170 30918
rect -136 30884 -124 30918
rect -182 30850 -124 30884
rect -182 30816 -170 30850
rect -136 30816 -124 30850
rect -182 30782 -124 30816
rect -182 30748 -170 30782
rect -136 30748 -124 30782
rect -182 30714 -124 30748
rect -182 30680 -170 30714
rect -136 30680 -124 30714
rect -182 30646 -124 30680
rect -182 30612 -170 30646
rect -136 30612 -124 30646
rect -182 30578 -124 30612
rect -182 30544 -170 30578
rect -136 30544 -124 30578
rect -182 30510 -124 30544
rect -182 30476 -170 30510
rect -136 30476 -124 30510
rect -182 30442 -124 30476
rect -182 30408 -170 30442
rect -136 30408 -124 30442
rect -182 30374 -124 30408
rect -182 30340 -170 30374
rect -136 30340 -124 30374
rect -182 30306 -124 30340
rect -182 30272 -170 30306
rect -136 30272 -124 30306
rect -182 30238 -124 30272
rect -182 30204 -170 30238
rect -136 30204 -124 30238
rect -182 30170 -124 30204
rect -182 30136 -170 30170
rect -136 30136 -124 30170
rect -182 30102 -124 30136
rect -182 30068 -170 30102
rect -136 30068 -124 30102
rect -182 30034 -124 30068
rect -182 30000 -170 30034
rect -136 30000 -124 30034
rect -182 29959 -124 30000
rect -24 30918 34 30959
rect -24 30884 -12 30918
rect 22 30884 34 30918
rect -24 30850 34 30884
rect -24 30816 -12 30850
rect 22 30816 34 30850
rect -24 30782 34 30816
rect -24 30748 -12 30782
rect 22 30748 34 30782
rect -24 30714 34 30748
rect -24 30680 -12 30714
rect 22 30680 34 30714
rect -24 30646 34 30680
rect -24 30612 -12 30646
rect 22 30612 34 30646
rect -24 30578 34 30612
rect -24 30544 -12 30578
rect 22 30544 34 30578
rect -24 30510 34 30544
rect -24 30476 -12 30510
rect 22 30476 34 30510
rect -24 30442 34 30476
rect -24 30408 -12 30442
rect 22 30408 34 30442
rect -24 30374 34 30408
rect -24 30340 -12 30374
rect 22 30340 34 30374
rect -24 30306 34 30340
rect -24 30272 -12 30306
rect 22 30272 34 30306
rect -24 30238 34 30272
rect -24 30204 -12 30238
rect 22 30204 34 30238
rect -24 30170 34 30204
rect -24 30136 -12 30170
rect 22 30136 34 30170
rect -24 30102 34 30136
rect -24 30068 -12 30102
rect 22 30068 34 30102
rect -24 30034 34 30068
rect -24 30000 -12 30034
rect 22 30000 34 30034
rect -24 29959 34 30000
rect 134 30918 192 30959
rect 134 30884 146 30918
rect 180 30884 192 30918
rect 134 30850 192 30884
rect 134 30816 146 30850
rect 180 30816 192 30850
rect 134 30782 192 30816
rect 134 30748 146 30782
rect 180 30748 192 30782
rect 134 30714 192 30748
rect 134 30680 146 30714
rect 180 30680 192 30714
rect 134 30646 192 30680
rect 134 30612 146 30646
rect 180 30612 192 30646
rect 134 30578 192 30612
rect 134 30544 146 30578
rect 180 30544 192 30578
rect 134 30510 192 30544
rect 134 30476 146 30510
rect 180 30476 192 30510
rect 134 30442 192 30476
rect 134 30408 146 30442
rect 180 30408 192 30442
rect 134 30374 192 30408
rect 134 30340 146 30374
rect 180 30340 192 30374
rect 134 30306 192 30340
rect 134 30272 146 30306
rect 180 30272 192 30306
rect 134 30238 192 30272
rect 134 30204 146 30238
rect 180 30204 192 30238
rect 134 30170 192 30204
rect 134 30136 146 30170
rect 180 30136 192 30170
rect 134 30102 192 30136
rect 134 30068 146 30102
rect 180 30068 192 30102
rect 134 30034 192 30068
rect 134 30000 146 30034
rect 180 30000 192 30034
rect 134 29959 192 30000
rect 292 30918 350 30959
rect 292 30884 304 30918
rect 338 30884 350 30918
rect 292 30850 350 30884
rect 292 30816 304 30850
rect 338 30816 350 30850
rect 292 30782 350 30816
rect 292 30748 304 30782
rect 338 30748 350 30782
rect 292 30714 350 30748
rect 292 30680 304 30714
rect 338 30680 350 30714
rect 292 30646 350 30680
rect 292 30612 304 30646
rect 338 30612 350 30646
rect 292 30578 350 30612
rect 292 30544 304 30578
rect 338 30544 350 30578
rect 292 30510 350 30544
rect 292 30476 304 30510
rect 338 30476 350 30510
rect 292 30442 350 30476
rect 292 30408 304 30442
rect 338 30408 350 30442
rect 292 30374 350 30408
rect 292 30340 304 30374
rect 338 30340 350 30374
rect 292 30306 350 30340
rect 292 30272 304 30306
rect 338 30272 350 30306
rect 292 30238 350 30272
rect 292 30204 304 30238
rect 338 30204 350 30238
rect 292 30170 350 30204
rect 292 30136 304 30170
rect 338 30136 350 30170
rect 292 30102 350 30136
rect 292 30068 304 30102
rect 338 30068 350 30102
rect 292 30034 350 30068
rect 292 30000 304 30034
rect 338 30000 350 30034
rect 292 29959 350 30000
rect 450 30918 508 30959
rect 450 30884 462 30918
rect 496 30884 508 30918
rect 450 30850 508 30884
rect 450 30816 462 30850
rect 496 30816 508 30850
rect 450 30782 508 30816
rect 450 30748 462 30782
rect 496 30748 508 30782
rect 450 30714 508 30748
rect 450 30680 462 30714
rect 496 30680 508 30714
rect 450 30646 508 30680
rect 450 30612 462 30646
rect 496 30612 508 30646
rect 450 30578 508 30612
rect 450 30544 462 30578
rect 496 30544 508 30578
rect 450 30510 508 30544
rect 450 30476 462 30510
rect 496 30476 508 30510
rect 450 30442 508 30476
rect 450 30408 462 30442
rect 496 30408 508 30442
rect 450 30374 508 30408
rect 450 30340 462 30374
rect 496 30340 508 30374
rect 450 30306 508 30340
rect 450 30272 462 30306
rect 496 30272 508 30306
rect 450 30238 508 30272
rect 450 30204 462 30238
rect 496 30204 508 30238
rect 450 30170 508 30204
rect 450 30136 462 30170
rect 496 30136 508 30170
rect 450 30102 508 30136
rect 450 30068 462 30102
rect 496 30068 508 30102
rect 450 30034 508 30068
rect 450 30000 462 30034
rect 496 30000 508 30034
rect 450 29959 508 30000
rect 608 30918 666 30959
rect 608 30884 620 30918
rect 654 30884 666 30918
rect 608 30850 666 30884
rect 608 30816 620 30850
rect 654 30816 666 30850
rect 608 30782 666 30816
rect 608 30748 620 30782
rect 654 30748 666 30782
rect 608 30714 666 30748
rect 608 30680 620 30714
rect 654 30680 666 30714
rect 608 30646 666 30680
rect 608 30612 620 30646
rect 654 30612 666 30646
rect 608 30578 666 30612
rect 608 30544 620 30578
rect 654 30544 666 30578
rect 608 30510 666 30544
rect 608 30476 620 30510
rect 654 30476 666 30510
rect 608 30442 666 30476
rect 608 30408 620 30442
rect 654 30408 666 30442
rect 608 30374 666 30408
rect 608 30340 620 30374
rect 654 30340 666 30374
rect 608 30306 666 30340
rect 608 30272 620 30306
rect 654 30272 666 30306
rect 608 30238 666 30272
rect 608 30204 620 30238
rect 654 30204 666 30238
rect 608 30170 666 30204
rect 608 30136 620 30170
rect 654 30136 666 30170
rect 608 30102 666 30136
rect 608 30068 620 30102
rect 654 30068 666 30102
rect 608 30034 666 30068
rect 608 30000 620 30034
rect 654 30000 666 30034
rect 608 29959 666 30000
rect 766 30918 824 30959
rect 766 30884 778 30918
rect 812 30884 824 30918
rect 766 30850 824 30884
rect 766 30816 778 30850
rect 812 30816 824 30850
rect 766 30782 824 30816
rect 766 30748 778 30782
rect 812 30748 824 30782
rect 766 30714 824 30748
rect 766 30680 778 30714
rect 812 30680 824 30714
rect 766 30646 824 30680
rect 766 30612 778 30646
rect 812 30612 824 30646
rect 766 30578 824 30612
rect 766 30544 778 30578
rect 812 30544 824 30578
rect 766 30510 824 30544
rect 766 30476 778 30510
rect 812 30476 824 30510
rect 766 30442 824 30476
rect 766 30408 778 30442
rect 812 30408 824 30442
rect 766 30374 824 30408
rect 766 30340 778 30374
rect 812 30340 824 30374
rect 766 30306 824 30340
rect 766 30272 778 30306
rect 812 30272 824 30306
rect 766 30238 824 30272
rect 766 30204 778 30238
rect 812 30204 824 30238
rect 766 30170 824 30204
rect 766 30136 778 30170
rect 812 30136 824 30170
rect 766 30102 824 30136
rect 766 30068 778 30102
rect 812 30068 824 30102
rect 766 30034 824 30068
rect 766 30000 778 30034
rect 812 30000 824 30034
rect 766 29959 824 30000
rect 924 30918 982 30959
rect 924 30884 936 30918
rect 970 30884 982 30918
rect 924 30850 982 30884
rect 924 30816 936 30850
rect 970 30816 982 30850
rect 924 30782 982 30816
rect 924 30748 936 30782
rect 970 30748 982 30782
rect 924 30714 982 30748
rect 924 30680 936 30714
rect 970 30680 982 30714
rect 924 30646 982 30680
rect 924 30612 936 30646
rect 970 30612 982 30646
rect 924 30578 982 30612
rect 924 30544 936 30578
rect 970 30544 982 30578
rect 924 30510 982 30544
rect 924 30476 936 30510
rect 970 30476 982 30510
rect 924 30442 982 30476
rect 924 30408 936 30442
rect 970 30408 982 30442
rect 924 30374 982 30408
rect 924 30340 936 30374
rect 970 30340 982 30374
rect 924 30306 982 30340
rect 924 30272 936 30306
rect 970 30272 982 30306
rect 924 30238 982 30272
rect 924 30204 936 30238
rect 970 30204 982 30238
rect 924 30170 982 30204
rect 924 30136 936 30170
rect 970 30136 982 30170
rect 924 30102 982 30136
rect 924 30068 936 30102
rect 970 30068 982 30102
rect 924 30034 982 30068
rect 924 30000 936 30034
rect 970 30000 982 30034
rect 924 29959 982 30000
rect 1082 30918 1140 30959
rect 1082 30884 1094 30918
rect 1128 30884 1140 30918
rect 1082 30850 1140 30884
rect 1082 30816 1094 30850
rect 1128 30816 1140 30850
rect 1082 30782 1140 30816
rect 1082 30748 1094 30782
rect 1128 30748 1140 30782
rect 1082 30714 1140 30748
rect 1082 30680 1094 30714
rect 1128 30680 1140 30714
rect 1082 30646 1140 30680
rect 1082 30612 1094 30646
rect 1128 30612 1140 30646
rect 1082 30578 1140 30612
rect 1082 30544 1094 30578
rect 1128 30544 1140 30578
rect 1082 30510 1140 30544
rect 1082 30476 1094 30510
rect 1128 30476 1140 30510
rect 1082 30442 1140 30476
rect 1082 30408 1094 30442
rect 1128 30408 1140 30442
rect 1082 30374 1140 30408
rect 1082 30340 1094 30374
rect 1128 30340 1140 30374
rect 1082 30306 1140 30340
rect 1082 30272 1094 30306
rect 1128 30272 1140 30306
rect 1082 30238 1140 30272
rect 1082 30204 1094 30238
rect 1128 30204 1140 30238
rect 1082 30170 1140 30204
rect 1082 30136 1094 30170
rect 1128 30136 1140 30170
rect 1082 30102 1140 30136
rect 1082 30068 1094 30102
rect 1128 30068 1140 30102
rect 1082 30034 1140 30068
rect 1082 30000 1094 30034
rect 1128 30000 1140 30034
rect 1082 29959 1140 30000
rect 1240 30918 1298 30959
rect 1240 30884 1252 30918
rect 1286 30884 1298 30918
rect 1240 30850 1298 30884
rect 1240 30816 1252 30850
rect 1286 30816 1298 30850
rect 1240 30782 1298 30816
rect 1240 30748 1252 30782
rect 1286 30748 1298 30782
rect 1240 30714 1298 30748
rect 1240 30680 1252 30714
rect 1286 30680 1298 30714
rect 1240 30646 1298 30680
rect 1240 30612 1252 30646
rect 1286 30612 1298 30646
rect 1240 30578 1298 30612
rect 1240 30544 1252 30578
rect 1286 30544 1298 30578
rect 1240 30510 1298 30544
rect 1240 30476 1252 30510
rect 1286 30476 1298 30510
rect 1240 30442 1298 30476
rect 1240 30408 1252 30442
rect 1286 30408 1298 30442
rect 1240 30374 1298 30408
rect 1240 30340 1252 30374
rect 1286 30340 1298 30374
rect 1240 30306 1298 30340
rect 1240 30272 1252 30306
rect 1286 30272 1298 30306
rect 1240 30238 1298 30272
rect 1240 30204 1252 30238
rect 1286 30204 1298 30238
rect 1240 30170 1298 30204
rect 1240 30136 1252 30170
rect 1286 30136 1298 30170
rect 1240 30102 1298 30136
rect 1240 30068 1252 30102
rect 1286 30068 1298 30102
rect 1240 30034 1298 30068
rect 1240 30000 1252 30034
rect 1286 30000 1298 30034
rect 1240 29959 1298 30000
rect 1398 30918 1456 30959
rect 1398 30884 1410 30918
rect 1444 30884 1456 30918
rect 1398 30850 1456 30884
rect 1398 30816 1410 30850
rect 1444 30816 1456 30850
rect 1398 30782 1456 30816
rect 1398 30748 1410 30782
rect 1444 30748 1456 30782
rect 1398 30714 1456 30748
rect 1398 30680 1410 30714
rect 1444 30680 1456 30714
rect 1398 30646 1456 30680
rect 1398 30612 1410 30646
rect 1444 30612 1456 30646
rect 1398 30578 1456 30612
rect 1398 30544 1410 30578
rect 1444 30544 1456 30578
rect 1398 30510 1456 30544
rect 1398 30476 1410 30510
rect 1444 30476 1456 30510
rect 1398 30442 1456 30476
rect 1398 30408 1410 30442
rect 1444 30408 1456 30442
rect 1398 30374 1456 30408
rect 1398 30340 1410 30374
rect 1444 30340 1456 30374
rect 1398 30306 1456 30340
rect 1398 30272 1410 30306
rect 1444 30272 1456 30306
rect 1398 30238 1456 30272
rect 1398 30204 1410 30238
rect 1444 30204 1456 30238
rect 1398 30170 1456 30204
rect 1398 30136 1410 30170
rect 1444 30136 1456 30170
rect 1398 30102 1456 30136
rect 1398 30068 1410 30102
rect 1444 30068 1456 30102
rect 1398 30034 1456 30068
rect 1398 30000 1410 30034
rect 1444 30000 1456 30034
rect 1398 29959 1456 30000
rect 1556 30918 1614 30959
rect 1556 30884 1568 30918
rect 1602 30884 1614 30918
rect 1556 30850 1614 30884
rect 1556 30816 1568 30850
rect 1602 30816 1614 30850
rect 1556 30782 1614 30816
rect 1556 30748 1568 30782
rect 1602 30748 1614 30782
rect 1556 30714 1614 30748
rect 1556 30680 1568 30714
rect 1602 30680 1614 30714
rect 1556 30646 1614 30680
rect 1556 30612 1568 30646
rect 1602 30612 1614 30646
rect 1556 30578 1614 30612
rect 1556 30544 1568 30578
rect 1602 30544 1614 30578
rect 1556 30510 1614 30544
rect 1556 30476 1568 30510
rect 1602 30476 1614 30510
rect 1556 30442 1614 30476
rect 1556 30408 1568 30442
rect 1602 30408 1614 30442
rect 1556 30374 1614 30408
rect 1556 30340 1568 30374
rect 1602 30340 1614 30374
rect 1556 30306 1614 30340
rect 1556 30272 1568 30306
rect 1602 30272 1614 30306
rect 1556 30238 1614 30272
rect 1556 30204 1568 30238
rect 1602 30204 1614 30238
rect 1556 30170 1614 30204
rect 1556 30136 1568 30170
rect 1602 30136 1614 30170
rect 1556 30102 1614 30136
rect 1556 30068 1568 30102
rect 1602 30068 1614 30102
rect 1556 30034 1614 30068
rect 1556 30000 1568 30034
rect 1602 30000 1614 30034
rect 1556 29959 1614 30000
rect 1714 30918 1772 30959
rect 1714 30884 1726 30918
rect 1760 30884 1772 30918
rect 1714 30850 1772 30884
rect 1714 30816 1726 30850
rect 1760 30816 1772 30850
rect 1714 30782 1772 30816
rect 1714 30748 1726 30782
rect 1760 30748 1772 30782
rect 1714 30714 1772 30748
rect 1714 30680 1726 30714
rect 1760 30680 1772 30714
rect 1714 30646 1772 30680
rect 1714 30612 1726 30646
rect 1760 30612 1772 30646
rect 1714 30578 1772 30612
rect 1714 30544 1726 30578
rect 1760 30544 1772 30578
rect 1714 30510 1772 30544
rect 1714 30476 1726 30510
rect 1760 30476 1772 30510
rect 1714 30442 1772 30476
rect 1714 30408 1726 30442
rect 1760 30408 1772 30442
rect 1714 30374 1772 30408
rect 1714 30340 1726 30374
rect 1760 30340 1772 30374
rect 1714 30306 1772 30340
rect 1714 30272 1726 30306
rect 1760 30272 1772 30306
rect 1714 30238 1772 30272
rect 1714 30204 1726 30238
rect 1760 30204 1772 30238
rect 1714 30170 1772 30204
rect 1714 30136 1726 30170
rect 1760 30136 1772 30170
rect 1714 30102 1772 30136
rect 1714 30068 1726 30102
rect 1760 30068 1772 30102
rect 1714 30034 1772 30068
rect 1714 30000 1726 30034
rect 1760 30000 1772 30034
rect 1714 29959 1772 30000
rect 1872 30918 1930 30959
rect 1872 30884 1884 30918
rect 1918 30884 1930 30918
rect 1872 30850 1930 30884
rect 1872 30816 1884 30850
rect 1918 30816 1930 30850
rect 1872 30782 1930 30816
rect 1872 30748 1884 30782
rect 1918 30748 1930 30782
rect 1872 30714 1930 30748
rect 1872 30680 1884 30714
rect 1918 30680 1930 30714
rect 1872 30646 1930 30680
rect 1872 30612 1884 30646
rect 1918 30612 1930 30646
rect 1872 30578 1930 30612
rect 1872 30544 1884 30578
rect 1918 30544 1930 30578
rect 1872 30510 1930 30544
rect 1872 30476 1884 30510
rect 1918 30476 1930 30510
rect 1872 30442 1930 30476
rect 1872 30408 1884 30442
rect 1918 30408 1930 30442
rect 1872 30374 1930 30408
rect 1872 30340 1884 30374
rect 1918 30340 1930 30374
rect 1872 30306 1930 30340
rect 1872 30272 1884 30306
rect 1918 30272 1930 30306
rect 1872 30238 1930 30272
rect 1872 30204 1884 30238
rect 1918 30204 1930 30238
rect 1872 30170 1930 30204
rect 1872 30136 1884 30170
rect 1918 30136 1930 30170
rect 1872 30102 1930 30136
rect 1872 30068 1884 30102
rect 1918 30068 1930 30102
rect 1872 30034 1930 30068
rect 1872 30000 1884 30034
rect 1918 30000 1930 30034
rect 1872 29959 1930 30000
rect 2030 30918 2088 30959
rect 2030 30884 2042 30918
rect 2076 30884 2088 30918
rect 2030 30850 2088 30884
rect 2030 30816 2042 30850
rect 2076 30816 2088 30850
rect 2030 30782 2088 30816
rect 2030 30748 2042 30782
rect 2076 30748 2088 30782
rect 2030 30714 2088 30748
rect 2030 30680 2042 30714
rect 2076 30680 2088 30714
rect 2030 30646 2088 30680
rect 2030 30612 2042 30646
rect 2076 30612 2088 30646
rect 2030 30578 2088 30612
rect 2030 30544 2042 30578
rect 2076 30544 2088 30578
rect 2030 30510 2088 30544
rect 2030 30476 2042 30510
rect 2076 30476 2088 30510
rect 2030 30442 2088 30476
rect 2030 30408 2042 30442
rect 2076 30408 2088 30442
rect 2030 30374 2088 30408
rect 2030 30340 2042 30374
rect 2076 30340 2088 30374
rect 2030 30306 2088 30340
rect 2030 30272 2042 30306
rect 2076 30272 2088 30306
rect 2030 30238 2088 30272
rect 2030 30204 2042 30238
rect 2076 30204 2088 30238
rect 2030 30170 2088 30204
rect 2030 30136 2042 30170
rect 2076 30136 2088 30170
rect 2030 30102 2088 30136
rect 2030 30068 2042 30102
rect 2076 30068 2088 30102
rect 2030 30034 2088 30068
rect 2030 30000 2042 30034
rect 2076 30000 2088 30034
rect 2030 29959 2088 30000
rect 2188 30918 2246 30959
rect 2188 30884 2200 30918
rect 2234 30884 2246 30918
rect 2188 30850 2246 30884
rect 2188 30816 2200 30850
rect 2234 30816 2246 30850
rect 2188 30782 2246 30816
rect 2188 30748 2200 30782
rect 2234 30748 2246 30782
rect 2188 30714 2246 30748
rect 2188 30680 2200 30714
rect 2234 30680 2246 30714
rect 2188 30646 2246 30680
rect 2188 30612 2200 30646
rect 2234 30612 2246 30646
rect 2188 30578 2246 30612
rect 2188 30544 2200 30578
rect 2234 30544 2246 30578
rect 2188 30510 2246 30544
rect 2188 30476 2200 30510
rect 2234 30476 2246 30510
rect 2188 30442 2246 30476
rect 2188 30408 2200 30442
rect 2234 30408 2246 30442
rect 2188 30374 2246 30408
rect 2188 30340 2200 30374
rect 2234 30340 2246 30374
rect 2188 30306 2246 30340
rect 2188 30272 2200 30306
rect 2234 30272 2246 30306
rect 2188 30238 2246 30272
rect 2188 30204 2200 30238
rect 2234 30204 2246 30238
rect 2188 30170 2246 30204
rect 2188 30136 2200 30170
rect 2234 30136 2246 30170
rect 2188 30102 2246 30136
rect 2188 30068 2200 30102
rect 2234 30068 2246 30102
rect 2188 30034 2246 30068
rect 2188 30000 2200 30034
rect 2234 30000 2246 30034
rect 2188 29959 2246 30000
rect 2346 30918 2404 30959
rect 2346 30884 2358 30918
rect 2392 30884 2404 30918
rect 2346 30850 2404 30884
rect 2346 30816 2358 30850
rect 2392 30816 2404 30850
rect 2346 30782 2404 30816
rect 2346 30748 2358 30782
rect 2392 30748 2404 30782
rect 2346 30714 2404 30748
rect 2346 30680 2358 30714
rect 2392 30680 2404 30714
rect 2346 30646 2404 30680
rect 2346 30612 2358 30646
rect 2392 30612 2404 30646
rect 2346 30578 2404 30612
rect 2346 30544 2358 30578
rect 2392 30544 2404 30578
rect 2346 30510 2404 30544
rect 2346 30476 2358 30510
rect 2392 30476 2404 30510
rect 2346 30442 2404 30476
rect 2346 30408 2358 30442
rect 2392 30408 2404 30442
rect 2346 30374 2404 30408
rect 2346 30340 2358 30374
rect 2392 30340 2404 30374
rect 2346 30306 2404 30340
rect 2346 30272 2358 30306
rect 2392 30272 2404 30306
rect 2346 30238 2404 30272
rect 2346 30204 2358 30238
rect 2392 30204 2404 30238
rect 2346 30170 2404 30204
rect 2346 30136 2358 30170
rect 2392 30136 2404 30170
rect 2346 30102 2404 30136
rect 2346 30068 2358 30102
rect 2392 30068 2404 30102
rect 2346 30034 2404 30068
rect 2346 30000 2358 30034
rect 2392 30000 2404 30034
rect 2346 29959 2404 30000
rect 2504 30918 2562 30959
rect 2504 30884 2516 30918
rect 2550 30884 2562 30918
rect 2504 30850 2562 30884
rect 2504 30816 2516 30850
rect 2550 30816 2562 30850
rect 2504 30782 2562 30816
rect 2504 30748 2516 30782
rect 2550 30748 2562 30782
rect 2504 30714 2562 30748
rect 2504 30680 2516 30714
rect 2550 30680 2562 30714
rect 2504 30646 2562 30680
rect 2504 30612 2516 30646
rect 2550 30612 2562 30646
rect 2504 30578 2562 30612
rect 2504 30544 2516 30578
rect 2550 30544 2562 30578
rect 2504 30510 2562 30544
rect 2504 30476 2516 30510
rect 2550 30476 2562 30510
rect 2504 30442 2562 30476
rect 2504 30408 2516 30442
rect 2550 30408 2562 30442
rect 2504 30374 2562 30408
rect 2504 30340 2516 30374
rect 2550 30340 2562 30374
rect 2504 30306 2562 30340
rect 2504 30272 2516 30306
rect 2550 30272 2562 30306
rect 2504 30238 2562 30272
rect 2504 30204 2516 30238
rect 2550 30204 2562 30238
rect 2504 30170 2562 30204
rect 2504 30136 2516 30170
rect 2550 30136 2562 30170
rect 2504 30102 2562 30136
rect 2504 30068 2516 30102
rect 2550 30068 2562 30102
rect 2504 30034 2562 30068
rect 2504 30000 2516 30034
rect 2550 30000 2562 30034
rect 2504 29959 2562 30000
rect 2662 30918 2720 30959
rect 2662 30884 2674 30918
rect 2708 30884 2720 30918
rect 2662 30850 2720 30884
rect 2662 30816 2674 30850
rect 2708 30816 2720 30850
rect 2662 30782 2720 30816
rect 2662 30748 2674 30782
rect 2708 30748 2720 30782
rect 2662 30714 2720 30748
rect 2662 30680 2674 30714
rect 2708 30680 2720 30714
rect 2662 30646 2720 30680
rect 2662 30612 2674 30646
rect 2708 30612 2720 30646
rect 2662 30578 2720 30612
rect 2662 30544 2674 30578
rect 2708 30544 2720 30578
rect 2662 30510 2720 30544
rect 2662 30476 2674 30510
rect 2708 30476 2720 30510
rect 2662 30442 2720 30476
rect 2662 30408 2674 30442
rect 2708 30408 2720 30442
rect 2662 30374 2720 30408
rect 2662 30340 2674 30374
rect 2708 30340 2720 30374
rect 2662 30306 2720 30340
rect 2662 30272 2674 30306
rect 2708 30272 2720 30306
rect 2662 30238 2720 30272
rect 2662 30204 2674 30238
rect 2708 30204 2720 30238
rect 2662 30170 2720 30204
rect 2662 30136 2674 30170
rect 2708 30136 2720 30170
rect 2662 30102 2720 30136
rect 2662 30068 2674 30102
rect 2708 30068 2720 30102
rect 2662 30034 2720 30068
rect 2662 30000 2674 30034
rect 2708 30000 2720 30034
rect 2662 29959 2720 30000
rect 2820 30918 2878 30959
rect 2820 30884 2832 30918
rect 2866 30884 2878 30918
rect 2820 30850 2878 30884
rect 2820 30816 2832 30850
rect 2866 30816 2878 30850
rect 2820 30782 2878 30816
rect 2820 30748 2832 30782
rect 2866 30748 2878 30782
rect 2820 30714 2878 30748
rect 2820 30680 2832 30714
rect 2866 30680 2878 30714
rect 2820 30646 2878 30680
rect 2820 30612 2832 30646
rect 2866 30612 2878 30646
rect 2820 30578 2878 30612
rect 2820 30544 2832 30578
rect 2866 30544 2878 30578
rect 2820 30510 2878 30544
rect 2820 30476 2832 30510
rect 2866 30476 2878 30510
rect 2820 30442 2878 30476
rect 2820 30408 2832 30442
rect 2866 30408 2878 30442
rect 2820 30374 2878 30408
rect 2820 30340 2832 30374
rect 2866 30340 2878 30374
rect 2820 30306 2878 30340
rect 2820 30272 2832 30306
rect 2866 30272 2878 30306
rect 2820 30238 2878 30272
rect 2820 30204 2832 30238
rect 2866 30204 2878 30238
rect 2820 30170 2878 30204
rect 2820 30136 2832 30170
rect 2866 30136 2878 30170
rect 2820 30102 2878 30136
rect 2820 30068 2832 30102
rect 2866 30068 2878 30102
rect 2820 30034 2878 30068
rect 2820 30000 2832 30034
rect 2866 30000 2878 30034
rect 2820 29959 2878 30000
rect 2978 30918 3036 30959
rect 2978 30884 2990 30918
rect 3024 30884 3036 30918
rect 2978 30850 3036 30884
rect 2978 30816 2990 30850
rect 3024 30816 3036 30850
rect 2978 30782 3036 30816
rect 2978 30748 2990 30782
rect 3024 30748 3036 30782
rect 2978 30714 3036 30748
rect 2978 30680 2990 30714
rect 3024 30680 3036 30714
rect 2978 30646 3036 30680
rect 2978 30612 2990 30646
rect 3024 30612 3036 30646
rect 2978 30578 3036 30612
rect 2978 30544 2990 30578
rect 3024 30544 3036 30578
rect 2978 30510 3036 30544
rect 2978 30476 2990 30510
rect 3024 30476 3036 30510
rect 2978 30442 3036 30476
rect 2978 30408 2990 30442
rect 3024 30408 3036 30442
rect 2978 30374 3036 30408
rect 2978 30340 2990 30374
rect 3024 30340 3036 30374
rect 2978 30306 3036 30340
rect 2978 30272 2990 30306
rect 3024 30272 3036 30306
rect 2978 30238 3036 30272
rect 2978 30204 2990 30238
rect 3024 30204 3036 30238
rect 2978 30170 3036 30204
rect 2978 30136 2990 30170
rect 3024 30136 3036 30170
rect 2978 30102 3036 30136
rect 2978 30068 2990 30102
rect 3024 30068 3036 30102
rect 2978 30034 3036 30068
rect 2978 30000 2990 30034
rect 3024 30000 3036 30034
rect 2978 29959 3036 30000
rect 3136 30918 3194 30959
rect 3136 30884 3148 30918
rect 3182 30884 3194 30918
rect 3136 30850 3194 30884
rect 3136 30816 3148 30850
rect 3182 30816 3194 30850
rect 3136 30782 3194 30816
rect 3136 30748 3148 30782
rect 3182 30748 3194 30782
rect 3136 30714 3194 30748
rect 3136 30680 3148 30714
rect 3182 30680 3194 30714
rect 3136 30646 3194 30680
rect 3136 30612 3148 30646
rect 3182 30612 3194 30646
rect 3136 30578 3194 30612
rect 3136 30544 3148 30578
rect 3182 30544 3194 30578
rect 3136 30510 3194 30544
rect 3136 30476 3148 30510
rect 3182 30476 3194 30510
rect 3136 30442 3194 30476
rect 3136 30408 3148 30442
rect 3182 30408 3194 30442
rect 3136 30374 3194 30408
rect 3136 30340 3148 30374
rect 3182 30340 3194 30374
rect 3136 30306 3194 30340
rect 3136 30272 3148 30306
rect 3182 30272 3194 30306
rect 3136 30238 3194 30272
rect 3136 30204 3148 30238
rect 3182 30204 3194 30238
rect 3136 30170 3194 30204
rect 3136 30136 3148 30170
rect 3182 30136 3194 30170
rect 3136 30102 3194 30136
rect 3136 30068 3148 30102
rect 3182 30068 3194 30102
rect 3136 30034 3194 30068
rect 3136 30000 3148 30034
rect 3182 30000 3194 30034
rect 3136 29959 3194 30000
rect -1684 29248 -1626 29289
rect -1684 29214 -1672 29248
rect -1638 29214 -1626 29248
rect -1684 29180 -1626 29214
rect -1684 29146 -1672 29180
rect -1638 29146 -1626 29180
rect -1684 29112 -1626 29146
rect -1684 29078 -1672 29112
rect -1638 29078 -1626 29112
rect -1684 29044 -1626 29078
rect -1684 29010 -1672 29044
rect -1638 29010 -1626 29044
rect -1684 28976 -1626 29010
rect -1684 28942 -1672 28976
rect -1638 28942 -1626 28976
rect -1684 28908 -1626 28942
rect -1684 28874 -1672 28908
rect -1638 28874 -1626 28908
rect -1684 28840 -1626 28874
rect -1684 28806 -1672 28840
rect -1638 28806 -1626 28840
rect -1684 28772 -1626 28806
rect -1684 28738 -1672 28772
rect -1638 28738 -1626 28772
rect -1684 28704 -1626 28738
rect -1684 28670 -1672 28704
rect -1638 28670 -1626 28704
rect -1684 28636 -1626 28670
rect -1684 28602 -1672 28636
rect -1638 28602 -1626 28636
rect -1684 28568 -1626 28602
rect -1684 28534 -1672 28568
rect -1638 28534 -1626 28568
rect -1684 28500 -1626 28534
rect -1684 28466 -1672 28500
rect -1638 28466 -1626 28500
rect -1684 28432 -1626 28466
rect -1684 28398 -1672 28432
rect -1638 28398 -1626 28432
rect -1684 28364 -1626 28398
rect -1684 28330 -1672 28364
rect -1638 28330 -1626 28364
rect -1684 28289 -1626 28330
rect -1526 29248 -1468 29289
rect -1526 29214 -1514 29248
rect -1480 29214 -1468 29248
rect -1526 29180 -1468 29214
rect -1526 29146 -1514 29180
rect -1480 29146 -1468 29180
rect -1526 29112 -1468 29146
rect -1526 29078 -1514 29112
rect -1480 29078 -1468 29112
rect -1526 29044 -1468 29078
rect -1526 29010 -1514 29044
rect -1480 29010 -1468 29044
rect -1526 28976 -1468 29010
rect -1526 28942 -1514 28976
rect -1480 28942 -1468 28976
rect -1526 28908 -1468 28942
rect -1526 28874 -1514 28908
rect -1480 28874 -1468 28908
rect -1526 28840 -1468 28874
rect -1526 28806 -1514 28840
rect -1480 28806 -1468 28840
rect -1526 28772 -1468 28806
rect -1526 28738 -1514 28772
rect -1480 28738 -1468 28772
rect -1526 28704 -1468 28738
rect -1526 28670 -1514 28704
rect -1480 28670 -1468 28704
rect -1526 28636 -1468 28670
rect -1526 28602 -1514 28636
rect -1480 28602 -1468 28636
rect -1526 28568 -1468 28602
rect -1526 28534 -1514 28568
rect -1480 28534 -1468 28568
rect -1526 28500 -1468 28534
rect -1526 28466 -1514 28500
rect -1480 28466 -1468 28500
rect -1526 28432 -1468 28466
rect -1526 28398 -1514 28432
rect -1480 28398 -1468 28432
rect -1526 28364 -1468 28398
rect -1526 28330 -1514 28364
rect -1480 28330 -1468 28364
rect -1526 28289 -1468 28330
rect -1368 29248 -1310 29289
rect -1368 29214 -1356 29248
rect -1322 29214 -1310 29248
rect -1368 29180 -1310 29214
rect -1368 29146 -1356 29180
rect -1322 29146 -1310 29180
rect -1368 29112 -1310 29146
rect -1368 29078 -1356 29112
rect -1322 29078 -1310 29112
rect -1368 29044 -1310 29078
rect -1368 29010 -1356 29044
rect -1322 29010 -1310 29044
rect -1368 28976 -1310 29010
rect -1368 28942 -1356 28976
rect -1322 28942 -1310 28976
rect -1368 28908 -1310 28942
rect -1368 28874 -1356 28908
rect -1322 28874 -1310 28908
rect -1368 28840 -1310 28874
rect -1368 28806 -1356 28840
rect -1322 28806 -1310 28840
rect -1368 28772 -1310 28806
rect -1368 28738 -1356 28772
rect -1322 28738 -1310 28772
rect -1368 28704 -1310 28738
rect -1368 28670 -1356 28704
rect -1322 28670 -1310 28704
rect -1368 28636 -1310 28670
rect -1368 28602 -1356 28636
rect -1322 28602 -1310 28636
rect -1368 28568 -1310 28602
rect -1368 28534 -1356 28568
rect -1322 28534 -1310 28568
rect -1368 28500 -1310 28534
rect -1368 28466 -1356 28500
rect -1322 28466 -1310 28500
rect -1368 28432 -1310 28466
rect -1368 28398 -1356 28432
rect -1322 28398 -1310 28432
rect -1368 28364 -1310 28398
rect -1368 28330 -1356 28364
rect -1322 28330 -1310 28364
rect -1368 28289 -1310 28330
rect -1210 29248 -1152 29289
rect -1210 29214 -1198 29248
rect -1164 29214 -1152 29248
rect -1210 29180 -1152 29214
rect -1210 29146 -1198 29180
rect -1164 29146 -1152 29180
rect -1210 29112 -1152 29146
rect -1210 29078 -1198 29112
rect -1164 29078 -1152 29112
rect -1210 29044 -1152 29078
rect -1210 29010 -1198 29044
rect -1164 29010 -1152 29044
rect -1210 28976 -1152 29010
rect -1210 28942 -1198 28976
rect -1164 28942 -1152 28976
rect -1210 28908 -1152 28942
rect -1210 28874 -1198 28908
rect -1164 28874 -1152 28908
rect -1210 28840 -1152 28874
rect -1210 28806 -1198 28840
rect -1164 28806 -1152 28840
rect -1210 28772 -1152 28806
rect -1210 28738 -1198 28772
rect -1164 28738 -1152 28772
rect -1210 28704 -1152 28738
rect -1210 28670 -1198 28704
rect -1164 28670 -1152 28704
rect -1210 28636 -1152 28670
rect -1210 28602 -1198 28636
rect -1164 28602 -1152 28636
rect -1210 28568 -1152 28602
rect -1210 28534 -1198 28568
rect -1164 28534 -1152 28568
rect -1210 28500 -1152 28534
rect -1210 28466 -1198 28500
rect -1164 28466 -1152 28500
rect -1210 28432 -1152 28466
rect -1210 28398 -1198 28432
rect -1164 28398 -1152 28432
rect -1210 28364 -1152 28398
rect -1210 28330 -1198 28364
rect -1164 28330 -1152 28364
rect -1210 28289 -1152 28330
rect -1052 29248 -994 29289
rect -1052 29214 -1040 29248
rect -1006 29214 -994 29248
rect -1052 29180 -994 29214
rect -1052 29146 -1040 29180
rect -1006 29146 -994 29180
rect -1052 29112 -994 29146
rect -1052 29078 -1040 29112
rect -1006 29078 -994 29112
rect -1052 29044 -994 29078
rect -1052 29010 -1040 29044
rect -1006 29010 -994 29044
rect -1052 28976 -994 29010
rect -1052 28942 -1040 28976
rect -1006 28942 -994 28976
rect -1052 28908 -994 28942
rect -1052 28874 -1040 28908
rect -1006 28874 -994 28908
rect -1052 28840 -994 28874
rect -1052 28806 -1040 28840
rect -1006 28806 -994 28840
rect -1052 28772 -994 28806
rect -1052 28738 -1040 28772
rect -1006 28738 -994 28772
rect -1052 28704 -994 28738
rect -1052 28670 -1040 28704
rect -1006 28670 -994 28704
rect -1052 28636 -994 28670
rect -1052 28602 -1040 28636
rect -1006 28602 -994 28636
rect -1052 28568 -994 28602
rect -1052 28534 -1040 28568
rect -1006 28534 -994 28568
rect -1052 28500 -994 28534
rect -1052 28466 -1040 28500
rect -1006 28466 -994 28500
rect -1052 28432 -994 28466
rect -1052 28398 -1040 28432
rect -1006 28398 -994 28432
rect -1052 28364 -994 28398
rect -1052 28330 -1040 28364
rect -1006 28330 -994 28364
rect -1052 28289 -994 28330
rect -894 29248 -836 29289
rect -894 29214 -882 29248
rect -848 29214 -836 29248
rect -894 29180 -836 29214
rect -894 29146 -882 29180
rect -848 29146 -836 29180
rect -894 29112 -836 29146
rect -894 29078 -882 29112
rect -848 29078 -836 29112
rect -894 29044 -836 29078
rect -894 29010 -882 29044
rect -848 29010 -836 29044
rect -894 28976 -836 29010
rect -894 28942 -882 28976
rect -848 28942 -836 28976
rect -894 28908 -836 28942
rect -894 28874 -882 28908
rect -848 28874 -836 28908
rect -894 28840 -836 28874
rect -894 28806 -882 28840
rect -848 28806 -836 28840
rect -894 28772 -836 28806
rect -894 28738 -882 28772
rect -848 28738 -836 28772
rect -894 28704 -836 28738
rect -894 28670 -882 28704
rect -848 28670 -836 28704
rect -894 28636 -836 28670
rect -894 28602 -882 28636
rect -848 28602 -836 28636
rect -894 28568 -836 28602
rect -894 28534 -882 28568
rect -848 28534 -836 28568
rect -894 28500 -836 28534
rect -894 28466 -882 28500
rect -848 28466 -836 28500
rect -894 28432 -836 28466
rect -894 28398 -882 28432
rect -848 28398 -836 28432
rect -894 28364 -836 28398
rect -894 28330 -882 28364
rect -848 28330 -836 28364
rect -894 28289 -836 28330
rect -736 29248 -678 29289
rect -736 29214 -724 29248
rect -690 29214 -678 29248
rect -736 29180 -678 29214
rect -736 29146 -724 29180
rect -690 29146 -678 29180
rect -736 29112 -678 29146
rect -736 29078 -724 29112
rect -690 29078 -678 29112
rect -736 29044 -678 29078
rect -736 29010 -724 29044
rect -690 29010 -678 29044
rect -736 28976 -678 29010
rect -736 28942 -724 28976
rect -690 28942 -678 28976
rect -736 28908 -678 28942
rect -736 28874 -724 28908
rect -690 28874 -678 28908
rect -736 28840 -678 28874
rect -736 28806 -724 28840
rect -690 28806 -678 28840
rect -736 28772 -678 28806
rect -736 28738 -724 28772
rect -690 28738 -678 28772
rect -736 28704 -678 28738
rect -736 28670 -724 28704
rect -690 28670 -678 28704
rect -736 28636 -678 28670
rect -736 28602 -724 28636
rect -690 28602 -678 28636
rect -736 28568 -678 28602
rect -736 28534 -724 28568
rect -690 28534 -678 28568
rect -736 28500 -678 28534
rect -736 28466 -724 28500
rect -690 28466 -678 28500
rect -736 28432 -678 28466
rect -736 28398 -724 28432
rect -690 28398 -678 28432
rect -736 28364 -678 28398
rect -736 28330 -724 28364
rect -690 28330 -678 28364
rect -736 28289 -678 28330
rect -578 29248 -520 29289
rect -578 29214 -566 29248
rect -532 29214 -520 29248
rect -578 29180 -520 29214
rect -578 29146 -566 29180
rect -532 29146 -520 29180
rect -578 29112 -520 29146
rect -578 29078 -566 29112
rect -532 29078 -520 29112
rect -578 29044 -520 29078
rect -578 29010 -566 29044
rect -532 29010 -520 29044
rect -578 28976 -520 29010
rect -578 28942 -566 28976
rect -532 28942 -520 28976
rect -578 28908 -520 28942
rect -578 28874 -566 28908
rect -532 28874 -520 28908
rect -578 28840 -520 28874
rect -578 28806 -566 28840
rect -532 28806 -520 28840
rect -578 28772 -520 28806
rect -578 28738 -566 28772
rect -532 28738 -520 28772
rect -578 28704 -520 28738
rect -578 28670 -566 28704
rect -532 28670 -520 28704
rect -578 28636 -520 28670
rect -578 28602 -566 28636
rect -532 28602 -520 28636
rect -578 28568 -520 28602
rect -578 28534 -566 28568
rect -532 28534 -520 28568
rect -578 28500 -520 28534
rect -578 28466 -566 28500
rect -532 28466 -520 28500
rect -578 28432 -520 28466
rect -578 28398 -566 28432
rect -532 28398 -520 28432
rect -578 28364 -520 28398
rect -578 28330 -566 28364
rect -532 28330 -520 28364
rect -578 28289 -520 28330
rect -420 29248 -362 29289
rect -420 29214 -408 29248
rect -374 29214 -362 29248
rect -420 29180 -362 29214
rect -420 29146 -408 29180
rect -374 29146 -362 29180
rect -420 29112 -362 29146
rect -420 29078 -408 29112
rect -374 29078 -362 29112
rect -420 29044 -362 29078
rect -420 29010 -408 29044
rect -374 29010 -362 29044
rect -420 28976 -362 29010
rect -420 28942 -408 28976
rect -374 28942 -362 28976
rect -420 28908 -362 28942
rect -420 28874 -408 28908
rect -374 28874 -362 28908
rect -420 28840 -362 28874
rect -420 28806 -408 28840
rect -374 28806 -362 28840
rect -420 28772 -362 28806
rect -420 28738 -408 28772
rect -374 28738 -362 28772
rect -420 28704 -362 28738
rect -420 28670 -408 28704
rect -374 28670 -362 28704
rect -420 28636 -362 28670
rect -420 28602 -408 28636
rect -374 28602 -362 28636
rect -420 28568 -362 28602
rect -420 28534 -408 28568
rect -374 28534 -362 28568
rect -420 28500 -362 28534
rect -420 28466 -408 28500
rect -374 28466 -362 28500
rect -420 28432 -362 28466
rect -420 28398 -408 28432
rect -374 28398 -362 28432
rect -420 28364 -362 28398
rect -420 28330 -408 28364
rect -374 28330 -362 28364
rect -420 28289 -362 28330
rect -262 29248 -204 29289
rect -262 29214 -250 29248
rect -216 29214 -204 29248
rect -262 29180 -204 29214
rect -262 29146 -250 29180
rect -216 29146 -204 29180
rect -262 29112 -204 29146
rect -262 29078 -250 29112
rect -216 29078 -204 29112
rect -262 29044 -204 29078
rect -262 29010 -250 29044
rect -216 29010 -204 29044
rect -262 28976 -204 29010
rect -262 28942 -250 28976
rect -216 28942 -204 28976
rect -262 28908 -204 28942
rect -262 28874 -250 28908
rect -216 28874 -204 28908
rect -262 28840 -204 28874
rect -262 28806 -250 28840
rect -216 28806 -204 28840
rect -262 28772 -204 28806
rect -262 28738 -250 28772
rect -216 28738 -204 28772
rect -262 28704 -204 28738
rect -262 28670 -250 28704
rect -216 28670 -204 28704
rect -262 28636 -204 28670
rect -262 28602 -250 28636
rect -216 28602 -204 28636
rect -262 28568 -204 28602
rect -262 28534 -250 28568
rect -216 28534 -204 28568
rect -262 28500 -204 28534
rect -262 28466 -250 28500
rect -216 28466 -204 28500
rect -262 28432 -204 28466
rect -262 28398 -250 28432
rect -216 28398 -204 28432
rect -262 28364 -204 28398
rect -262 28330 -250 28364
rect -216 28330 -204 28364
rect -262 28289 -204 28330
rect -104 29248 -46 29289
rect -104 29214 -92 29248
rect -58 29214 -46 29248
rect -104 29180 -46 29214
rect -104 29146 -92 29180
rect -58 29146 -46 29180
rect -104 29112 -46 29146
rect -104 29078 -92 29112
rect -58 29078 -46 29112
rect -104 29044 -46 29078
rect -104 29010 -92 29044
rect -58 29010 -46 29044
rect -104 28976 -46 29010
rect -104 28942 -92 28976
rect -58 28942 -46 28976
rect -104 28908 -46 28942
rect -104 28874 -92 28908
rect -58 28874 -46 28908
rect -104 28840 -46 28874
rect -104 28806 -92 28840
rect -58 28806 -46 28840
rect -104 28772 -46 28806
rect -104 28738 -92 28772
rect -58 28738 -46 28772
rect -104 28704 -46 28738
rect -104 28670 -92 28704
rect -58 28670 -46 28704
rect -104 28636 -46 28670
rect -104 28602 -92 28636
rect -58 28602 -46 28636
rect -104 28568 -46 28602
rect -104 28534 -92 28568
rect -58 28534 -46 28568
rect -104 28500 -46 28534
rect -104 28466 -92 28500
rect -58 28466 -46 28500
rect -104 28432 -46 28466
rect -104 28398 -92 28432
rect -58 28398 -46 28432
rect -104 28364 -46 28398
rect -104 28330 -92 28364
rect -58 28330 -46 28364
rect -104 28289 -46 28330
rect 54 29248 112 29289
rect 54 29214 66 29248
rect 100 29214 112 29248
rect 54 29180 112 29214
rect 54 29146 66 29180
rect 100 29146 112 29180
rect 54 29112 112 29146
rect 54 29078 66 29112
rect 100 29078 112 29112
rect 54 29044 112 29078
rect 54 29010 66 29044
rect 100 29010 112 29044
rect 54 28976 112 29010
rect 54 28942 66 28976
rect 100 28942 112 28976
rect 54 28908 112 28942
rect 54 28874 66 28908
rect 100 28874 112 28908
rect 54 28840 112 28874
rect 54 28806 66 28840
rect 100 28806 112 28840
rect 54 28772 112 28806
rect 54 28738 66 28772
rect 100 28738 112 28772
rect 54 28704 112 28738
rect 54 28670 66 28704
rect 100 28670 112 28704
rect 54 28636 112 28670
rect 54 28602 66 28636
rect 100 28602 112 28636
rect 54 28568 112 28602
rect 54 28534 66 28568
rect 100 28534 112 28568
rect 54 28500 112 28534
rect 54 28466 66 28500
rect 100 28466 112 28500
rect 54 28432 112 28466
rect 54 28398 66 28432
rect 100 28398 112 28432
rect 54 28364 112 28398
rect 54 28330 66 28364
rect 100 28330 112 28364
rect 54 28289 112 28330
rect 212 29248 270 29289
rect 212 29214 224 29248
rect 258 29214 270 29248
rect 212 29180 270 29214
rect 212 29146 224 29180
rect 258 29146 270 29180
rect 212 29112 270 29146
rect 212 29078 224 29112
rect 258 29078 270 29112
rect 212 29044 270 29078
rect 212 29010 224 29044
rect 258 29010 270 29044
rect 212 28976 270 29010
rect 212 28942 224 28976
rect 258 28942 270 28976
rect 212 28908 270 28942
rect 212 28874 224 28908
rect 258 28874 270 28908
rect 212 28840 270 28874
rect 212 28806 224 28840
rect 258 28806 270 28840
rect 212 28772 270 28806
rect 212 28738 224 28772
rect 258 28738 270 28772
rect 212 28704 270 28738
rect 212 28670 224 28704
rect 258 28670 270 28704
rect 212 28636 270 28670
rect 212 28602 224 28636
rect 258 28602 270 28636
rect 212 28568 270 28602
rect 212 28534 224 28568
rect 258 28534 270 28568
rect 212 28500 270 28534
rect 212 28466 224 28500
rect 258 28466 270 28500
rect 212 28432 270 28466
rect 212 28398 224 28432
rect 258 28398 270 28432
rect 212 28364 270 28398
rect 212 28330 224 28364
rect 258 28330 270 28364
rect 212 28289 270 28330
rect 370 29248 428 29289
rect 370 29214 382 29248
rect 416 29214 428 29248
rect 370 29180 428 29214
rect 370 29146 382 29180
rect 416 29146 428 29180
rect 370 29112 428 29146
rect 370 29078 382 29112
rect 416 29078 428 29112
rect 370 29044 428 29078
rect 370 29010 382 29044
rect 416 29010 428 29044
rect 370 28976 428 29010
rect 370 28942 382 28976
rect 416 28942 428 28976
rect 370 28908 428 28942
rect 370 28874 382 28908
rect 416 28874 428 28908
rect 370 28840 428 28874
rect 370 28806 382 28840
rect 416 28806 428 28840
rect 370 28772 428 28806
rect 370 28738 382 28772
rect 416 28738 428 28772
rect 370 28704 428 28738
rect 370 28670 382 28704
rect 416 28670 428 28704
rect 370 28636 428 28670
rect 370 28602 382 28636
rect 416 28602 428 28636
rect 370 28568 428 28602
rect 370 28534 382 28568
rect 416 28534 428 28568
rect 370 28500 428 28534
rect 370 28466 382 28500
rect 416 28466 428 28500
rect 370 28432 428 28466
rect 370 28398 382 28432
rect 416 28398 428 28432
rect 370 28364 428 28398
rect 370 28330 382 28364
rect 416 28330 428 28364
rect 370 28289 428 28330
rect 528 29248 586 29289
rect 528 29214 540 29248
rect 574 29214 586 29248
rect 528 29180 586 29214
rect 528 29146 540 29180
rect 574 29146 586 29180
rect 528 29112 586 29146
rect 528 29078 540 29112
rect 574 29078 586 29112
rect 528 29044 586 29078
rect 528 29010 540 29044
rect 574 29010 586 29044
rect 528 28976 586 29010
rect 528 28942 540 28976
rect 574 28942 586 28976
rect 528 28908 586 28942
rect 528 28874 540 28908
rect 574 28874 586 28908
rect 528 28840 586 28874
rect 528 28806 540 28840
rect 574 28806 586 28840
rect 528 28772 586 28806
rect 528 28738 540 28772
rect 574 28738 586 28772
rect 528 28704 586 28738
rect 528 28670 540 28704
rect 574 28670 586 28704
rect 528 28636 586 28670
rect 528 28602 540 28636
rect 574 28602 586 28636
rect 528 28568 586 28602
rect 528 28534 540 28568
rect 574 28534 586 28568
rect 528 28500 586 28534
rect 528 28466 540 28500
rect 574 28466 586 28500
rect 528 28432 586 28466
rect 528 28398 540 28432
rect 574 28398 586 28432
rect 528 28364 586 28398
rect 528 28330 540 28364
rect 574 28330 586 28364
rect 528 28289 586 28330
rect 686 29248 744 29289
rect 686 29214 698 29248
rect 732 29214 744 29248
rect 686 29180 744 29214
rect 686 29146 698 29180
rect 732 29146 744 29180
rect 686 29112 744 29146
rect 686 29078 698 29112
rect 732 29078 744 29112
rect 686 29044 744 29078
rect 686 29010 698 29044
rect 732 29010 744 29044
rect 686 28976 744 29010
rect 686 28942 698 28976
rect 732 28942 744 28976
rect 686 28908 744 28942
rect 686 28874 698 28908
rect 732 28874 744 28908
rect 686 28840 744 28874
rect 686 28806 698 28840
rect 732 28806 744 28840
rect 686 28772 744 28806
rect 686 28738 698 28772
rect 732 28738 744 28772
rect 686 28704 744 28738
rect 686 28670 698 28704
rect 732 28670 744 28704
rect 686 28636 744 28670
rect 686 28602 698 28636
rect 732 28602 744 28636
rect 686 28568 744 28602
rect 686 28534 698 28568
rect 732 28534 744 28568
rect 686 28500 744 28534
rect 686 28466 698 28500
rect 732 28466 744 28500
rect 686 28432 744 28466
rect 686 28398 698 28432
rect 732 28398 744 28432
rect 686 28364 744 28398
rect 686 28330 698 28364
rect 732 28330 744 28364
rect 686 28289 744 28330
rect 844 29248 902 29289
rect 844 29214 856 29248
rect 890 29214 902 29248
rect 844 29180 902 29214
rect 844 29146 856 29180
rect 890 29146 902 29180
rect 844 29112 902 29146
rect 844 29078 856 29112
rect 890 29078 902 29112
rect 844 29044 902 29078
rect 844 29010 856 29044
rect 890 29010 902 29044
rect 844 28976 902 29010
rect 844 28942 856 28976
rect 890 28942 902 28976
rect 844 28908 902 28942
rect 844 28874 856 28908
rect 890 28874 902 28908
rect 844 28840 902 28874
rect 844 28806 856 28840
rect 890 28806 902 28840
rect 844 28772 902 28806
rect 844 28738 856 28772
rect 890 28738 902 28772
rect 844 28704 902 28738
rect 844 28670 856 28704
rect 890 28670 902 28704
rect 844 28636 902 28670
rect 844 28602 856 28636
rect 890 28602 902 28636
rect 844 28568 902 28602
rect 844 28534 856 28568
rect 890 28534 902 28568
rect 844 28500 902 28534
rect 844 28466 856 28500
rect 890 28466 902 28500
rect 844 28432 902 28466
rect 844 28398 856 28432
rect 890 28398 902 28432
rect 844 28364 902 28398
rect 844 28330 856 28364
rect 890 28330 902 28364
rect 844 28289 902 28330
rect 1002 29248 1060 29289
rect 1002 29214 1014 29248
rect 1048 29214 1060 29248
rect 1002 29180 1060 29214
rect 1002 29146 1014 29180
rect 1048 29146 1060 29180
rect 1002 29112 1060 29146
rect 1002 29078 1014 29112
rect 1048 29078 1060 29112
rect 1002 29044 1060 29078
rect 1002 29010 1014 29044
rect 1048 29010 1060 29044
rect 1002 28976 1060 29010
rect 1002 28942 1014 28976
rect 1048 28942 1060 28976
rect 1002 28908 1060 28942
rect 1002 28874 1014 28908
rect 1048 28874 1060 28908
rect 1002 28840 1060 28874
rect 1002 28806 1014 28840
rect 1048 28806 1060 28840
rect 1002 28772 1060 28806
rect 1002 28738 1014 28772
rect 1048 28738 1060 28772
rect 1002 28704 1060 28738
rect 1002 28670 1014 28704
rect 1048 28670 1060 28704
rect 1002 28636 1060 28670
rect 1002 28602 1014 28636
rect 1048 28602 1060 28636
rect 1002 28568 1060 28602
rect 1002 28534 1014 28568
rect 1048 28534 1060 28568
rect 1002 28500 1060 28534
rect 1002 28466 1014 28500
rect 1048 28466 1060 28500
rect 1002 28432 1060 28466
rect 1002 28398 1014 28432
rect 1048 28398 1060 28432
rect 1002 28364 1060 28398
rect 1002 28330 1014 28364
rect 1048 28330 1060 28364
rect 1002 28289 1060 28330
rect 1160 29248 1218 29289
rect 1160 29214 1172 29248
rect 1206 29214 1218 29248
rect 1160 29180 1218 29214
rect 1160 29146 1172 29180
rect 1206 29146 1218 29180
rect 1160 29112 1218 29146
rect 1160 29078 1172 29112
rect 1206 29078 1218 29112
rect 1160 29044 1218 29078
rect 1160 29010 1172 29044
rect 1206 29010 1218 29044
rect 1160 28976 1218 29010
rect 1160 28942 1172 28976
rect 1206 28942 1218 28976
rect 1160 28908 1218 28942
rect 1160 28874 1172 28908
rect 1206 28874 1218 28908
rect 1160 28840 1218 28874
rect 1160 28806 1172 28840
rect 1206 28806 1218 28840
rect 1160 28772 1218 28806
rect 1160 28738 1172 28772
rect 1206 28738 1218 28772
rect 1160 28704 1218 28738
rect 1160 28670 1172 28704
rect 1206 28670 1218 28704
rect 1160 28636 1218 28670
rect 1160 28602 1172 28636
rect 1206 28602 1218 28636
rect 1160 28568 1218 28602
rect 1160 28534 1172 28568
rect 1206 28534 1218 28568
rect 1160 28500 1218 28534
rect 1160 28466 1172 28500
rect 1206 28466 1218 28500
rect 1160 28432 1218 28466
rect 1160 28398 1172 28432
rect 1206 28398 1218 28432
rect 1160 28364 1218 28398
rect 1160 28330 1172 28364
rect 1206 28330 1218 28364
rect 1160 28289 1218 28330
rect 1318 29248 1376 29289
rect 1318 29214 1330 29248
rect 1364 29214 1376 29248
rect 1318 29180 1376 29214
rect 1318 29146 1330 29180
rect 1364 29146 1376 29180
rect 1318 29112 1376 29146
rect 1318 29078 1330 29112
rect 1364 29078 1376 29112
rect 1318 29044 1376 29078
rect 1318 29010 1330 29044
rect 1364 29010 1376 29044
rect 1318 28976 1376 29010
rect 1318 28942 1330 28976
rect 1364 28942 1376 28976
rect 1318 28908 1376 28942
rect 1318 28874 1330 28908
rect 1364 28874 1376 28908
rect 1318 28840 1376 28874
rect 1318 28806 1330 28840
rect 1364 28806 1376 28840
rect 1318 28772 1376 28806
rect 1318 28738 1330 28772
rect 1364 28738 1376 28772
rect 1318 28704 1376 28738
rect 1318 28670 1330 28704
rect 1364 28670 1376 28704
rect 1318 28636 1376 28670
rect 1318 28602 1330 28636
rect 1364 28602 1376 28636
rect 1318 28568 1376 28602
rect 1318 28534 1330 28568
rect 1364 28534 1376 28568
rect 1318 28500 1376 28534
rect 1318 28466 1330 28500
rect 1364 28466 1376 28500
rect 1318 28432 1376 28466
rect 1318 28398 1330 28432
rect 1364 28398 1376 28432
rect 1318 28364 1376 28398
rect 1318 28330 1330 28364
rect 1364 28330 1376 28364
rect 1318 28289 1376 28330
rect 1476 29248 1534 29289
rect 1476 29214 1488 29248
rect 1522 29214 1534 29248
rect 1476 29180 1534 29214
rect 1476 29146 1488 29180
rect 1522 29146 1534 29180
rect 1476 29112 1534 29146
rect 1476 29078 1488 29112
rect 1522 29078 1534 29112
rect 1476 29044 1534 29078
rect 1476 29010 1488 29044
rect 1522 29010 1534 29044
rect 1476 28976 1534 29010
rect 1476 28942 1488 28976
rect 1522 28942 1534 28976
rect 1476 28908 1534 28942
rect 1476 28874 1488 28908
rect 1522 28874 1534 28908
rect 1476 28840 1534 28874
rect 1476 28806 1488 28840
rect 1522 28806 1534 28840
rect 1476 28772 1534 28806
rect 1476 28738 1488 28772
rect 1522 28738 1534 28772
rect 1476 28704 1534 28738
rect 1476 28670 1488 28704
rect 1522 28670 1534 28704
rect 1476 28636 1534 28670
rect 1476 28602 1488 28636
rect 1522 28602 1534 28636
rect 1476 28568 1534 28602
rect 1476 28534 1488 28568
rect 1522 28534 1534 28568
rect 1476 28500 1534 28534
rect 1476 28466 1488 28500
rect 1522 28466 1534 28500
rect 1476 28432 1534 28466
rect 1476 28398 1488 28432
rect 1522 28398 1534 28432
rect 1476 28364 1534 28398
rect 1476 28330 1488 28364
rect 1522 28330 1534 28364
rect 1476 28289 1534 28330
rect 1634 29248 1692 29289
rect 1634 29214 1646 29248
rect 1680 29214 1692 29248
rect 1634 29180 1692 29214
rect 1634 29146 1646 29180
rect 1680 29146 1692 29180
rect 1634 29112 1692 29146
rect 1634 29078 1646 29112
rect 1680 29078 1692 29112
rect 1634 29044 1692 29078
rect 1634 29010 1646 29044
rect 1680 29010 1692 29044
rect 1634 28976 1692 29010
rect 1634 28942 1646 28976
rect 1680 28942 1692 28976
rect 1634 28908 1692 28942
rect 1634 28874 1646 28908
rect 1680 28874 1692 28908
rect 1634 28840 1692 28874
rect 1634 28806 1646 28840
rect 1680 28806 1692 28840
rect 1634 28772 1692 28806
rect 1634 28738 1646 28772
rect 1680 28738 1692 28772
rect 1634 28704 1692 28738
rect 1634 28670 1646 28704
rect 1680 28670 1692 28704
rect 1634 28636 1692 28670
rect 1634 28602 1646 28636
rect 1680 28602 1692 28636
rect 1634 28568 1692 28602
rect 1634 28534 1646 28568
rect 1680 28534 1692 28568
rect 1634 28500 1692 28534
rect 1634 28466 1646 28500
rect 1680 28466 1692 28500
rect 1634 28432 1692 28466
rect 1634 28398 1646 28432
rect 1680 28398 1692 28432
rect 1634 28364 1692 28398
rect 1634 28330 1646 28364
rect 1680 28330 1692 28364
rect 1634 28289 1692 28330
rect -1684 27708 -1626 27749
rect -1684 27674 -1672 27708
rect -1638 27674 -1626 27708
rect -1684 27640 -1626 27674
rect -1684 27606 -1672 27640
rect -1638 27606 -1626 27640
rect -1684 27572 -1626 27606
rect -1684 27538 -1672 27572
rect -1638 27538 -1626 27572
rect -1684 27504 -1626 27538
rect -1684 27470 -1672 27504
rect -1638 27470 -1626 27504
rect -1684 27436 -1626 27470
rect -1684 27402 -1672 27436
rect -1638 27402 -1626 27436
rect -1684 27368 -1626 27402
rect -1684 27334 -1672 27368
rect -1638 27334 -1626 27368
rect -1684 27300 -1626 27334
rect -1684 27266 -1672 27300
rect -1638 27266 -1626 27300
rect -1684 27232 -1626 27266
rect -1684 27198 -1672 27232
rect -1638 27198 -1626 27232
rect -1684 27164 -1626 27198
rect -1684 27130 -1672 27164
rect -1638 27130 -1626 27164
rect -1684 27096 -1626 27130
rect -1684 27062 -1672 27096
rect -1638 27062 -1626 27096
rect -1684 27028 -1626 27062
rect -1684 26994 -1672 27028
rect -1638 26994 -1626 27028
rect -1684 26960 -1626 26994
rect -1684 26926 -1672 26960
rect -1638 26926 -1626 26960
rect -1684 26892 -1626 26926
rect -1684 26858 -1672 26892
rect -1638 26858 -1626 26892
rect -1684 26824 -1626 26858
rect -1684 26790 -1672 26824
rect -1638 26790 -1626 26824
rect -1684 26749 -1626 26790
rect -1526 27708 -1468 27749
rect -1526 27674 -1514 27708
rect -1480 27674 -1468 27708
rect -1526 27640 -1468 27674
rect -1526 27606 -1514 27640
rect -1480 27606 -1468 27640
rect -1526 27572 -1468 27606
rect -1526 27538 -1514 27572
rect -1480 27538 -1468 27572
rect -1526 27504 -1468 27538
rect -1526 27470 -1514 27504
rect -1480 27470 -1468 27504
rect -1526 27436 -1468 27470
rect -1526 27402 -1514 27436
rect -1480 27402 -1468 27436
rect -1526 27368 -1468 27402
rect -1526 27334 -1514 27368
rect -1480 27334 -1468 27368
rect -1526 27300 -1468 27334
rect -1526 27266 -1514 27300
rect -1480 27266 -1468 27300
rect -1526 27232 -1468 27266
rect -1526 27198 -1514 27232
rect -1480 27198 -1468 27232
rect -1526 27164 -1468 27198
rect -1526 27130 -1514 27164
rect -1480 27130 -1468 27164
rect -1526 27096 -1468 27130
rect -1526 27062 -1514 27096
rect -1480 27062 -1468 27096
rect -1526 27028 -1468 27062
rect -1526 26994 -1514 27028
rect -1480 26994 -1468 27028
rect -1526 26960 -1468 26994
rect -1526 26926 -1514 26960
rect -1480 26926 -1468 26960
rect -1526 26892 -1468 26926
rect -1526 26858 -1514 26892
rect -1480 26858 -1468 26892
rect -1526 26824 -1468 26858
rect -1526 26790 -1514 26824
rect -1480 26790 -1468 26824
rect -1526 26749 -1468 26790
rect -1368 27708 -1310 27749
rect -1368 27674 -1356 27708
rect -1322 27674 -1310 27708
rect -1368 27640 -1310 27674
rect -1368 27606 -1356 27640
rect -1322 27606 -1310 27640
rect -1368 27572 -1310 27606
rect -1368 27538 -1356 27572
rect -1322 27538 -1310 27572
rect -1368 27504 -1310 27538
rect -1368 27470 -1356 27504
rect -1322 27470 -1310 27504
rect -1368 27436 -1310 27470
rect -1368 27402 -1356 27436
rect -1322 27402 -1310 27436
rect -1368 27368 -1310 27402
rect -1368 27334 -1356 27368
rect -1322 27334 -1310 27368
rect -1368 27300 -1310 27334
rect -1368 27266 -1356 27300
rect -1322 27266 -1310 27300
rect -1368 27232 -1310 27266
rect -1368 27198 -1356 27232
rect -1322 27198 -1310 27232
rect -1368 27164 -1310 27198
rect -1368 27130 -1356 27164
rect -1322 27130 -1310 27164
rect -1368 27096 -1310 27130
rect -1368 27062 -1356 27096
rect -1322 27062 -1310 27096
rect -1368 27028 -1310 27062
rect -1368 26994 -1356 27028
rect -1322 26994 -1310 27028
rect -1368 26960 -1310 26994
rect -1368 26926 -1356 26960
rect -1322 26926 -1310 26960
rect -1368 26892 -1310 26926
rect -1368 26858 -1356 26892
rect -1322 26858 -1310 26892
rect -1368 26824 -1310 26858
rect -1368 26790 -1356 26824
rect -1322 26790 -1310 26824
rect -1368 26749 -1310 26790
rect -1210 27708 -1152 27749
rect -1210 27674 -1198 27708
rect -1164 27674 -1152 27708
rect -1210 27640 -1152 27674
rect -1210 27606 -1198 27640
rect -1164 27606 -1152 27640
rect -1210 27572 -1152 27606
rect -1210 27538 -1198 27572
rect -1164 27538 -1152 27572
rect -1210 27504 -1152 27538
rect -1210 27470 -1198 27504
rect -1164 27470 -1152 27504
rect -1210 27436 -1152 27470
rect -1210 27402 -1198 27436
rect -1164 27402 -1152 27436
rect -1210 27368 -1152 27402
rect -1210 27334 -1198 27368
rect -1164 27334 -1152 27368
rect -1210 27300 -1152 27334
rect -1210 27266 -1198 27300
rect -1164 27266 -1152 27300
rect -1210 27232 -1152 27266
rect -1210 27198 -1198 27232
rect -1164 27198 -1152 27232
rect -1210 27164 -1152 27198
rect -1210 27130 -1198 27164
rect -1164 27130 -1152 27164
rect -1210 27096 -1152 27130
rect -1210 27062 -1198 27096
rect -1164 27062 -1152 27096
rect -1210 27028 -1152 27062
rect -1210 26994 -1198 27028
rect -1164 26994 -1152 27028
rect -1210 26960 -1152 26994
rect -1210 26926 -1198 26960
rect -1164 26926 -1152 26960
rect -1210 26892 -1152 26926
rect -1210 26858 -1198 26892
rect -1164 26858 -1152 26892
rect -1210 26824 -1152 26858
rect -1210 26790 -1198 26824
rect -1164 26790 -1152 26824
rect -1210 26749 -1152 26790
rect -1052 27708 -994 27749
rect -1052 27674 -1040 27708
rect -1006 27674 -994 27708
rect -1052 27640 -994 27674
rect -1052 27606 -1040 27640
rect -1006 27606 -994 27640
rect -1052 27572 -994 27606
rect -1052 27538 -1040 27572
rect -1006 27538 -994 27572
rect -1052 27504 -994 27538
rect -1052 27470 -1040 27504
rect -1006 27470 -994 27504
rect -1052 27436 -994 27470
rect -1052 27402 -1040 27436
rect -1006 27402 -994 27436
rect -1052 27368 -994 27402
rect -1052 27334 -1040 27368
rect -1006 27334 -994 27368
rect -1052 27300 -994 27334
rect -1052 27266 -1040 27300
rect -1006 27266 -994 27300
rect -1052 27232 -994 27266
rect -1052 27198 -1040 27232
rect -1006 27198 -994 27232
rect -1052 27164 -994 27198
rect -1052 27130 -1040 27164
rect -1006 27130 -994 27164
rect -1052 27096 -994 27130
rect -1052 27062 -1040 27096
rect -1006 27062 -994 27096
rect -1052 27028 -994 27062
rect -1052 26994 -1040 27028
rect -1006 26994 -994 27028
rect -1052 26960 -994 26994
rect -1052 26926 -1040 26960
rect -1006 26926 -994 26960
rect -1052 26892 -994 26926
rect -1052 26858 -1040 26892
rect -1006 26858 -994 26892
rect -1052 26824 -994 26858
rect -1052 26790 -1040 26824
rect -1006 26790 -994 26824
rect -1052 26749 -994 26790
rect -894 27708 -836 27749
rect -894 27674 -882 27708
rect -848 27674 -836 27708
rect -894 27640 -836 27674
rect -894 27606 -882 27640
rect -848 27606 -836 27640
rect -894 27572 -836 27606
rect -894 27538 -882 27572
rect -848 27538 -836 27572
rect -894 27504 -836 27538
rect -894 27470 -882 27504
rect -848 27470 -836 27504
rect -894 27436 -836 27470
rect -894 27402 -882 27436
rect -848 27402 -836 27436
rect -894 27368 -836 27402
rect -894 27334 -882 27368
rect -848 27334 -836 27368
rect -894 27300 -836 27334
rect -894 27266 -882 27300
rect -848 27266 -836 27300
rect -894 27232 -836 27266
rect -894 27198 -882 27232
rect -848 27198 -836 27232
rect -894 27164 -836 27198
rect -894 27130 -882 27164
rect -848 27130 -836 27164
rect -894 27096 -836 27130
rect -894 27062 -882 27096
rect -848 27062 -836 27096
rect -894 27028 -836 27062
rect -894 26994 -882 27028
rect -848 26994 -836 27028
rect -894 26960 -836 26994
rect -894 26926 -882 26960
rect -848 26926 -836 26960
rect -894 26892 -836 26926
rect -894 26858 -882 26892
rect -848 26858 -836 26892
rect -894 26824 -836 26858
rect -894 26790 -882 26824
rect -848 26790 -836 26824
rect -894 26749 -836 26790
rect -736 27708 -678 27749
rect -736 27674 -724 27708
rect -690 27674 -678 27708
rect -736 27640 -678 27674
rect -736 27606 -724 27640
rect -690 27606 -678 27640
rect -736 27572 -678 27606
rect -736 27538 -724 27572
rect -690 27538 -678 27572
rect -736 27504 -678 27538
rect -736 27470 -724 27504
rect -690 27470 -678 27504
rect -736 27436 -678 27470
rect -736 27402 -724 27436
rect -690 27402 -678 27436
rect -736 27368 -678 27402
rect -736 27334 -724 27368
rect -690 27334 -678 27368
rect -736 27300 -678 27334
rect -736 27266 -724 27300
rect -690 27266 -678 27300
rect -736 27232 -678 27266
rect -736 27198 -724 27232
rect -690 27198 -678 27232
rect -736 27164 -678 27198
rect -736 27130 -724 27164
rect -690 27130 -678 27164
rect -736 27096 -678 27130
rect -736 27062 -724 27096
rect -690 27062 -678 27096
rect -736 27028 -678 27062
rect -736 26994 -724 27028
rect -690 26994 -678 27028
rect -736 26960 -678 26994
rect -736 26926 -724 26960
rect -690 26926 -678 26960
rect -736 26892 -678 26926
rect -736 26858 -724 26892
rect -690 26858 -678 26892
rect -736 26824 -678 26858
rect -736 26790 -724 26824
rect -690 26790 -678 26824
rect -736 26749 -678 26790
rect -578 27708 -520 27749
rect -578 27674 -566 27708
rect -532 27674 -520 27708
rect -578 27640 -520 27674
rect -578 27606 -566 27640
rect -532 27606 -520 27640
rect -578 27572 -520 27606
rect -578 27538 -566 27572
rect -532 27538 -520 27572
rect -578 27504 -520 27538
rect -578 27470 -566 27504
rect -532 27470 -520 27504
rect -578 27436 -520 27470
rect -578 27402 -566 27436
rect -532 27402 -520 27436
rect -578 27368 -520 27402
rect -578 27334 -566 27368
rect -532 27334 -520 27368
rect -578 27300 -520 27334
rect -578 27266 -566 27300
rect -532 27266 -520 27300
rect -578 27232 -520 27266
rect -578 27198 -566 27232
rect -532 27198 -520 27232
rect -578 27164 -520 27198
rect -578 27130 -566 27164
rect -532 27130 -520 27164
rect -578 27096 -520 27130
rect -578 27062 -566 27096
rect -532 27062 -520 27096
rect -578 27028 -520 27062
rect -578 26994 -566 27028
rect -532 26994 -520 27028
rect -578 26960 -520 26994
rect -578 26926 -566 26960
rect -532 26926 -520 26960
rect -578 26892 -520 26926
rect -578 26858 -566 26892
rect -532 26858 -520 26892
rect -578 26824 -520 26858
rect -578 26790 -566 26824
rect -532 26790 -520 26824
rect -578 26749 -520 26790
rect -420 27708 -362 27749
rect -420 27674 -408 27708
rect -374 27674 -362 27708
rect -420 27640 -362 27674
rect -420 27606 -408 27640
rect -374 27606 -362 27640
rect -420 27572 -362 27606
rect -420 27538 -408 27572
rect -374 27538 -362 27572
rect -420 27504 -362 27538
rect -420 27470 -408 27504
rect -374 27470 -362 27504
rect -420 27436 -362 27470
rect -420 27402 -408 27436
rect -374 27402 -362 27436
rect -420 27368 -362 27402
rect -420 27334 -408 27368
rect -374 27334 -362 27368
rect -420 27300 -362 27334
rect -420 27266 -408 27300
rect -374 27266 -362 27300
rect -420 27232 -362 27266
rect -420 27198 -408 27232
rect -374 27198 -362 27232
rect -420 27164 -362 27198
rect -420 27130 -408 27164
rect -374 27130 -362 27164
rect -420 27096 -362 27130
rect -420 27062 -408 27096
rect -374 27062 -362 27096
rect -420 27028 -362 27062
rect -420 26994 -408 27028
rect -374 26994 -362 27028
rect -420 26960 -362 26994
rect -420 26926 -408 26960
rect -374 26926 -362 26960
rect -420 26892 -362 26926
rect -420 26858 -408 26892
rect -374 26858 -362 26892
rect -420 26824 -362 26858
rect -420 26790 -408 26824
rect -374 26790 -362 26824
rect -420 26749 -362 26790
rect -262 27708 -204 27749
rect -262 27674 -250 27708
rect -216 27674 -204 27708
rect -262 27640 -204 27674
rect -262 27606 -250 27640
rect -216 27606 -204 27640
rect -262 27572 -204 27606
rect -262 27538 -250 27572
rect -216 27538 -204 27572
rect -262 27504 -204 27538
rect -262 27470 -250 27504
rect -216 27470 -204 27504
rect -262 27436 -204 27470
rect -262 27402 -250 27436
rect -216 27402 -204 27436
rect -262 27368 -204 27402
rect -262 27334 -250 27368
rect -216 27334 -204 27368
rect -262 27300 -204 27334
rect -262 27266 -250 27300
rect -216 27266 -204 27300
rect -262 27232 -204 27266
rect -262 27198 -250 27232
rect -216 27198 -204 27232
rect -262 27164 -204 27198
rect -262 27130 -250 27164
rect -216 27130 -204 27164
rect -262 27096 -204 27130
rect -262 27062 -250 27096
rect -216 27062 -204 27096
rect -262 27028 -204 27062
rect -262 26994 -250 27028
rect -216 26994 -204 27028
rect -262 26960 -204 26994
rect -262 26926 -250 26960
rect -216 26926 -204 26960
rect -262 26892 -204 26926
rect -262 26858 -250 26892
rect -216 26858 -204 26892
rect -262 26824 -204 26858
rect -262 26790 -250 26824
rect -216 26790 -204 26824
rect -262 26749 -204 26790
rect -104 27708 -46 27749
rect -104 27674 -92 27708
rect -58 27674 -46 27708
rect -104 27640 -46 27674
rect -104 27606 -92 27640
rect -58 27606 -46 27640
rect -104 27572 -46 27606
rect -104 27538 -92 27572
rect -58 27538 -46 27572
rect -104 27504 -46 27538
rect -104 27470 -92 27504
rect -58 27470 -46 27504
rect -104 27436 -46 27470
rect -104 27402 -92 27436
rect -58 27402 -46 27436
rect -104 27368 -46 27402
rect -104 27334 -92 27368
rect -58 27334 -46 27368
rect -104 27300 -46 27334
rect -104 27266 -92 27300
rect -58 27266 -46 27300
rect -104 27232 -46 27266
rect -104 27198 -92 27232
rect -58 27198 -46 27232
rect -104 27164 -46 27198
rect -104 27130 -92 27164
rect -58 27130 -46 27164
rect -104 27096 -46 27130
rect -104 27062 -92 27096
rect -58 27062 -46 27096
rect -104 27028 -46 27062
rect -104 26994 -92 27028
rect -58 26994 -46 27028
rect -104 26960 -46 26994
rect -104 26926 -92 26960
rect -58 26926 -46 26960
rect -104 26892 -46 26926
rect -104 26858 -92 26892
rect -58 26858 -46 26892
rect -104 26824 -46 26858
rect -104 26790 -92 26824
rect -58 26790 -46 26824
rect -104 26749 -46 26790
rect 54 27708 112 27749
rect 54 27674 66 27708
rect 100 27674 112 27708
rect 54 27640 112 27674
rect 54 27606 66 27640
rect 100 27606 112 27640
rect 54 27572 112 27606
rect 54 27538 66 27572
rect 100 27538 112 27572
rect 54 27504 112 27538
rect 54 27470 66 27504
rect 100 27470 112 27504
rect 54 27436 112 27470
rect 54 27402 66 27436
rect 100 27402 112 27436
rect 54 27368 112 27402
rect 54 27334 66 27368
rect 100 27334 112 27368
rect 54 27300 112 27334
rect 54 27266 66 27300
rect 100 27266 112 27300
rect 54 27232 112 27266
rect 54 27198 66 27232
rect 100 27198 112 27232
rect 54 27164 112 27198
rect 54 27130 66 27164
rect 100 27130 112 27164
rect 54 27096 112 27130
rect 54 27062 66 27096
rect 100 27062 112 27096
rect 54 27028 112 27062
rect 54 26994 66 27028
rect 100 26994 112 27028
rect 54 26960 112 26994
rect 54 26926 66 26960
rect 100 26926 112 26960
rect 54 26892 112 26926
rect 54 26858 66 26892
rect 100 26858 112 26892
rect 54 26824 112 26858
rect 54 26790 66 26824
rect 100 26790 112 26824
rect 54 26749 112 26790
rect 212 27708 270 27749
rect 212 27674 224 27708
rect 258 27674 270 27708
rect 212 27640 270 27674
rect 212 27606 224 27640
rect 258 27606 270 27640
rect 212 27572 270 27606
rect 212 27538 224 27572
rect 258 27538 270 27572
rect 212 27504 270 27538
rect 212 27470 224 27504
rect 258 27470 270 27504
rect 212 27436 270 27470
rect 212 27402 224 27436
rect 258 27402 270 27436
rect 212 27368 270 27402
rect 212 27334 224 27368
rect 258 27334 270 27368
rect 212 27300 270 27334
rect 212 27266 224 27300
rect 258 27266 270 27300
rect 212 27232 270 27266
rect 212 27198 224 27232
rect 258 27198 270 27232
rect 212 27164 270 27198
rect 212 27130 224 27164
rect 258 27130 270 27164
rect 212 27096 270 27130
rect 212 27062 224 27096
rect 258 27062 270 27096
rect 212 27028 270 27062
rect 212 26994 224 27028
rect 258 26994 270 27028
rect 212 26960 270 26994
rect 212 26926 224 26960
rect 258 26926 270 26960
rect 212 26892 270 26926
rect 212 26858 224 26892
rect 258 26858 270 26892
rect 212 26824 270 26858
rect 212 26790 224 26824
rect 258 26790 270 26824
rect 212 26749 270 26790
rect 370 27708 428 27749
rect 370 27674 382 27708
rect 416 27674 428 27708
rect 370 27640 428 27674
rect 370 27606 382 27640
rect 416 27606 428 27640
rect 370 27572 428 27606
rect 370 27538 382 27572
rect 416 27538 428 27572
rect 370 27504 428 27538
rect 370 27470 382 27504
rect 416 27470 428 27504
rect 370 27436 428 27470
rect 370 27402 382 27436
rect 416 27402 428 27436
rect 370 27368 428 27402
rect 370 27334 382 27368
rect 416 27334 428 27368
rect 370 27300 428 27334
rect 370 27266 382 27300
rect 416 27266 428 27300
rect 370 27232 428 27266
rect 370 27198 382 27232
rect 416 27198 428 27232
rect 370 27164 428 27198
rect 370 27130 382 27164
rect 416 27130 428 27164
rect 370 27096 428 27130
rect 370 27062 382 27096
rect 416 27062 428 27096
rect 370 27028 428 27062
rect 370 26994 382 27028
rect 416 26994 428 27028
rect 370 26960 428 26994
rect 370 26926 382 26960
rect 416 26926 428 26960
rect 370 26892 428 26926
rect 370 26858 382 26892
rect 416 26858 428 26892
rect 370 26824 428 26858
rect 370 26790 382 26824
rect 416 26790 428 26824
rect 370 26749 428 26790
rect 528 27708 586 27749
rect 528 27674 540 27708
rect 574 27674 586 27708
rect 528 27640 586 27674
rect 528 27606 540 27640
rect 574 27606 586 27640
rect 528 27572 586 27606
rect 528 27538 540 27572
rect 574 27538 586 27572
rect 528 27504 586 27538
rect 528 27470 540 27504
rect 574 27470 586 27504
rect 528 27436 586 27470
rect 528 27402 540 27436
rect 574 27402 586 27436
rect 528 27368 586 27402
rect 528 27334 540 27368
rect 574 27334 586 27368
rect 528 27300 586 27334
rect 528 27266 540 27300
rect 574 27266 586 27300
rect 528 27232 586 27266
rect 528 27198 540 27232
rect 574 27198 586 27232
rect 528 27164 586 27198
rect 528 27130 540 27164
rect 574 27130 586 27164
rect 528 27096 586 27130
rect 528 27062 540 27096
rect 574 27062 586 27096
rect 528 27028 586 27062
rect 528 26994 540 27028
rect 574 26994 586 27028
rect 528 26960 586 26994
rect 528 26926 540 26960
rect 574 26926 586 26960
rect 528 26892 586 26926
rect 528 26858 540 26892
rect 574 26858 586 26892
rect 528 26824 586 26858
rect 528 26790 540 26824
rect 574 26790 586 26824
rect 528 26749 586 26790
rect 686 27708 744 27749
rect 686 27674 698 27708
rect 732 27674 744 27708
rect 686 27640 744 27674
rect 686 27606 698 27640
rect 732 27606 744 27640
rect 686 27572 744 27606
rect 686 27538 698 27572
rect 732 27538 744 27572
rect 686 27504 744 27538
rect 686 27470 698 27504
rect 732 27470 744 27504
rect 686 27436 744 27470
rect 686 27402 698 27436
rect 732 27402 744 27436
rect 686 27368 744 27402
rect 686 27334 698 27368
rect 732 27334 744 27368
rect 686 27300 744 27334
rect 686 27266 698 27300
rect 732 27266 744 27300
rect 686 27232 744 27266
rect 686 27198 698 27232
rect 732 27198 744 27232
rect 686 27164 744 27198
rect 686 27130 698 27164
rect 732 27130 744 27164
rect 686 27096 744 27130
rect 686 27062 698 27096
rect 732 27062 744 27096
rect 686 27028 744 27062
rect 686 26994 698 27028
rect 732 26994 744 27028
rect 686 26960 744 26994
rect 686 26926 698 26960
rect 732 26926 744 26960
rect 686 26892 744 26926
rect 686 26858 698 26892
rect 732 26858 744 26892
rect 686 26824 744 26858
rect 686 26790 698 26824
rect 732 26790 744 26824
rect 686 26749 744 26790
rect 844 27708 902 27749
rect 844 27674 856 27708
rect 890 27674 902 27708
rect 844 27640 902 27674
rect 844 27606 856 27640
rect 890 27606 902 27640
rect 844 27572 902 27606
rect 844 27538 856 27572
rect 890 27538 902 27572
rect 844 27504 902 27538
rect 844 27470 856 27504
rect 890 27470 902 27504
rect 844 27436 902 27470
rect 844 27402 856 27436
rect 890 27402 902 27436
rect 844 27368 902 27402
rect 844 27334 856 27368
rect 890 27334 902 27368
rect 844 27300 902 27334
rect 844 27266 856 27300
rect 890 27266 902 27300
rect 844 27232 902 27266
rect 844 27198 856 27232
rect 890 27198 902 27232
rect 844 27164 902 27198
rect 844 27130 856 27164
rect 890 27130 902 27164
rect 844 27096 902 27130
rect 844 27062 856 27096
rect 890 27062 902 27096
rect 844 27028 902 27062
rect 844 26994 856 27028
rect 890 26994 902 27028
rect 844 26960 902 26994
rect 844 26926 856 26960
rect 890 26926 902 26960
rect 844 26892 902 26926
rect 844 26858 856 26892
rect 890 26858 902 26892
rect 844 26824 902 26858
rect 844 26790 856 26824
rect 890 26790 902 26824
rect 844 26749 902 26790
rect 1002 27708 1060 27749
rect 1002 27674 1014 27708
rect 1048 27674 1060 27708
rect 1002 27640 1060 27674
rect 1002 27606 1014 27640
rect 1048 27606 1060 27640
rect 1002 27572 1060 27606
rect 1002 27538 1014 27572
rect 1048 27538 1060 27572
rect 1002 27504 1060 27538
rect 1002 27470 1014 27504
rect 1048 27470 1060 27504
rect 1002 27436 1060 27470
rect 1002 27402 1014 27436
rect 1048 27402 1060 27436
rect 1002 27368 1060 27402
rect 1002 27334 1014 27368
rect 1048 27334 1060 27368
rect 1002 27300 1060 27334
rect 1002 27266 1014 27300
rect 1048 27266 1060 27300
rect 1002 27232 1060 27266
rect 1002 27198 1014 27232
rect 1048 27198 1060 27232
rect 1002 27164 1060 27198
rect 1002 27130 1014 27164
rect 1048 27130 1060 27164
rect 1002 27096 1060 27130
rect 1002 27062 1014 27096
rect 1048 27062 1060 27096
rect 1002 27028 1060 27062
rect 1002 26994 1014 27028
rect 1048 26994 1060 27028
rect 1002 26960 1060 26994
rect 1002 26926 1014 26960
rect 1048 26926 1060 26960
rect 1002 26892 1060 26926
rect 1002 26858 1014 26892
rect 1048 26858 1060 26892
rect 1002 26824 1060 26858
rect 1002 26790 1014 26824
rect 1048 26790 1060 26824
rect 1002 26749 1060 26790
rect 1160 27708 1218 27749
rect 1160 27674 1172 27708
rect 1206 27674 1218 27708
rect 1160 27640 1218 27674
rect 1160 27606 1172 27640
rect 1206 27606 1218 27640
rect 1160 27572 1218 27606
rect 1160 27538 1172 27572
rect 1206 27538 1218 27572
rect 1160 27504 1218 27538
rect 1160 27470 1172 27504
rect 1206 27470 1218 27504
rect 1160 27436 1218 27470
rect 1160 27402 1172 27436
rect 1206 27402 1218 27436
rect 1160 27368 1218 27402
rect 1160 27334 1172 27368
rect 1206 27334 1218 27368
rect 1160 27300 1218 27334
rect 1160 27266 1172 27300
rect 1206 27266 1218 27300
rect 1160 27232 1218 27266
rect 1160 27198 1172 27232
rect 1206 27198 1218 27232
rect 1160 27164 1218 27198
rect 1160 27130 1172 27164
rect 1206 27130 1218 27164
rect 1160 27096 1218 27130
rect 1160 27062 1172 27096
rect 1206 27062 1218 27096
rect 1160 27028 1218 27062
rect 1160 26994 1172 27028
rect 1206 26994 1218 27028
rect 1160 26960 1218 26994
rect 1160 26926 1172 26960
rect 1206 26926 1218 26960
rect 1160 26892 1218 26926
rect 1160 26858 1172 26892
rect 1206 26858 1218 26892
rect 1160 26824 1218 26858
rect 1160 26790 1172 26824
rect 1206 26790 1218 26824
rect 1160 26749 1218 26790
rect 1318 27708 1376 27749
rect 1318 27674 1330 27708
rect 1364 27674 1376 27708
rect 1318 27640 1376 27674
rect 1318 27606 1330 27640
rect 1364 27606 1376 27640
rect 1318 27572 1376 27606
rect 1318 27538 1330 27572
rect 1364 27538 1376 27572
rect 1318 27504 1376 27538
rect 1318 27470 1330 27504
rect 1364 27470 1376 27504
rect 1318 27436 1376 27470
rect 1318 27402 1330 27436
rect 1364 27402 1376 27436
rect 1318 27368 1376 27402
rect 1318 27334 1330 27368
rect 1364 27334 1376 27368
rect 1318 27300 1376 27334
rect 1318 27266 1330 27300
rect 1364 27266 1376 27300
rect 1318 27232 1376 27266
rect 1318 27198 1330 27232
rect 1364 27198 1376 27232
rect 1318 27164 1376 27198
rect 1318 27130 1330 27164
rect 1364 27130 1376 27164
rect 1318 27096 1376 27130
rect 1318 27062 1330 27096
rect 1364 27062 1376 27096
rect 1318 27028 1376 27062
rect 1318 26994 1330 27028
rect 1364 26994 1376 27028
rect 1318 26960 1376 26994
rect 1318 26926 1330 26960
rect 1364 26926 1376 26960
rect 1318 26892 1376 26926
rect 1318 26858 1330 26892
rect 1364 26858 1376 26892
rect 1318 26824 1376 26858
rect 1318 26790 1330 26824
rect 1364 26790 1376 26824
rect 1318 26749 1376 26790
rect 1476 27708 1534 27749
rect 1476 27674 1488 27708
rect 1522 27674 1534 27708
rect 1476 27640 1534 27674
rect 1476 27606 1488 27640
rect 1522 27606 1534 27640
rect 1476 27572 1534 27606
rect 1476 27538 1488 27572
rect 1522 27538 1534 27572
rect 1476 27504 1534 27538
rect 1476 27470 1488 27504
rect 1522 27470 1534 27504
rect 1476 27436 1534 27470
rect 1476 27402 1488 27436
rect 1522 27402 1534 27436
rect 1476 27368 1534 27402
rect 1476 27334 1488 27368
rect 1522 27334 1534 27368
rect 1476 27300 1534 27334
rect 1476 27266 1488 27300
rect 1522 27266 1534 27300
rect 1476 27232 1534 27266
rect 1476 27198 1488 27232
rect 1522 27198 1534 27232
rect 1476 27164 1534 27198
rect 1476 27130 1488 27164
rect 1522 27130 1534 27164
rect 1476 27096 1534 27130
rect 1476 27062 1488 27096
rect 1522 27062 1534 27096
rect 1476 27028 1534 27062
rect 1476 26994 1488 27028
rect 1522 26994 1534 27028
rect 1476 26960 1534 26994
rect 1476 26926 1488 26960
rect 1522 26926 1534 26960
rect 1476 26892 1534 26926
rect 1476 26858 1488 26892
rect 1522 26858 1534 26892
rect 1476 26824 1534 26858
rect 1476 26790 1488 26824
rect 1522 26790 1534 26824
rect 1476 26749 1534 26790
rect 1634 27708 1692 27749
rect 1634 27674 1646 27708
rect 1680 27674 1692 27708
rect 1634 27640 1692 27674
rect 1634 27606 1646 27640
rect 1680 27606 1692 27640
rect 1634 27572 1692 27606
rect 1634 27538 1646 27572
rect 1680 27538 1692 27572
rect 1634 27504 1692 27538
rect 1634 27470 1646 27504
rect 1680 27470 1692 27504
rect 1634 27436 1692 27470
rect 1634 27402 1646 27436
rect 1680 27402 1692 27436
rect 1634 27368 1692 27402
rect 1634 27334 1646 27368
rect 1680 27334 1692 27368
rect 1634 27300 1692 27334
rect 1634 27266 1646 27300
rect 1680 27266 1692 27300
rect 1634 27232 1692 27266
rect 1634 27198 1646 27232
rect 1680 27198 1692 27232
rect 1634 27164 1692 27198
rect 1634 27130 1646 27164
rect 1680 27130 1692 27164
rect 1634 27096 1692 27130
rect 1634 27062 1646 27096
rect 1680 27062 1692 27096
rect 1634 27028 1692 27062
rect 1634 26994 1646 27028
rect 1680 26994 1692 27028
rect 1634 26960 1692 26994
rect 1634 26926 1646 26960
rect 1680 26926 1692 26960
rect 1634 26892 1692 26926
rect 1634 26858 1646 26892
rect 1680 26858 1692 26892
rect 1634 26824 1692 26858
rect 1634 26790 1646 26824
rect 1680 26790 1692 26824
rect 1634 26749 1692 26790
rect -3591 19432 -2591 19444
rect -3591 19398 -3579 19432
rect -2603 19398 -2591 19432
rect -3591 19386 -2591 19398
rect -2355 19432 -1355 19444
rect -2355 19398 -2343 19432
rect -1367 19398 -1355 19432
rect -2355 19386 -1355 19398
rect -1119 19432 -119 19444
rect -1119 19398 -1107 19432
rect -131 19398 -119 19432
rect -1119 19386 -119 19398
rect 117 19432 1117 19444
rect 117 19398 129 19432
rect 1105 19398 1117 19432
rect 117 19386 1117 19398
rect 1353 19432 2353 19444
rect 1353 19398 1365 19432
rect 2341 19398 2353 19432
rect 1353 19386 2353 19398
rect 2589 19432 3589 19444
rect 2589 19398 2601 19432
rect 3577 19398 3589 19432
rect 2589 19386 3589 19398
rect -3591 19174 -2591 19186
rect -3591 19140 -3579 19174
rect -2603 19140 -2591 19174
rect -3591 19128 -2591 19140
rect -2355 19174 -1355 19186
rect -2355 19140 -2343 19174
rect -1367 19140 -1355 19174
rect -2355 19128 -1355 19140
rect -1119 19174 -119 19186
rect -1119 19140 -1107 19174
rect -131 19140 -119 19174
rect -1119 19128 -119 19140
rect 117 19174 1117 19186
rect 117 19140 129 19174
rect 1105 19140 1117 19174
rect 117 19128 1117 19140
rect 1353 19174 2353 19186
rect 1353 19140 1365 19174
rect 2341 19140 2353 19174
rect 1353 19128 2353 19140
rect 2589 19174 3589 19186
rect 2589 19140 2601 19174
rect 3577 19140 3589 19174
rect 2589 19128 3589 19140
rect -3591 18842 -2591 18854
rect -3591 18808 -3579 18842
rect -2603 18808 -2591 18842
rect -3591 18796 -2591 18808
rect -2355 18842 -1355 18854
rect -2355 18808 -2343 18842
rect -1367 18808 -1355 18842
rect -2355 18796 -1355 18808
rect -1119 18842 -119 18854
rect -1119 18808 -1107 18842
rect -131 18808 -119 18842
rect -1119 18796 -119 18808
rect 117 18842 1117 18854
rect 117 18808 129 18842
rect 1105 18808 1117 18842
rect 117 18796 1117 18808
rect 1353 18842 2353 18854
rect 1353 18808 1365 18842
rect 2341 18808 2353 18842
rect 1353 18796 2353 18808
rect 2589 18842 3589 18854
rect 2589 18808 2601 18842
rect 3577 18808 3589 18842
rect 2589 18796 3589 18808
rect -3591 18584 -2591 18596
rect -3591 18550 -3579 18584
rect -2603 18550 -2591 18584
rect -3591 18538 -2591 18550
rect -2355 18584 -1355 18596
rect -2355 18550 -2343 18584
rect -1367 18550 -1355 18584
rect -2355 18538 -1355 18550
rect -1119 18584 -119 18596
rect -1119 18550 -1107 18584
rect -131 18550 -119 18584
rect -1119 18538 -119 18550
rect 117 18584 1117 18596
rect 117 18550 129 18584
rect 1105 18550 1117 18584
rect 117 18538 1117 18550
rect 1353 18584 2353 18596
rect 1353 18550 1365 18584
rect 2341 18550 2353 18584
rect 1353 18538 2353 18550
rect 2589 18584 3589 18596
rect 2589 18550 2601 18584
rect 3577 18550 3589 18584
rect 2589 18538 3589 18550
<< ndiffc >>
rect -571 26106 -537 26140
rect -571 26038 -537 26072
rect -571 25970 -537 26004
rect -571 25902 -537 25936
rect -571 25834 -537 25868
rect -571 25766 -537 25800
rect -571 25698 -537 25732
rect -571 25630 -537 25664
rect -571 25562 -537 25596
rect -571 25494 -537 25528
rect -571 25426 -537 25460
rect -571 25358 -537 25392
rect -571 25290 -537 25324
rect -571 25222 -537 25256
rect -413 26106 -379 26140
rect -413 26038 -379 26072
rect -413 25970 -379 26004
rect -413 25902 -379 25936
rect -413 25834 -379 25868
rect -413 25766 -379 25800
rect -413 25698 -379 25732
rect -413 25630 -379 25664
rect -413 25562 -379 25596
rect -413 25494 -379 25528
rect -413 25426 -379 25460
rect -413 25358 -379 25392
rect -413 25290 -379 25324
rect -413 25222 -379 25256
rect -255 26106 -221 26140
rect -255 26038 -221 26072
rect -255 25970 -221 26004
rect -255 25902 -221 25936
rect -255 25834 -221 25868
rect -255 25766 -221 25800
rect -255 25698 -221 25732
rect -255 25630 -221 25664
rect -255 25562 -221 25596
rect -255 25494 -221 25528
rect -255 25426 -221 25460
rect -255 25358 -221 25392
rect -255 25290 -221 25324
rect -255 25222 -221 25256
rect -97 26106 -63 26140
rect -97 26038 -63 26072
rect -97 25970 -63 26004
rect -97 25902 -63 25936
rect -97 25834 -63 25868
rect -97 25766 -63 25800
rect -97 25698 -63 25732
rect -97 25630 -63 25664
rect -97 25562 -63 25596
rect -97 25494 -63 25528
rect -97 25426 -63 25460
rect -97 25358 -63 25392
rect -97 25290 -63 25324
rect -97 25222 -63 25256
rect 61 26106 95 26140
rect 61 26038 95 26072
rect 61 25970 95 26004
rect 61 25902 95 25936
rect 61 25834 95 25868
rect 61 25766 95 25800
rect 61 25698 95 25732
rect 61 25630 95 25664
rect 61 25562 95 25596
rect 61 25494 95 25528
rect 61 25426 95 25460
rect 61 25358 95 25392
rect 61 25290 95 25324
rect 61 25222 95 25256
rect 219 26106 253 26140
rect 219 26038 253 26072
rect 219 25970 253 26004
rect 219 25902 253 25936
rect 219 25834 253 25868
rect 219 25766 253 25800
rect 219 25698 253 25732
rect 219 25630 253 25664
rect 219 25562 253 25596
rect 219 25494 253 25528
rect 219 25426 253 25460
rect 219 25358 253 25392
rect 219 25290 253 25324
rect 219 25222 253 25256
rect 377 26106 411 26140
rect 377 26038 411 26072
rect 377 25970 411 26004
rect 377 25902 411 25936
rect 377 25834 411 25868
rect 377 25766 411 25800
rect 377 25698 411 25732
rect 377 25630 411 25664
rect 377 25562 411 25596
rect 377 25494 411 25528
rect 377 25426 411 25460
rect 377 25358 411 25392
rect 377 25290 411 25324
rect 377 25222 411 25256
rect 535 26106 569 26140
rect 535 26038 569 26072
rect 535 25970 569 26004
rect 535 25902 569 25936
rect 535 25834 569 25868
rect 535 25766 569 25800
rect 535 25698 569 25732
rect 535 25630 569 25664
rect 535 25562 569 25596
rect 535 25494 569 25528
rect 535 25426 569 25460
rect 535 25358 569 25392
rect 535 25290 569 25324
rect 535 25222 569 25256
rect -571 24586 -537 24620
rect -571 24518 -537 24552
rect -571 24450 -537 24484
rect -571 24382 -537 24416
rect -571 24314 -537 24348
rect -571 24246 -537 24280
rect -571 24178 -537 24212
rect -571 24110 -537 24144
rect -571 24042 -537 24076
rect -571 23974 -537 24008
rect -571 23906 -537 23940
rect -571 23838 -537 23872
rect -571 23770 -537 23804
rect -571 23702 -537 23736
rect -413 24586 -379 24620
rect -413 24518 -379 24552
rect -413 24450 -379 24484
rect -413 24382 -379 24416
rect -413 24314 -379 24348
rect -413 24246 -379 24280
rect -413 24178 -379 24212
rect -413 24110 -379 24144
rect -413 24042 -379 24076
rect -413 23974 -379 24008
rect -413 23906 -379 23940
rect -413 23838 -379 23872
rect -413 23770 -379 23804
rect -413 23702 -379 23736
rect -255 24586 -221 24620
rect -255 24518 -221 24552
rect -255 24450 -221 24484
rect -255 24382 -221 24416
rect -255 24314 -221 24348
rect -255 24246 -221 24280
rect -255 24178 -221 24212
rect -255 24110 -221 24144
rect -255 24042 -221 24076
rect -255 23974 -221 24008
rect -255 23906 -221 23940
rect -255 23838 -221 23872
rect -255 23770 -221 23804
rect -255 23702 -221 23736
rect -97 24586 -63 24620
rect -97 24518 -63 24552
rect -97 24450 -63 24484
rect -97 24382 -63 24416
rect -97 24314 -63 24348
rect -97 24246 -63 24280
rect -97 24178 -63 24212
rect -97 24110 -63 24144
rect -97 24042 -63 24076
rect -97 23974 -63 24008
rect -97 23906 -63 23940
rect -97 23838 -63 23872
rect -97 23770 -63 23804
rect -97 23702 -63 23736
rect 61 24586 95 24620
rect 61 24518 95 24552
rect 61 24450 95 24484
rect 61 24382 95 24416
rect 61 24314 95 24348
rect 61 24246 95 24280
rect 61 24178 95 24212
rect 61 24110 95 24144
rect 61 24042 95 24076
rect 61 23974 95 24008
rect 61 23906 95 23940
rect 61 23838 95 23872
rect 61 23770 95 23804
rect 61 23702 95 23736
rect 219 24586 253 24620
rect 219 24518 253 24552
rect 219 24450 253 24484
rect 219 24382 253 24416
rect 219 24314 253 24348
rect 219 24246 253 24280
rect 219 24178 253 24212
rect 219 24110 253 24144
rect 219 24042 253 24076
rect 219 23974 253 24008
rect 219 23906 253 23940
rect 219 23838 253 23872
rect 219 23770 253 23804
rect 219 23702 253 23736
rect 377 24586 411 24620
rect 377 24518 411 24552
rect 377 24450 411 24484
rect 377 24382 411 24416
rect 377 24314 411 24348
rect 377 24246 411 24280
rect 377 24178 411 24212
rect 377 24110 411 24144
rect 377 24042 411 24076
rect 377 23974 411 24008
rect 377 23906 411 23940
rect 377 23838 411 23872
rect 377 23770 411 23804
rect 377 23702 411 23736
rect 535 24586 569 24620
rect 535 24518 569 24552
rect 535 24450 569 24484
rect 535 24382 569 24416
rect 535 24314 569 24348
rect 535 24246 569 24280
rect 535 24178 569 24212
rect 535 24110 569 24144
rect 535 24042 569 24076
rect 535 23974 569 24008
rect 535 23906 569 23940
rect 535 23838 569 23872
rect 535 23770 569 23804
rect 535 23702 569 23736
rect -1562 23065 -1528 23099
rect -1562 22997 -1528 23031
rect -1562 22929 -1528 22963
rect -1562 22861 -1528 22895
rect -1562 22793 -1528 22827
rect -1562 22725 -1528 22759
rect -1562 22657 -1528 22691
rect -1562 22589 -1528 22623
rect -1562 22521 -1528 22555
rect -1562 22453 -1528 22487
rect -1562 22385 -1528 22419
rect -1562 22317 -1528 22351
rect -1562 22249 -1528 22283
rect -1562 22181 -1528 22215
rect -1304 23065 -1270 23099
rect -1304 22997 -1270 23031
rect -1304 22929 -1270 22963
rect -1304 22861 -1270 22895
rect -1304 22793 -1270 22827
rect -1304 22725 -1270 22759
rect -1304 22657 -1270 22691
rect -1304 22589 -1270 22623
rect -1304 22521 -1270 22555
rect -1304 22453 -1270 22487
rect -1304 22385 -1270 22419
rect -1304 22317 -1270 22351
rect -1304 22249 -1270 22283
rect -1304 22181 -1270 22215
rect -1046 23065 -1012 23099
rect -1046 22997 -1012 23031
rect -1046 22929 -1012 22963
rect -1046 22861 -1012 22895
rect -1046 22793 -1012 22827
rect -1046 22725 -1012 22759
rect -1046 22657 -1012 22691
rect -1046 22589 -1012 22623
rect -1046 22521 -1012 22555
rect -1046 22453 -1012 22487
rect -1046 22385 -1012 22419
rect -1046 22317 -1012 22351
rect -1046 22249 -1012 22283
rect -1046 22181 -1012 22215
rect -788 23065 -754 23099
rect -788 22997 -754 23031
rect -788 22929 -754 22963
rect -788 22861 -754 22895
rect -788 22793 -754 22827
rect -788 22725 -754 22759
rect -788 22657 -754 22691
rect -788 22589 -754 22623
rect -788 22521 -754 22555
rect -788 22453 -754 22487
rect -788 22385 -754 22419
rect -788 22317 -754 22351
rect -788 22249 -754 22283
rect -788 22181 -754 22215
rect -530 23065 -496 23099
rect -530 22997 -496 23031
rect -530 22929 -496 22963
rect -530 22861 -496 22895
rect -530 22793 -496 22827
rect -530 22725 -496 22759
rect -530 22657 -496 22691
rect -530 22589 -496 22623
rect -530 22521 -496 22555
rect -530 22453 -496 22487
rect -530 22385 -496 22419
rect -530 22317 -496 22351
rect -530 22249 -496 22283
rect -530 22181 -496 22215
rect -272 23065 -238 23099
rect -272 22997 -238 23031
rect -272 22929 -238 22963
rect -272 22861 -238 22895
rect -272 22793 -238 22827
rect -272 22725 -238 22759
rect -272 22657 -238 22691
rect -272 22589 -238 22623
rect -272 22521 -238 22555
rect -272 22453 -238 22487
rect -272 22385 -238 22419
rect -272 22317 -238 22351
rect -272 22249 -238 22283
rect -272 22181 -238 22215
rect -14 23065 20 23099
rect -14 22997 20 23031
rect -14 22929 20 22963
rect -14 22861 20 22895
rect -14 22793 20 22827
rect -14 22725 20 22759
rect -14 22657 20 22691
rect -14 22589 20 22623
rect -14 22521 20 22555
rect -14 22453 20 22487
rect -14 22385 20 22419
rect -14 22317 20 22351
rect -14 22249 20 22283
rect -14 22181 20 22215
rect 244 23065 278 23099
rect 244 22997 278 23031
rect 244 22929 278 22963
rect 244 22861 278 22895
rect 244 22793 278 22827
rect 244 22725 278 22759
rect 244 22657 278 22691
rect 244 22589 278 22623
rect 244 22521 278 22555
rect 244 22453 278 22487
rect 244 22385 278 22419
rect 244 22317 278 22351
rect 244 22249 278 22283
rect 244 22181 278 22215
rect 502 23065 536 23099
rect 502 22997 536 23031
rect 502 22929 536 22963
rect 502 22861 536 22895
rect 502 22793 536 22827
rect 502 22725 536 22759
rect 502 22657 536 22691
rect 502 22589 536 22623
rect 502 22521 536 22555
rect 502 22453 536 22487
rect 502 22385 536 22419
rect 502 22317 536 22351
rect 502 22249 536 22283
rect 502 22181 536 22215
rect 760 23065 794 23099
rect 760 22997 794 23031
rect 760 22929 794 22963
rect 760 22861 794 22895
rect 760 22793 794 22827
rect 760 22725 794 22759
rect 760 22657 794 22691
rect 760 22589 794 22623
rect 760 22521 794 22555
rect 760 22453 794 22487
rect 760 22385 794 22419
rect 760 22317 794 22351
rect 760 22249 794 22283
rect 760 22181 794 22215
rect 1018 23065 1052 23099
rect 1018 22997 1052 23031
rect 1018 22929 1052 22963
rect 1018 22861 1052 22895
rect 1018 22793 1052 22827
rect 1018 22725 1052 22759
rect 1018 22657 1052 22691
rect 1018 22589 1052 22623
rect 1018 22521 1052 22555
rect 1018 22453 1052 22487
rect 1018 22385 1052 22419
rect 1018 22317 1052 22351
rect 1018 22249 1052 22283
rect 1018 22181 1052 22215
rect 1276 23065 1310 23099
rect 1276 22997 1310 23031
rect 1276 22929 1310 22963
rect 1276 22861 1310 22895
rect 1276 22793 1310 22827
rect 1276 22725 1310 22759
rect 1276 22657 1310 22691
rect 1276 22589 1310 22623
rect 1276 22521 1310 22555
rect 1276 22453 1310 22487
rect 1276 22385 1310 22419
rect 1276 22317 1310 22351
rect 1276 22249 1310 22283
rect 1276 22181 1310 22215
rect 1534 23065 1568 23099
rect 1534 22997 1568 23031
rect 1534 22929 1568 22963
rect 1534 22861 1568 22895
rect 1534 22793 1568 22827
rect 1534 22725 1568 22759
rect 1534 22657 1568 22691
rect 1534 22589 1568 22623
rect 1534 22521 1568 22555
rect 1534 22453 1568 22487
rect 1534 22385 1568 22419
rect 1534 22317 1568 22351
rect 1534 22249 1568 22283
rect 1534 22181 1568 22215
rect -1822 21545 -1788 21579
rect -1822 21477 -1788 21511
rect -1822 21409 -1788 21443
rect -1822 21341 -1788 21375
rect -1822 21273 -1788 21307
rect -1822 21205 -1788 21239
rect -1822 21137 -1788 21171
rect -1822 21069 -1788 21103
rect -1822 21001 -1788 21035
rect -1822 20933 -1788 20967
rect -1822 20865 -1788 20899
rect -1822 20797 -1788 20831
rect -1822 20729 -1788 20763
rect -1822 20661 -1788 20695
rect -1564 21545 -1530 21579
rect -1564 21477 -1530 21511
rect -1564 21409 -1530 21443
rect -1564 21341 -1530 21375
rect -1564 21273 -1530 21307
rect -1564 21205 -1530 21239
rect -1564 21137 -1530 21171
rect -1564 21069 -1530 21103
rect -1564 21001 -1530 21035
rect -1564 20933 -1530 20967
rect -1564 20865 -1530 20899
rect -1564 20797 -1530 20831
rect -1564 20729 -1530 20763
rect -1564 20661 -1530 20695
rect -1306 21545 -1272 21579
rect -1306 21477 -1272 21511
rect -1306 21409 -1272 21443
rect -1306 21341 -1272 21375
rect -1306 21273 -1272 21307
rect -1306 21205 -1272 21239
rect -1306 21137 -1272 21171
rect -1306 21069 -1272 21103
rect -1306 21001 -1272 21035
rect -1306 20933 -1272 20967
rect -1306 20865 -1272 20899
rect -1306 20797 -1272 20831
rect -1306 20729 -1272 20763
rect -1306 20661 -1272 20695
rect -1048 21545 -1014 21579
rect -1048 21477 -1014 21511
rect -1048 21409 -1014 21443
rect -1048 21341 -1014 21375
rect -1048 21273 -1014 21307
rect -1048 21205 -1014 21239
rect -1048 21137 -1014 21171
rect -1048 21069 -1014 21103
rect -1048 21001 -1014 21035
rect -1048 20933 -1014 20967
rect -1048 20865 -1014 20899
rect -1048 20797 -1014 20831
rect -1048 20729 -1014 20763
rect -1048 20661 -1014 20695
rect -790 21545 -756 21579
rect -790 21477 -756 21511
rect -790 21409 -756 21443
rect -790 21341 -756 21375
rect -790 21273 -756 21307
rect -790 21205 -756 21239
rect -790 21137 -756 21171
rect -790 21069 -756 21103
rect -790 21001 -756 21035
rect -790 20933 -756 20967
rect -790 20865 -756 20899
rect -790 20797 -756 20831
rect -790 20729 -756 20763
rect -790 20661 -756 20695
rect -532 21545 -498 21579
rect -532 21477 -498 21511
rect -532 21409 -498 21443
rect -532 21341 -498 21375
rect -532 21273 -498 21307
rect -532 21205 -498 21239
rect -532 21137 -498 21171
rect -532 21069 -498 21103
rect -532 21001 -498 21035
rect -532 20933 -498 20967
rect -532 20865 -498 20899
rect -532 20797 -498 20831
rect -532 20729 -498 20763
rect -532 20661 -498 20695
rect -274 21545 -240 21579
rect -274 21477 -240 21511
rect -274 21409 -240 21443
rect -274 21341 -240 21375
rect -274 21273 -240 21307
rect -274 21205 -240 21239
rect -274 21137 -240 21171
rect -274 21069 -240 21103
rect -274 21001 -240 21035
rect -274 20933 -240 20967
rect -274 20865 -240 20899
rect -274 20797 -240 20831
rect -274 20729 -240 20763
rect -274 20661 -240 20695
rect -16 21545 18 21579
rect -16 21477 18 21511
rect -16 21409 18 21443
rect -16 21341 18 21375
rect -16 21273 18 21307
rect -16 21205 18 21239
rect -16 21137 18 21171
rect -16 21069 18 21103
rect -16 21001 18 21035
rect -16 20933 18 20967
rect -16 20865 18 20899
rect -16 20797 18 20831
rect -16 20729 18 20763
rect -16 20661 18 20695
rect 242 21545 276 21579
rect 242 21477 276 21511
rect 242 21409 276 21443
rect 242 21341 276 21375
rect 242 21273 276 21307
rect 242 21205 276 21239
rect 242 21137 276 21171
rect 242 21069 276 21103
rect 242 21001 276 21035
rect 242 20933 276 20967
rect 242 20865 276 20899
rect 242 20797 276 20831
rect 242 20729 276 20763
rect 242 20661 276 20695
rect 500 21545 534 21579
rect 500 21477 534 21511
rect 500 21409 534 21443
rect 500 21341 534 21375
rect 500 21273 534 21307
rect 500 21205 534 21239
rect 500 21137 534 21171
rect 500 21069 534 21103
rect 500 21001 534 21035
rect 500 20933 534 20967
rect 500 20865 534 20899
rect 500 20797 534 20831
rect 500 20729 534 20763
rect 500 20661 534 20695
rect 758 21545 792 21579
rect 758 21477 792 21511
rect 758 21409 792 21443
rect 758 21341 792 21375
rect 758 21273 792 21307
rect 758 21205 792 21239
rect 758 21137 792 21171
rect 758 21069 792 21103
rect 758 21001 792 21035
rect 758 20933 792 20967
rect 758 20865 792 20899
rect 758 20797 792 20831
rect 758 20729 792 20763
rect 758 20661 792 20695
rect 1016 21545 1050 21579
rect 1016 21477 1050 21511
rect 1016 21409 1050 21443
rect 1016 21341 1050 21375
rect 1016 21273 1050 21307
rect 1016 21205 1050 21239
rect 1016 21137 1050 21171
rect 1016 21069 1050 21103
rect 1016 21001 1050 21035
rect 1016 20933 1050 20967
rect 1016 20865 1050 20899
rect 1016 20797 1050 20831
rect 1016 20729 1050 20763
rect 1016 20661 1050 20695
rect 1274 21545 1308 21579
rect 1274 21477 1308 21511
rect 1274 21409 1308 21443
rect 1274 21341 1308 21375
rect 1274 21273 1308 21307
rect 1274 21205 1308 21239
rect 1274 21137 1308 21171
rect 1274 21069 1308 21103
rect 1274 21001 1308 21035
rect 1274 20933 1308 20967
rect 1274 20865 1308 20899
rect 1274 20797 1308 20831
rect 1274 20729 1308 20763
rect 1274 20661 1308 20695
rect 1532 21545 1566 21579
rect 1532 21477 1566 21511
rect 1532 21409 1566 21443
rect 1532 21341 1566 21375
rect 1532 21273 1566 21307
rect 1532 21205 1566 21239
rect 1532 21137 1566 21171
rect 1532 21069 1566 21103
rect 1532 21001 1566 21035
rect 1532 20933 1566 20967
rect 1532 20865 1566 20899
rect 1532 20797 1566 20831
rect 1532 20729 1566 20763
rect 1532 20661 1566 20695
rect 1790 21545 1824 21579
rect 1790 21477 1824 21511
rect 1790 21409 1824 21443
rect 1790 21341 1824 21375
rect 1790 21273 1824 21307
rect 1790 21205 1824 21239
rect 1790 21137 1824 21171
rect 1790 21069 1824 21103
rect 1790 21001 1824 21035
rect 1790 20933 1824 20967
rect 1790 20865 1824 20899
rect 1790 20797 1824 20831
rect 1790 20729 1824 20763
rect 1790 20661 1824 20695
rect -818 18018 -592 18052
rect -350 18018 -124 18052
rect 118 18018 344 18052
rect 586 18018 812 18052
rect -818 17760 -592 17794
rect -350 17760 -124 17794
rect 118 17760 344 17794
rect 586 17760 812 17794
rect -598 17393 -122 17427
rect 120 17393 596 17427
rect -598 17235 -122 17269
rect 120 17235 596 17269
rect -3533 16868 -2557 16902
rect -2315 16868 -1339 16902
rect -1097 16868 -121 16902
rect 121 16868 1097 16902
rect 1339 16868 2315 16902
rect 2557 16868 3533 16902
rect -3533 16610 -2557 16644
rect -2315 16610 -1339 16644
rect -1097 16610 -121 16644
rect 121 16610 1097 16644
rect 1339 16610 2315 16644
rect 2557 16610 3533 16644
<< pdiffc >>
rect -3172 30884 -3138 30918
rect -3172 30816 -3138 30850
rect -3172 30748 -3138 30782
rect -3172 30680 -3138 30714
rect -3172 30612 -3138 30646
rect -3172 30544 -3138 30578
rect -3172 30476 -3138 30510
rect -3172 30408 -3138 30442
rect -3172 30340 -3138 30374
rect -3172 30272 -3138 30306
rect -3172 30204 -3138 30238
rect -3172 30136 -3138 30170
rect -3172 30068 -3138 30102
rect -3172 30000 -3138 30034
rect -3014 30884 -2980 30918
rect -3014 30816 -2980 30850
rect -3014 30748 -2980 30782
rect -3014 30680 -2980 30714
rect -3014 30612 -2980 30646
rect -3014 30544 -2980 30578
rect -3014 30476 -2980 30510
rect -3014 30408 -2980 30442
rect -3014 30340 -2980 30374
rect -3014 30272 -2980 30306
rect -3014 30204 -2980 30238
rect -3014 30136 -2980 30170
rect -3014 30068 -2980 30102
rect -3014 30000 -2980 30034
rect -2856 30884 -2822 30918
rect -2856 30816 -2822 30850
rect -2856 30748 -2822 30782
rect -2856 30680 -2822 30714
rect -2856 30612 -2822 30646
rect -2856 30544 -2822 30578
rect -2856 30476 -2822 30510
rect -2856 30408 -2822 30442
rect -2856 30340 -2822 30374
rect -2856 30272 -2822 30306
rect -2856 30204 -2822 30238
rect -2856 30136 -2822 30170
rect -2856 30068 -2822 30102
rect -2856 30000 -2822 30034
rect -2698 30884 -2664 30918
rect -2698 30816 -2664 30850
rect -2698 30748 -2664 30782
rect -2698 30680 -2664 30714
rect -2698 30612 -2664 30646
rect -2698 30544 -2664 30578
rect -2698 30476 -2664 30510
rect -2698 30408 -2664 30442
rect -2698 30340 -2664 30374
rect -2698 30272 -2664 30306
rect -2698 30204 -2664 30238
rect -2698 30136 -2664 30170
rect -2698 30068 -2664 30102
rect -2698 30000 -2664 30034
rect -2540 30884 -2506 30918
rect -2540 30816 -2506 30850
rect -2540 30748 -2506 30782
rect -2540 30680 -2506 30714
rect -2540 30612 -2506 30646
rect -2540 30544 -2506 30578
rect -2540 30476 -2506 30510
rect -2540 30408 -2506 30442
rect -2540 30340 -2506 30374
rect -2540 30272 -2506 30306
rect -2540 30204 -2506 30238
rect -2540 30136 -2506 30170
rect -2540 30068 -2506 30102
rect -2540 30000 -2506 30034
rect -2382 30884 -2348 30918
rect -2382 30816 -2348 30850
rect -2382 30748 -2348 30782
rect -2382 30680 -2348 30714
rect -2382 30612 -2348 30646
rect -2382 30544 -2348 30578
rect -2382 30476 -2348 30510
rect -2382 30408 -2348 30442
rect -2382 30340 -2348 30374
rect -2382 30272 -2348 30306
rect -2382 30204 -2348 30238
rect -2382 30136 -2348 30170
rect -2382 30068 -2348 30102
rect -2382 30000 -2348 30034
rect -2224 30884 -2190 30918
rect -2224 30816 -2190 30850
rect -2224 30748 -2190 30782
rect -2224 30680 -2190 30714
rect -2224 30612 -2190 30646
rect -2224 30544 -2190 30578
rect -2224 30476 -2190 30510
rect -2224 30408 -2190 30442
rect -2224 30340 -2190 30374
rect -2224 30272 -2190 30306
rect -2224 30204 -2190 30238
rect -2224 30136 -2190 30170
rect -2224 30068 -2190 30102
rect -2224 30000 -2190 30034
rect -2066 30884 -2032 30918
rect -2066 30816 -2032 30850
rect -2066 30748 -2032 30782
rect -2066 30680 -2032 30714
rect -2066 30612 -2032 30646
rect -2066 30544 -2032 30578
rect -2066 30476 -2032 30510
rect -2066 30408 -2032 30442
rect -2066 30340 -2032 30374
rect -2066 30272 -2032 30306
rect -2066 30204 -2032 30238
rect -2066 30136 -2032 30170
rect -2066 30068 -2032 30102
rect -2066 30000 -2032 30034
rect -1908 30884 -1874 30918
rect -1908 30816 -1874 30850
rect -1908 30748 -1874 30782
rect -1908 30680 -1874 30714
rect -1908 30612 -1874 30646
rect -1908 30544 -1874 30578
rect -1908 30476 -1874 30510
rect -1908 30408 -1874 30442
rect -1908 30340 -1874 30374
rect -1908 30272 -1874 30306
rect -1908 30204 -1874 30238
rect -1908 30136 -1874 30170
rect -1908 30068 -1874 30102
rect -1908 30000 -1874 30034
rect -1750 30884 -1716 30918
rect -1750 30816 -1716 30850
rect -1750 30748 -1716 30782
rect -1750 30680 -1716 30714
rect -1750 30612 -1716 30646
rect -1750 30544 -1716 30578
rect -1750 30476 -1716 30510
rect -1750 30408 -1716 30442
rect -1750 30340 -1716 30374
rect -1750 30272 -1716 30306
rect -1750 30204 -1716 30238
rect -1750 30136 -1716 30170
rect -1750 30068 -1716 30102
rect -1750 30000 -1716 30034
rect -1592 30884 -1558 30918
rect -1592 30816 -1558 30850
rect -1592 30748 -1558 30782
rect -1592 30680 -1558 30714
rect -1592 30612 -1558 30646
rect -1592 30544 -1558 30578
rect -1592 30476 -1558 30510
rect -1592 30408 -1558 30442
rect -1592 30340 -1558 30374
rect -1592 30272 -1558 30306
rect -1592 30204 -1558 30238
rect -1592 30136 -1558 30170
rect -1592 30068 -1558 30102
rect -1592 30000 -1558 30034
rect -1434 30884 -1400 30918
rect -1434 30816 -1400 30850
rect -1434 30748 -1400 30782
rect -1434 30680 -1400 30714
rect -1434 30612 -1400 30646
rect -1434 30544 -1400 30578
rect -1434 30476 -1400 30510
rect -1434 30408 -1400 30442
rect -1434 30340 -1400 30374
rect -1434 30272 -1400 30306
rect -1434 30204 -1400 30238
rect -1434 30136 -1400 30170
rect -1434 30068 -1400 30102
rect -1434 30000 -1400 30034
rect -1276 30884 -1242 30918
rect -1276 30816 -1242 30850
rect -1276 30748 -1242 30782
rect -1276 30680 -1242 30714
rect -1276 30612 -1242 30646
rect -1276 30544 -1242 30578
rect -1276 30476 -1242 30510
rect -1276 30408 -1242 30442
rect -1276 30340 -1242 30374
rect -1276 30272 -1242 30306
rect -1276 30204 -1242 30238
rect -1276 30136 -1242 30170
rect -1276 30068 -1242 30102
rect -1276 30000 -1242 30034
rect -1118 30884 -1084 30918
rect -1118 30816 -1084 30850
rect -1118 30748 -1084 30782
rect -1118 30680 -1084 30714
rect -1118 30612 -1084 30646
rect -1118 30544 -1084 30578
rect -1118 30476 -1084 30510
rect -1118 30408 -1084 30442
rect -1118 30340 -1084 30374
rect -1118 30272 -1084 30306
rect -1118 30204 -1084 30238
rect -1118 30136 -1084 30170
rect -1118 30068 -1084 30102
rect -1118 30000 -1084 30034
rect -960 30884 -926 30918
rect -960 30816 -926 30850
rect -960 30748 -926 30782
rect -960 30680 -926 30714
rect -960 30612 -926 30646
rect -960 30544 -926 30578
rect -960 30476 -926 30510
rect -960 30408 -926 30442
rect -960 30340 -926 30374
rect -960 30272 -926 30306
rect -960 30204 -926 30238
rect -960 30136 -926 30170
rect -960 30068 -926 30102
rect -960 30000 -926 30034
rect -802 30884 -768 30918
rect -802 30816 -768 30850
rect -802 30748 -768 30782
rect -802 30680 -768 30714
rect -802 30612 -768 30646
rect -802 30544 -768 30578
rect -802 30476 -768 30510
rect -802 30408 -768 30442
rect -802 30340 -768 30374
rect -802 30272 -768 30306
rect -802 30204 -768 30238
rect -802 30136 -768 30170
rect -802 30068 -768 30102
rect -802 30000 -768 30034
rect -644 30884 -610 30918
rect -644 30816 -610 30850
rect -644 30748 -610 30782
rect -644 30680 -610 30714
rect -644 30612 -610 30646
rect -644 30544 -610 30578
rect -644 30476 -610 30510
rect -644 30408 -610 30442
rect -644 30340 -610 30374
rect -644 30272 -610 30306
rect -644 30204 -610 30238
rect -644 30136 -610 30170
rect -644 30068 -610 30102
rect -644 30000 -610 30034
rect -486 30884 -452 30918
rect -486 30816 -452 30850
rect -486 30748 -452 30782
rect -486 30680 -452 30714
rect -486 30612 -452 30646
rect -486 30544 -452 30578
rect -486 30476 -452 30510
rect -486 30408 -452 30442
rect -486 30340 -452 30374
rect -486 30272 -452 30306
rect -486 30204 -452 30238
rect -486 30136 -452 30170
rect -486 30068 -452 30102
rect -486 30000 -452 30034
rect -328 30884 -294 30918
rect -328 30816 -294 30850
rect -328 30748 -294 30782
rect -328 30680 -294 30714
rect -328 30612 -294 30646
rect -328 30544 -294 30578
rect -328 30476 -294 30510
rect -328 30408 -294 30442
rect -328 30340 -294 30374
rect -328 30272 -294 30306
rect -328 30204 -294 30238
rect -328 30136 -294 30170
rect -328 30068 -294 30102
rect -328 30000 -294 30034
rect -170 30884 -136 30918
rect -170 30816 -136 30850
rect -170 30748 -136 30782
rect -170 30680 -136 30714
rect -170 30612 -136 30646
rect -170 30544 -136 30578
rect -170 30476 -136 30510
rect -170 30408 -136 30442
rect -170 30340 -136 30374
rect -170 30272 -136 30306
rect -170 30204 -136 30238
rect -170 30136 -136 30170
rect -170 30068 -136 30102
rect -170 30000 -136 30034
rect -12 30884 22 30918
rect -12 30816 22 30850
rect -12 30748 22 30782
rect -12 30680 22 30714
rect -12 30612 22 30646
rect -12 30544 22 30578
rect -12 30476 22 30510
rect -12 30408 22 30442
rect -12 30340 22 30374
rect -12 30272 22 30306
rect -12 30204 22 30238
rect -12 30136 22 30170
rect -12 30068 22 30102
rect -12 30000 22 30034
rect 146 30884 180 30918
rect 146 30816 180 30850
rect 146 30748 180 30782
rect 146 30680 180 30714
rect 146 30612 180 30646
rect 146 30544 180 30578
rect 146 30476 180 30510
rect 146 30408 180 30442
rect 146 30340 180 30374
rect 146 30272 180 30306
rect 146 30204 180 30238
rect 146 30136 180 30170
rect 146 30068 180 30102
rect 146 30000 180 30034
rect 304 30884 338 30918
rect 304 30816 338 30850
rect 304 30748 338 30782
rect 304 30680 338 30714
rect 304 30612 338 30646
rect 304 30544 338 30578
rect 304 30476 338 30510
rect 304 30408 338 30442
rect 304 30340 338 30374
rect 304 30272 338 30306
rect 304 30204 338 30238
rect 304 30136 338 30170
rect 304 30068 338 30102
rect 304 30000 338 30034
rect 462 30884 496 30918
rect 462 30816 496 30850
rect 462 30748 496 30782
rect 462 30680 496 30714
rect 462 30612 496 30646
rect 462 30544 496 30578
rect 462 30476 496 30510
rect 462 30408 496 30442
rect 462 30340 496 30374
rect 462 30272 496 30306
rect 462 30204 496 30238
rect 462 30136 496 30170
rect 462 30068 496 30102
rect 462 30000 496 30034
rect 620 30884 654 30918
rect 620 30816 654 30850
rect 620 30748 654 30782
rect 620 30680 654 30714
rect 620 30612 654 30646
rect 620 30544 654 30578
rect 620 30476 654 30510
rect 620 30408 654 30442
rect 620 30340 654 30374
rect 620 30272 654 30306
rect 620 30204 654 30238
rect 620 30136 654 30170
rect 620 30068 654 30102
rect 620 30000 654 30034
rect 778 30884 812 30918
rect 778 30816 812 30850
rect 778 30748 812 30782
rect 778 30680 812 30714
rect 778 30612 812 30646
rect 778 30544 812 30578
rect 778 30476 812 30510
rect 778 30408 812 30442
rect 778 30340 812 30374
rect 778 30272 812 30306
rect 778 30204 812 30238
rect 778 30136 812 30170
rect 778 30068 812 30102
rect 778 30000 812 30034
rect 936 30884 970 30918
rect 936 30816 970 30850
rect 936 30748 970 30782
rect 936 30680 970 30714
rect 936 30612 970 30646
rect 936 30544 970 30578
rect 936 30476 970 30510
rect 936 30408 970 30442
rect 936 30340 970 30374
rect 936 30272 970 30306
rect 936 30204 970 30238
rect 936 30136 970 30170
rect 936 30068 970 30102
rect 936 30000 970 30034
rect 1094 30884 1128 30918
rect 1094 30816 1128 30850
rect 1094 30748 1128 30782
rect 1094 30680 1128 30714
rect 1094 30612 1128 30646
rect 1094 30544 1128 30578
rect 1094 30476 1128 30510
rect 1094 30408 1128 30442
rect 1094 30340 1128 30374
rect 1094 30272 1128 30306
rect 1094 30204 1128 30238
rect 1094 30136 1128 30170
rect 1094 30068 1128 30102
rect 1094 30000 1128 30034
rect 1252 30884 1286 30918
rect 1252 30816 1286 30850
rect 1252 30748 1286 30782
rect 1252 30680 1286 30714
rect 1252 30612 1286 30646
rect 1252 30544 1286 30578
rect 1252 30476 1286 30510
rect 1252 30408 1286 30442
rect 1252 30340 1286 30374
rect 1252 30272 1286 30306
rect 1252 30204 1286 30238
rect 1252 30136 1286 30170
rect 1252 30068 1286 30102
rect 1252 30000 1286 30034
rect 1410 30884 1444 30918
rect 1410 30816 1444 30850
rect 1410 30748 1444 30782
rect 1410 30680 1444 30714
rect 1410 30612 1444 30646
rect 1410 30544 1444 30578
rect 1410 30476 1444 30510
rect 1410 30408 1444 30442
rect 1410 30340 1444 30374
rect 1410 30272 1444 30306
rect 1410 30204 1444 30238
rect 1410 30136 1444 30170
rect 1410 30068 1444 30102
rect 1410 30000 1444 30034
rect 1568 30884 1602 30918
rect 1568 30816 1602 30850
rect 1568 30748 1602 30782
rect 1568 30680 1602 30714
rect 1568 30612 1602 30646
rect 1568 30544 1602 30578
rect 1568 30476 1602 30510
rect 1568 30408 1602 30442
rect 1568 30340 1602 30374
rect 1568 30272 1602 30306
rect 1568 30204 1602 30238
rect 1568 30136 1602 30170
rect 1568 30068 1602 30102
rect 1568 30000 1602 30034
rect 1726 30884 1760 30918
rect 1726 30816 1760 30850
rect 1726 30748 1760 30782
rect 1726 30680 1760 30714
rect 1726 30612 1760 30646
rect 1726 30544 1760 30578
rect 1726 30476 1760 30510
rect 1726 30408 1760 30442
rect 1726 30340 1760 30374
rect 1726 30272 1760 30306
rect 1726 30204 1760 30238
rect 1726 30136 1760 30170
rect 1726 30068 1760 30102
rect 1726 30000 1760 30034
rect 1884 30884 1918 30918
rect 1884 30816 1918 30850
rect 1884 30748 1918 30782
rect 1884 30680 1918 30714
rect 1884 30612 1918 30646
rect 1884 30544 1918 30578
rect 1884 30476 1918 30510
rect 1884 30408 1918 30442
rect 1884 30340 1918 30374
rect 1884 30272 1918 30306
rect 1884 30204 1918 30238
rect 1884 30136 1918 30170
rect 1884 30068 1918 30102
rect 1884 30000 1918 30034
rect 2042 30884 2076 30918
rect 2042 30816 2076 30850
rect 2042 30748 2076 30782
rect 2042 30680 2076 30714
rect 2042 30612 2076 30646
rect 2042 30544 2076 30578
rect 2042 30476 2076 30510
rect 2042 30408 2076 30442
rect 2042 30340 2076 30374
rect 2042 30272 2076 30306
rect 2042 30204 2076 30238
rect 2042 30136 2076 30170
rect 2042 30068 2076 30102
rect 2042 30000 2076 30034
rect 2200 30884 2234 30918
rect 2200 30816 2234 30850
rect 2200 30748 2234 30782
rect 2200 30680 2234 30714
rect 2200 30612 2234 30646
rect 2200 30544 2234 30578
rect 2200 30476 2234 30510
rect 2200 30408 2234 30442
rect 2200 30340 2234 30374
rect 2200 30272 2234 30306
rect 2200 30204 2234 30238
rect 2200 30136 2234 30170
rect 2200 30068 2234 30102
rect 2200 30000 2234 30034
rect 2358 30884 2392 30918
rect 2358 30816 2392 30850
rect 2358 30748 2392 30782
rect 2358 30680 2392 30714
rect 2358 30612 2392 30646
rect 2358 30544 2392 30578
rect 2358 30476 2392 30510
rect 2358 30408 2392 30442
rect 2358 30340 2392 30374
rect 2358 30272 2392 30306
rect 2358 30204 2392 30238
rect 2358 30136 2392 30170
rect 2358 30068 2392 30102
rect 2358 30000 2392 30034
rect 2516 30884 2550 30918
rect 2516 30816 2550 30850
rect 2516 30748 2550 30782
rect 2516 30680 2550 30714
rect 2516 30612 2550 30646
rect 2516 30544 2550 30578
rect 2516 30476 2550 30510
rect 2516 30408 2550 30442
rect 2516 30340 2550 30374
rect 2516 30272 2550 30306
rect 2516 30204 2550 30238
rect 2516 30136 2550 30170
rect 2516 30068 2550 30102
rect 2516 30000 2550 30034
rect 2674 30884 2708 30918
rect 2674 30816 2708 30850
rect 2674 30748 2708 30782
rect 2674 30680 2708 30714
rect 2674 30612 2708 30646
rect 2674 30544 2708 30578
rect 2674 30476 2708 30510
rect 2674 30408 2708 30442
rect 2674 30340 2708 30374
rect 2674 30272 2708 30306
rect 2674 30204 2708 30238
rect 2674 30136 2708 30170
rect 2674 30068 2708 30102
rect 2674 30000 2708 30034
rect 2832 30884 2866 30918
rect 2832 30816 2866 30850
rect 2832 30748 2866 30782
rect 2832 30680 2866 30714
rect 2832 30612 2866 30646
rect 2832 30544 2866 30578
rect 2832 30476 2866 30510
rect 2832 30408 2866 30442
rect 2832 30340 2866 30374
rect 2832 30272 2866 30306
rect 2832 30204 2866 30238
rect 2832 30136 2866 30170
rect 2832 30068 2866 30102
rect 2832 30000 2866 30034
rect 2990 30884 3024 30918
rect 2990 30816 3024 30850
rect 2990 30748 3024 30782
rect 2990 30680 3024 30714
rect 2990 30612 3024 30646
rect 2990 30544 3024 30578
rect 2990 30476 3024 30510
rect 2990 30408 3024 30442
rect 2990 30340 3024 30374
rect 2990 30272 3024 30306
rect 2990 30204 3024 30238
rect 2990 30136 3024 30170
rect 2990 30068 3024 30102
rect 2990 30000 3024 30034
rect 3148 30884 3182 30918
rect 3148 30816 3182 30850
rect 3148 30748 3182 30782
rect 3148 30680 3182 30714
rect 3148 30612 3182 30646
rect 3148 30544 3182 30578
rect 3148 30476 3182 30510
rect 3148 30408 3182 30442
rect 3148 30340 3182 30374
rect 3148 30272 3182 30306
rect 3148 30204 3182 30238
rect 3148 30136 3182 30170
rect 3148 30068 3182 30102
rect 3148 30000 3182 30034
rect -1672 29214 -1638 29248
rect -1672 29146 -1638 29180
rect -1672 29078 -1638 29112
rect -1672 29010 -1638 29044
rect -1672 28942 -1638 28976
rect -1672 28874 -1638 28908
rect -1672 28806 -1638 28840
rect -1672 28738 -1638 28772
rect -1672 28670 -1638 28704
rect -1672 28602 -1638 28636
rect -1672 28534 -1638 28568
rect -1672 28466 -1638 28500
rect -1672 28398 -1638 28432
rect -1672 28330 -1638 28364
rect -1514 29214 -1480 29248
rect -1514 29146 -1480 29180
rect -1514 29078 -1480 29112
rect -1514 29010 -1480 29044
rect -1514 28942 -1480 28976
rect -1514 28874 -1480 28908
rect -1514 28806 -1480 28840
rect -1514 28738 -1480 28772
rect -1514 28670 -1480 28704
rect -1514 28602 -1480 28636
rect -1514 28534 -1480 28568
rect -1514 28466 -1480 28500
rect -1514 28398 -1480 28432
rect -1514 28330 -1480 28364
rect -1356 29214 -1322 29248
rect -1356 29146 -1322 29180
rect -1356 29078 -1322 29112
rect -1356 29010 -1322 29044
rect -1356 28942 -1322 28976
rect -1356 28874 -1322 28908
rect -1356 28806 -1322 28840
rect -1356 28738 -1322 28772
rect -1356 28670 -1322 28704
rect -1356 28602 -1322 28636
rect -1356 28534 -1322 28568
rect -1356 28466 -1322 28500
rect -1356 28398 -1322 28432
rect -1356 28330 -1322 28364
rect -1198 29214 -1164 29248
rect -1198 29146 -1164 29180
rect -1198 29078 -1164 29112
rect -1198 29010 -1164 29044
rect -1198 28942 -1164 28976
rect -1198 28874 -1164 28908
rect -1198 28806 -1164 28840
rect -1198 28738 -1164 28772
rect -1198 28670 -1164 28704
rect -1198 28602 -1164 28636
rect -1198 28534 -1164 28568
rect -1198 28466 -1164 28500
rect -1198 28398 -1164 28432
rect -1198 28330 -1164 28364
rect -1040 29214 -1006 29248
rect -1040 29146 -1006 29180
rect -1040 29078 -1006 29112
rect -1040 29010 -1006 29044
rect -1040 28942 -1006 28976
rect -1040 28874 -1006 28908
rect -1040 28806 -1006 28840
rect -1040 28738 -1006 28772
rect -1040 28670 -1006 28704
rect -1040 28602 -1006 28636
rect -1040 28534 -1006 28568
rect -1040 28466 -1006 28500
rect -1040 28398 -1006 28432
rect -1040 28330 -1006 28364
rect -882 29214 -848 29248
rect -882 29146 -848 29180
rect -882 29078 -848 29112
rect -882 29010 -848 29044
rect -882 28942 -848 28976
rect -882 28874 -848 28908
rect -882 28806 -848 28840
rect -882 28738 -848 28772
rect -882 28670 -848 28704
rect -882 28602 -848 28636
rect -882 28534 -848 28568
rect -882 28466 -848 28500
rect -882 28398 -848 28432
rect -882 28330 -848 28364
rect -724 29214 -690 29248
rect -724 29146 -690 29180
rect -724 29078 -690 29112
rect -724 29010 -690 29044
rect -724 28942 -690 28976
rect -724 28874 -690 28908
rect -724 28806 -690 28840
rect -724 28738 -690 28772
rect -724 28670 -690 28704
rect -724 28602 -690 28636
rect -724 28534 -690 28568
rect -724 28466 -690 28500
rect -724 28398 -690 28432
rect -724 28330 -690 28364
rect -566 29214 -532 29248
rect -566 29146 -532 29180
rect -566 29078 -532 29112
rect -566 29010 -532 29044
rect -566 28942 -532 28976
rect -566 28874 -532 28908
rect -566 28806 -532 28840
rect -566 28738 -532 28772
rect -566 28670 -532 28704
rect -566 28602 -532 28636
rect -566 28534 -532 28568
rect -566 28466 -532 28500
rect -566 28398 -532 28432
rect -566 28330 -532 28364
rect -408 29214 -374 29248
rect -408 29146 -374 29180
rect -408 29078 -374 29112
rect -408 29010 -374 29044
rect -408 28942 -374 28976
rect -408 28874 -374 28908
rect -408 28806 -374 28840
rect -408 28738 -374 28772
rect -408 28670 -374 28704
rect -408 28602 -374 28636
rect -408 28534 -374 28568
rect -408 28466 -374 28500
rect -408 28398 -374 28432
rect -408 28330 -374 28364
rect -250 29214 -216 29248
rect -250 29146 -216 29180
rect -250 29078 -216 29112
rect -250 29010 -216 29044
rect -250 28942 -216 28976
rect -250 28874 -216 28908
rect -250 28806 -216 28840
rect -250 28738 -216 28772
rect -250 28670 -216 28704
rect -250 28602 -216 28636
rect -250 28534 -216 28568
rect -250 28466 -216 28500
rect -250 28398 -216 28432
rect -250 28330 -216 28364
rect -92 29214 -58 29248
rect -92 29146 -58 29180
rect -92 29078 -58 29112
rect -92 29010 -58 29044
rect -92 28942 -58 28976
rect -92 28874 -58 28908
rect -92 28806 -58 28840
rect -92 28738 -58 28772
rect -92 28670 -58 28704
rect -92 28602 -58 28636
rect -92 28534 -58 28568
rect -92 28466 -58 28500
rect -92 28398 -58 28432
rect -92 28330 -58 28364
rect 66 29214 100 29248
rect 66 29146 100 29180
rect 66 29078 100 29112
rect 66 29010 100 29044
rect 66 28942 100 28976
rect 66 28874 100 28908
rect 66 28806 100 28840
rect 66 28738 100 28772
rect 66 28670 100 28704
rect 66 28602 100 28636
rect 66 28534 100 28568
rect 66 28466 100 28500
rect 66 28398 100 28432
rect 66 28330 100 28364
rect 224 29214 258 29248
rect 224 29146 258 29180
rect 224 29078 258 29112
rect 224 29010 258 29044
rect 224 28942 258 28976
rect 224 28874 258 28908
rect 224 28806 258 28840
rect 224 28738 258 28772
rect 224 28670 258 28704
rect 224 28602 258 28636
rect 224 28534 258 28568
rect 224 28466 258 28500
rect 224 28398 258 28432
rect 224 28330 258 28364
rect 382 29214 416 29248
rect 382 29146 416 29180
rect 382 29078 416 29112
rect 382 29010 416 29044
rect 382 28942 416 28976
rect 382 28874 416 28908
rect 382 28806 416 28840
rect 382 28738 416 28772
rect 382 28670 416 28704
rect 382 28602 416 28636
rect 382 28534 416 28568
rect 382 28466 416 28500
rect 382 28398 416 28432
rect 382 28330 416 28364
rect 540 29214 574 29248
rect 540 29146 574 29180
rect 540 29078 574 29112
rect 540 29010 574 29044
rect 540 28942 574 28976
rect 540 28874 574 28908
rect 540 28806 574 28840
rect 540 28738 574 28772
rect 540 28670 574 28704
rect 540 28602 574 28636
rect 540 28534 574 28568
rect 540 28466 574 28500
rect 540 28398 574 28432
rect 540 28330 574 28364
rect 698 29214 732 29248
rect 698 29146 732 29180
rect 698 29078 732 29112
rect 698 29010 732 29044
rect 698 28942 732 28976
rect 698 28874 732 28908
rect 698 28806 732 28840
rect 698 28738 732 28772
rect 698 28670 732 28704
rect 698 28602 732 28636
rect 698 28534 732 28568
rect 698 28466 732 28500
rect 698 28398 732 28432
rect 698 28330 732 28364
rect 856 29214 890 29248
rect 856 29146 890 29180
rect 856 29078 890 29112
rect 856 29010 890 29044
rect 856 28942 890 28976
rect 856 28874 890 28908
rect 856 28806 890 28840
rect 856 28738 890 28772
rect 856 28670 890 28704
rect 856 28602 890 28636
rect 856 28534 890 28568
rect 856 28466 890 28500
rect 856 28398 890 28432
rect 856 28330 890 28364
rect 1014 29214 1048 29248
rect 1014 29146 1048 29180
rect 1014 29078 1048 29112
rect 1014 29010 1048 29044
rect 1014 28942 1048 28976
rect 1014 28874 1048 28908
rect 1014 28806 1048 28840
rect 1014 28738 1048 28772
rect 1014 28670 1048 28704
rect 1014 28602 1048 28636
rect 1014 28534 1048 28568
rect 1014 28466 1048 28500
rect 1014 28398 1048 28432
rect 1014 28330 1048 28364
rect 1172 29214 1206 29248
rect 1172 29146 1206 29180
rect 1172 29078 1206 29112
rect 1172 29010 1206 29044
rect 1172 28942 1206 28976
rect 1172 28874 1206 28908
rect 1172 28806 1206 28840
rect 1172 28738 1206 28772
rect 1172 28670 1206 28704
rect 1172 28602 1206 28636
rect 1172 28534 1206 28568
rect 1172 28466 1206 28500
rect 1172 28398 1206 28432
rect 1172 28330 1206 28364
rect 1330 29214 1364 29248
rect 1330 29146 1364 29180
rect 1330 29078 1364 29112
rect 1330 29010 1364 29044
rect 1330 28942 1364 28976
rect 1330 28874 1364 28908
rect 1330 28806 1364 28840
rect 1330 28738 1364 28772
rect 1330 28670 1364 28704
rect 1330 28602 1364 28636
rect 1330 28534 1364 28568
rect 1330 28466 1364 28500
rect 1330 28398 1364 28432
rect 1330 28330 1364 28364
rect 1488 29214 1522 29248
rect 1488 29146 1522 29180
rect 1488 29078 1522 29112
rect 1488 29010 1522 29044
rect 1488 28942 1522 28976
rect 1488 28874 1522 28908
rect 1488 28806 1522 28840
rect 1488 28738 1522 28772
rect 1488 28670 1522 28704
rect 1488 28602 1522 28636
rect 1488 28534 1522 28568
rect 1488 28466 1522 28500
rect 1488 28398 1522 28432
rect 1488 28330 1522 28364
rect 1646 29214 1680 29248
rect 1646 29146 1680 29180
rect 1646 29078 1680 29112
rect 1646 29010 1680 29044
rect 1646 28942 1680 28976
rect 1646 28874 1680 28908
rect 1646 28806 1680 28840
rect 1646 28738 1680 28772
rect 1646 28670 1680 28704
rect 1646 28602 1680 28636
rect 1646 28534 1680 28568
rect 1646 28466 1680 28500
rect 1646 28398 1680 28432
rect 1646 28330 1680 28364
rect -1672 27674 -1638 27708
rect -1672 27606 -1638 27640
rect -1672 27538 -1638 27572
rect -1672 27470 -1638 27504
rect -1672 27402 -1638 27436
rect -1672 27334 -1638 27368
rect -1672 27266 -1638 27300
rect -1672 27198 -1638 27232
rect -1672 27130 -1638 27164
rect -1672 27062 -1638 27096
rect -1672 26994 -1638 27028
rect -1672 26926 -1638 26960
rect -1672 26858 -1638 26892
rect -1672 26790 -1638 26824
rect -1514 27674 -1480 27708
rect -1514 27606 -1480 27640
rect -1514 27538 -1480 27572
rect -1514 27470 -1480 27504
rect -1514 27402 -1480 27436
rect -1514 27334 -1480 27368
rect -1514 27266 -1480 27300
rect -1514 27198 -1480 27232
rect -1514 27130 -1480 27164
rect -1514 27062 -1480 27096
rect -1514 26994 -1480 27028
rect -1514 26926 -1480 26960
rect -1514 26858 -1480 26892
rect -1514 26790 -1480 26824
rect -1356 27674 -1322 27708
rect -1356 27606 -1322 27640
rect -1356 27538 -1322 27572
rect -1356 27470 -1322 27504
rect -1356 27402 -1322 27436
rect -1356 27334 -1322 27368
rect -1356 27266 -1322 27300
rect -1356 27198 -1322 27232
rect -1356 27130 -1322 27164
rect -1356 27062 -1322 27096
rect -1356 26994 -1322 27028
rect -1356 26926 -1322 26960
rect -1356 26858 -1322 26892
rect -1356 26790 -1322 26824
rect -1198 27674 -1164 27708
rect -1198 27606 -1164 27640
rect -1198 27538 -1164 27572
rect -1198 27470 -1164 27504
rect -1198 27402 -1164 27436
rect -1198 27334 -1164 27368
rect -1198 27266 -1164 27300
rect -1198 27198 -1164 27232
rect -1198 27130 -1164 27164
rect -1198 27062 -1164 27096
rect -1198 26994 -1164 27028
rect -1198 26926 -1164 26960
rect -1198 26858 -1164 26892
rect -1198 26790 -1164 26824
rect -1040 27674 -1006 27708
rect -1040 27606 -1006 27640
rect -1040 27538 -1006 27572
rect -1040 27470 -1006 27504
rect -1040 27402 -1006 27436
rect -1040 27334 -1006 27368
rect -1040 27266 -1006 27300
rect -1040 27198 -1006 27232
rect -1040 27130 -1006 27164
rect -1040 27062 -1006 27096
rect -1040 26994 -1006 27028
rect -1040 26926 -1006 26960
rect -1040 26858 -1006 26892
rect -1040 26790 -1006 26824
rect -882 27674 -848 27708
rect -882 27606 -848 27640
rect -882 27538 -848 27572
rect -882 27470 -848 27504
rect -882 27402 -848 27436
rect -882 27334 -848 27368
rect -882 27266 -848 27300
rect -882 27198 -848 27232
rect -882 27130 -848 27164
rect -882 27062 -848 27096
rect -882 26994 -848 27028
rect -882 26926 -848 26960
rect -882 26858 -848 26892
rect -882 26790 -848 26824
rect -724 27674 -690 27708
rect -724 27606 -690 27640
rect -724 27538 -690 27572
rect -724 27470 -690 27504
rect -724 27402 -690 27436
rect -724 27334 -690 27368
rect -724 27266 -690 27300
rect -724 27198 -690 27232
rect -724 27130 -690 27164
rect -724 27062 -690 27096
rect -724 26994 -690 27028
rect -724 26926 -690 26960
rect -724 26858 -690 26892
rect -724 26790 -690 26824
rect -566 27674 -532 27708
rect -566 27606 -532 27640
rect -566 27538 -532 27572
rect -566 27470 -532 27504
rect -566 27402 -532 27436
rect -566 27334 -532 27368
rect -566 27266 -532 27300
rect -566 27198 -532 27232
rect -566 27130 -532 27164
rect -566 27062 -532 27096
rect -566 26994 -532 27028
rect -566 26926 -532 26960
rect -566 26858 -532 26892
rect -566 26790 -532 26824
rect -408 27674 -374 27708
rect -408 27606 -374 27640
rect -408 27538 -374 27572
rect -408 27470 -374 27504
rect -408 27402 -374 27436
rect -408 27334 -374 27368
rect -408 27266 -374 27300
rect -408 27198 -374 27232
rect -408 27130 -374 27164
rect -408 27062 -374 27096
rect -408 26994 -374 27028
rect -408 26926 -374 26960
rect -408 26858 -374 26892
rect -408 26790 -374 26824
rect -250 27674 -216 27708
rect -250 27606 -216 27640
rect -250 27538 -216 27572
rect -250 27470 -216 27504
rect -250 27402 -216 27436
rect -250 27334 -216 27368
rect -250 27266 -216 27300
rect -250 27198 -216 27232
rect -250 27130 -216 27164
rect -250 27062 -216 27096
rect -250 26994 -216 27028
rect -250 26926 -216 26960
rect -250 26858 -216 26892
rect -250 26790 -216 26824
rect -92 27674 -58 27708
rect -92 27606 -58 27640
rect -92 27538 -58 27572
rect -92 27470 -58 27504
rect -92 27402 -58 27436
rect -92 27334 -58 27368
rect -92 27266 -58 27300
rect -92 27198 -58 27232
rect -92 27130 -58 27164
rect -92 27062 -58 27096
rect -92 26994 -58 27028
rect -92 26926 -58 26960
rect -92 26858 -58 26892
rect -92 26790 -58 26824
rect 66 27674 100 27708
rect 66 27606 100 27640
rect 66 27538 100 27572
rect 66 27470 100 27504
rect 66 27402 100 27436
rect 66 27334 100 27368
rect 66 27266 100 27300
rect 66 27198 100 27232
rect 66 27130 100 27164
rect 66 27062 100 27096
rect 66 26994 100 27028
rect 66 26926 100 26960
rect 66 26858 100 26892
rect 66 26790 100 26824
rect 224 27674 258 27708
rect 224 27606 258 27640
rect 224 27538 258 27572
rect 224 27470 258 27504
rect 224 27402 258 27436
rect 224 27334 258 27368
rect 224 27266 258 27300
rect 224 27198 258 27232
rect 224 27130 258 27164
rect 224 27062 258 27096
rect 224 26994 258 27028
rect 224 26926 258 26960
rect 224 26858 258 26892
rect 224 26790 258 26824
rect 382 27674 416 27708
rect 382 27606 416 27640
rect 382 27538 416 27572
rect 382 27470 416 27504
rect 382 27402 416 27436
rect 382 27334 416 27368
rect 382 27266 416 27300
rect 382 27198 416 27232
rect 382 27130 416 27164
rect 382 27062 416 27096
rect 382 26994 416 27028
rect 382 26926 416 26960
rect 382 26858 416 26892
rect 382 26790 416 26824
rect 540 27674 574 27708
rect 540 27606 574 27640
rect 540 27538 574 27572
rect 540 27470 574 27504
rect 540 27402 574 27436
rect 540 27334 574 27368
rect 540 27266 574 27300
rect 540 27198 574 27232
rect 540 27130 574 27164
rect 540 27062 574 27096
rect 540 26994 574 27028
rect 540 26926 574 26960
rect 540 26858 574 26892
rect 540 26790 574 26824
rect 698 27674 732 27708
rect 698 27606 732 27640
rect 698 27538 732 27572
rect 698 27470 732 27504
rect 698 27402 732 27436
rect 698 27334 732 27368
rect 698 27266 732 27300
rect 698 27198 732 27232
rect 698 27130 732 27164
rect 698 27062 732 27096
rect 698 26994 732 27028
rect 698 26926 732 26960
rect 698 26858 732 26892
rect 698 26790 732 26824
rect 856 27674 890 27708
rect 856 27606 890 27640
rect 856 27538 890 27572
rect 856 27470 890 27504
rect 856 27402 890 27436
rect 856 27334 890 27368
rect 856 27266 890 27300
rect 856 27198 890 27232
rect 856 27130 890 27164
rect 856 27062 890 27096
rect 856 26994 890 27028
rect 856 26926 890 26960
rect 856 26858 890 26892
rect 856 26790 890 26824
rect 1014 27674 1048 27708
rect 1014 27606 1048 27640
rect 1014 27538 1048 27572
rect 1014 27470 1048 27504
rect 1014 27402 1048 27436
rect 1014 27334 1048 27368
rect 1014 27266 1048 27300
rect 1014 27198 1048 27232
rect 1014 27130 1048 27164
rect 1014 27062 1048 27096
rect 1014 26994 1048 27028
rect 1014 26926 1048 26960
rect 1014 26858 1048 26892
rect 1014 26790 1048 26824
rect 1172 27674 1206 27708
rect 1172 27606 1206 27640
rect 1172 27538 1206 27572
rect 1172 27470 1206 27504
rect 1172 27402 1206 27436
rect 1172 27334 1206 27368
rect 1172 27266 1206 27300
rect 1172 27198 1206 27232
rect 1172 27130 1206 27164
rect 1172 27062 1206 27096
rect 1172 26994 1206 27028
rect 1172 26926 1206 26960
rect 1172 26858 1206 26892
rect 1172 26790 1206 26824
rect 1330 27674 1364 27708
rect 1330 27606 1364 27640
rect 1330 27538 1364 27572
rect 1330 27470 1364 27504
rect 1330 27402 1364 27436
rect 1330 27334 1364 27368
rect 1330 27266 1364 27300
rect 1330 27198 1364 27232
rect 1330 27130 1364 27164
rect 1330 27062 1364 27096
rect 1330 26994 1364 27028
rect 1330 26926 1364 26960
rect 1330 26858 1364 26892
rect 1330 26790 1364 26824
rect 1488 27674 1522 27708
rect 1488 27606 1522 27640
rect 1488 27538 1522 27572
rect 1488 27470 1522 27504
rect 1488 27402 1522 27436
rect 1488 27334 1522 27368
rect 1488 27266 1522 27300
rect 1488 27198 1522 27232
rect 1488 27130 1522 27164
rect 1488 27062 1522 27096
rect 1488 26994 1522 27028
rect 1488 26926 1522 26960
rect 1488 26858 1522 26892
rect 1488 26790 1522 26824
rect 1646 27674 1680 27708
rect 1646 27606 1680 27640
rect 1646 27538 1680 27572
rect 1646 27470 1680 27504
rect 1646 27402 1680 27436
rect 1646 27334 1680 27368
rect 1646 27266 1680 27300
rect 1646 27198 1680 27232
rect 1646 27130 1680 27164
rect 1646 27062 1680 27096
rect 1646 26994 1680 27028
rect 1646 26926 1680 26960
rect 1646 26858 1680 26892
rect 1646 26790 1680 26824
rect -3579 19398 -2603 19432
rect -2343 19398 -1367 19432
rect -1107 19398 -131 19432
rect 129 19398 1105 19432
rect 1365 19398 2341 19432
rect 2601 19398 3577 19432
rect -3579 19140 -2603 19174
rect -2343 19140 -1367 19174
rect -1107 19140 -131 19174
rect 129 19140 1105 19174
rect 1365 19140 2341 19174
rect 2601 19140 3577 19174
rect -3579 18808 -2603 18842
rect -2343 18808 -1367 18842
rect -1107 18808 -131 18842
rect 129 18808 1105 18842
rect 1365 18808 2341 18842
rect 2601 18808 3577 18842
rect -3579 18550 -2603 18584
rect -2343 18550 -1367 18584
rect -1107 18550 -131 18584
rect 129 18550 1105 18584
rect 1365 18550 2341 18584
rect 2601 18550 3577 18584
<< psubdiff >>
rect -7264 32038 -7168 32072
rect -4236 32038 -4140 32072
rect -7264 31976 -7230 32038
rect -4174 31976 -4140 32038
rect -7264 30700 -7230 30762
rect 4144 32008 4261 32042
rect 4295 32008 4329 32042
rect 4363 32008 4397 32042
rect 4431 32008 4465 32042
rect 4499 32008 4533 32042
rect 4567 32008 4601 32042
rect 4635 32008 4669 32042
rect 4703 32008 4737 32042
rect 4771 32008 4805 32042
rect 4839 32008 4873 32042
rect 4907 32008 4941 32042
rect 4975 32008 5009 32042
rect 5043 32008 5077 32042
rect 5111 32008 5145 32042
rect 5179 32008 5213 32042
rect 5247 32008 5281 32042
rect 5315 32008 5349 32042
rect 5383 32008 5417 32042
rect 5451 32008 5485 32042
rect 5519 32008 5553 32042
rect 5587 32008 5621 32042
rect 5655 32008 5689 32042
rect 5723 32008 5757 32042
rect 5791 32008 5825 32042
rect 5859 32008 5893 32042
rect 5927 32008 5961 32042
rect 5995 32008 6029 32042
rect 6063 32008 6097 32042
rect 6131 32008 6165 32042
rect 6199 32008 6233 32042
rect 6267 32008 6301 32042
rect 6335 32008 6369 32042
rect 6403 32008 6437 32042
rect 6471 32008 6505 32042
rect 6539 32008 6573 32042
rect 6607 32008 6641 32042
rect 6675 32008 6709 32042
rect 6743 32008 6777 32042
rect 6811 32008 6845 32042
rect 6879 32008 6913 32042
rect 6947 32008 6981 32042
rect 7015 32008 7049 32042
rect 7083 32008 7117 32042
rect 7151 32008 7268 32042
rect 4144 31934 4178 32008
rect 7234 31934 7268 32008
rect 4144 31866 4178 31900
rect 4144 31798 4178 31832
rect 4144 31730 4178 31764
rect 4144 31662 4178 31696
rect 4144 31594 4178 31628
rect 4144 31526 4178 31560
rect 4144 31458 4178 31492
rect 4144 31390 4178 31424
rect 4144 31322 4178 31356
rect 4144 31254 4178 31288
rect 4144 31186 4178 31220
rect -4174 30700 -4140 30762
rect -7264 30666 -7168 30700
rect -4236 30666 -4140 30700
rect -7264 30538 -7168 30572
rect -4236 30538 -4140 30572
rect -7264 30476 -7230 30538
rect -4174 30476 -4140 30538
rect -7264 29200 -7230 29262
rect 4144 31118 4178 31152
rect 4144 31050 4178 31084
rect 4144 30982 4178 31016
rect 4144 30914 4178 30948
rect 4144 30846 4178 30880
rect 4144 30778 4178 30812
rect 7234 31866 7268 31900
rect 7234 31798 7268 31832
rect 7234 31730 7268 31764
rect 7234 31662 7268 31696
rect 7234 31594 7268 31628
rect 7234 31526 7268 31560
rect 7234 31458 7268 31492
rect 7234 31390 7268 31424
rect 7234 31322 7268 31356
rect 7234 31254 7268 31288
rect 7234 31186 7268 31220
rect 7234 31118 7268 31152
rect 7234 31050 7268 31084
rect 7234 30982 7268 31016
rect 7234 30914 7268 30948
rect 7234 30846 7268 30880
rect 7234 30778 7268 30812
rect 4144 30670 4178 30744
rect 7234 30670 7268 30744
rect 4144 30636 4261 30670
rect 4295 30636 4329 30670
rect 4363 30636 4397 30670
rect 4431 30636 4465 30670
rect 4499 30636 4533 30670
rect 4567 30636 4601 30670
rect 4635 30636 4669 30670
rect 4703 30636 4737 30670
rect 4771 30636 4805 30670
rect 4839 30636 4873 30670
rect 4907 30636 4941 30670
rect 4975 30636 5009 30670
rect 5043 30636 5077 30670
rect 5111 30636 5145 30670
rect 5179 30636 5213 30670
rect 5247 30636 5281 30670
rect 5315 30636 5349 30670
rect 5383 30636 5417 30670
rect 5451 30636 5485 30670
rect 5519 30636 5553 30670
rect 5587 30636 5621 30670
rect 5655 30636 5689 30670
rect 5723 30636 5757 30670
rect 5791 30636 5825 30670
rect 5859 30636 5893 30670
rect 5927 30636 5961 30670
rect 5995 30636 6029 30670
rect 6063 30636 6097 30670
rect 6131 30636 6165 30670
rect 6199 30636 6233 30670
rect 6267 30636 6301 30670
rect 6335 30636 6369 30670
rect 6403 30636 6437 30670
rect 6471 30636 6505 30670
rect 6539 30636 6573 30670
rect 6607 30636 6641 30670
rect 6675 30636 6709 30670
rect 6743 30636 6777 30670
rect 6811 30636 6845 30670
rect 6879 30636 6913 30670
rect 6947 30636 6981 30670
rect 7015 30636 7049 30670
rect 7083 30636 7117 30670
rect 7151 30636 7268 30670
rect 4144 30528 4261 30562
rect 4295 30528 4329 30562
rect 4363 30528 4397 30562
rect 4431 30528 4465 30562
rect 4499 30528 4533 30562
rect 4567 30528 4601 30562
rect 4635 30528 4669 30562
rect 4703 30528 4737 30562
rect 4771 30528 4805 30562
rect 4839 30528 4873 30562
rect 4907 30528 4941 30562
rect 4975 30528 5009 30562
rect 5043 30528 5077 30562
rect 5111 30528 5145 30562
rect 5179 30528 5213 30562
rect 5247 30528 5281 30562
rect 5315 30528 5349 30562
rect 5383 30528 5417 30562
rect 5451 30528 5485 30562
rect 5519 30528 5553 30562
rect 5587 30528 5621 30562
rect 5655 30528 5689 30562
rect 5723 30528 5757 30562
rect 5791 30528 5825 30562
rect 5859 30528 5893 30562
rect 5927 30528 5961 30562
rect 5995 30528 6029 30562
rect 6063 30528 6097 30562
rect 6131 30528 6165 30562
rect 6199 30528 6233 30562
rect 6267 30528 6301 30562
rect 6335 30528 6369 30562
rect 6403 30528 6437 30562
rect 6471 30528 6505 30562
rect 6539 30528 6573 30562
rect 6607 30528 6641 30562
rect 6675 30528 6709 30562
rect 6743 30528 6777 30562
rect 6811 30528 6845 30562
rect 6879 30528 6913 30562
rect 6947 30528 6981 30562
rect 7015 30528 7049 30562
rect 7083 30528 7117 30562
rect 7151 30528 7268 30562
rect 4144 30454 4178 30528
rect 7234 30454 7268 30528
rect 4144 30386 4178 30420
rect 4144 30318 4178 30352
rect 4144 30250 4178 30284
rect 4144 30182 4178 30216
rect 4144 30114 4178 30148
rect 4144 30046 4178 30080
rect 4144 29978 4178 30012
rect 4144 29910 4178 29944
rect 4144 29842 4178 29876
rect 4144 29774 4178 29808
rect 4144 29706 4178 29740
rect 4144 29638 4178 29672
rect 4144 29570 4178 29604
rect 4144 29502 4178 29536
rect -4174 29200 -4140 29262
rect -7264 29166 -7168 29200
rect -4236 29166 -4140 29200
rect 4144 29434 4178 29468
rect 4144 29366 4178 29400
rect 4144 29298 4178 29332
rect 7234 30386 7268 30420
rect 7234 30318 7268 30352
rect 7234 30250 7268 30284
rect 7234 30182 7268 30216
rect 7234 30114 7268 30148
rect 7234 30046 7268 30080
rect 7234 29978 7268 30012
rect 7234 29910 7268 29944
rect 7234 29842 7268 29876
rect 7234 29774 7268 29808
rect 7234 29706 7268 29740
rect 7234 29638 7268 29672
rect 7234 29570 7268 29604
rect 7234 29502 7268 29536
rect 7234 29434 7268 29468
rect 7234 29366 7268 29400
rect 7234 29298 7268 29332
rect 4144 29190 4178 29264
rect 7234 29190 7268 29264
rect 4144 29156 4261 29190
rect 4295 29156 4329 29190
rect 4363 29156 4397 29190
rect 4431 29156 4465 29190
rect 4499 29156 4533 29190
rect 4567 29156 4601 29190
rect 4635 29156 4669 29190
rect 4703 29156 4737 29190
rect 4771 29156 4805 29190
rect 4839 29156 4873 29190
rect 4907 29156 4941 29190
rect 4975 29156 5009 29190
rect 5043 29156 5077 29190
rect 5111 29156 5145 29190
rect 5179 29156 5213 29190
rect 5247 29156 5281 29190
rect 5315 29156 5349 29190
rect 5383 29156 5417 29190
rect 5451 29156 5485 29190
rect 5519 29156 5553 29190
rect 5587 29156 5621 29190
rect 5655 29156 5689 29190
rect 5723 29156 5757 29190
rect 5791 29156 5825 29190
rect 5859 29156 5893 29190
rect 5927 29156 5961 29190
rect 5995 29156 6029 29190
rect 6063 29156 6097 29190
rect 6131 29156 6165 29190
rect 6199 29156 6233 29190
rect 6267 29156 6301 29190
rect 6335 29156 6369 29190
rect 6403 29156 6437 29190
rect 6471 29156 6505 29190
rect 6539 29156 6573 29190
rect 6607 29156 6641 29190
rect 6675 29156 6709 29190
rect 6743 29156 6777 29190
rect 6811 29156 6845 29190
rect 6879 29156 6913 29190
rect 6947 29156 6981 29190
rect 7015 29156 7049 29190
rect 7083 29156 7117 29190
rect 7151 29156 7268 29190
rect -685 26321 -562 26355
rect -528 26321 -494 26355
rect -460 26321 -426 26355
rect -392 26321 -358 26355
rect -324 26321 -290 26355
rect -256 26321 -222 26355
rect -188 26321 -154 26355
rect -120 26321 -86 26355
rect -52 26321 -18 26355
rect 16 26321 50 26355
rect 84 26321 118 26355
rect 152 26321 186 26355
rect 220 26321 254 26355
rect 288 26321 322 26355
rect 356 26321 390 26355
rect 424 26321 458 26355
rect 492 26321 526 26355
rect 560 26321 683 26355
rect -685 26242 -651 26321
rect -685 26174 -651 26208
rect 649 26242 683 26321
rect -685 26106 -651 26140
rect -685 26038 -651 26072
rect -685 25970 -651 26004
rect -685 25902 -651 25936
rect -685 25834 -651 25868
rect -685 25766 -651 25800
rect -685 25698 -651 25732
rect -685 25630 -651 25664
rect -685 25562 -651 25596
rect -685 25494 -651 25528
rect -685 25426 -651 25460
rect -685 25358 -651 25392
rect -685 25290 -651 25324
rect -685 25222 -651 25256
rect -685 25154 -651 25188
rect 649 26174 683 26208
rect 649 26106 683 26140
rect 649 26038 683 26072
rect 649 25970 683 26004
rect 649 25902 683 25936
rect 649 25834 683 25868
rect 649 25766 683 25800
rect 649 25698 683 25732
rect 649 25630 683 25664
rect 649 25562 683 25596
rect 649 25494 683 25528
rect 649 25426 683 25460
rect 649 25358 683 25392
rect 649 25290 683 25324
rect 649 25222 683 25256
rect -685 25041 -651 25120
rect 649 25154 683 25188
rect 649 25041 683 25120
rect -685 25007 -562 25041
rect -528 25007 -494 25041
rect -460 25007 -426 25041
rect -392 25007 -358 25041
rect -324 25007 -290 25041
rect -256 25007 -222 25041
rect -188 25007 -154 25041
rect -120 25007 -86 25041
rect -52 25007 -18 25041
rect 16 25007 50 25041
rect 84 25007 118 25041
rect 152 25007 186 25041
rect 220 25007 254 25041
rect 288 25007 322 25041
rect 356 25007 390 25041
rect 424 25007 458 25041
rect 492 25007 526 25041
rect 560 25007 683 25041
rect -685 24801 -562 24835
rect -528 24801 -494 24835
rect -460 24801 -426 24835
rect -392 24801 -358 24835
rect -324 24801 -290 24835
rect -256 24801 -222 24835
rect -188 24801 -154 24835
rect -120 24801 -86 24835
rect -52 24801 -18 24835
rect 16 24801 50 24835
rect 84 24801 118 24835
rect 152 24801 186 24835
rect 220 24801 254 24835
rect 288 24801 322 24835
rect 356 24801 390 24835
rect 424 24801 458 24835
rect 492 24801 526 24835
rect 560 24801 683 24835
rect -685 24722 -651 24801
rect -685 24654 -651 24688
rect 649 24722 683 24801
rect -685 24586 -651 24620
rect -685 24518 -651 24552
rect -685 24450 -651 24484
rect -685 24382 -651 24416
rect -685 24314 -651 24348
rect -685 24246 -651 24280
rect -685 24178 -651 24212
rect -685 24110 -651 24144
rect -685 24042 -651 24076
rect -685 23974 -651 24008
rect -685 23906 -651 23940
rect -685 23838 -651 23872
rect -685 23770 -651 23804
rect -685 23702 -651 23736
rect -685 23634 -651 23668
rect 649 24654 683 24688
rect 649 24586 683 24620
rect 649 24518 683 24552
rect 649 24450 683 24484
rect 649 24382 683 24416
rect 649 24314 683 24348
rect 649 24246 683 24280
rect 649 24178 683 24212
rect 649 24110 683 24144
rect 649 24042 683 24076
rect 649 23974 683 24008
rect 649 23906 683 23940
rect 649 23838 683 23872
rect 649 23770 683 23804
rect 649 23702 683 23736
rect -685 23521 -651 23600
rect 649 23634 683 23668
rect 649 23521 683 23600
rect -685 23487 -562 23521
rect -528 23487 -494 23521
rect -460 23487 -426 23521
rect -392 23487 -358 23521
rect -324 23487 -290 23521
rect -256 23487 -222 23521
rect -188 23487 -154 23521
rect -120 23487 -86 23521
rect -52 23487 -18 23521
rect 16 23487 50 23521
rect 84 23487 118 23521
rect 152 23487 186 23521
rect 220 23487 254 23521
rect 288 23487 322 23521
rect 356 23487 390 23521
rect 424 23487 458 23521
rect 492 23487 526 23521
rect 560 23487 683 23521
rect -1676 23280 -1578 23314
rect -1544 23280 -1510 23314
rect -1476 23280 -1442 23314
rect -1408 23280 -1374 23314
rect -1340 23280 -1306 23314
rect -1272 23280 -1238 23314
rect -1204 23280 -1170 23314
rect -1136 23280 -1102 23314
rect -1068 23280 -1034 23314
rect -1000 23280 -966 23314
rect -932 23280 -898 23314
rect -864 23280 -830 23314
rect -796 23280 -762 23314
rect -728 23280 -694 23314
rect -660 23280 -626 23314
rect -592 23280 -558 23314
rect -524 23280 -490 23314
rect -456 23280 -422 23314
rect -388 23280 -354 23314
rect -320 23280 -286 23314
rect -252 23280 -218 23314
rect -184 23280 -150 23314
rect -116 23280 -82 23314
rect -48 23280 -14 23314
rect 20 23280 54 23314
rect 88 23280 122 23314
rect 156 23280 190 23314
rect 224 23280 258 23314
rect 292 23280 326 23314
rect 360 23280 394 23314
rect 428 23280 462 23314
rect 496 23280 530 23314
rect 564 23280 598 23314
rect 632 23280 666 23314
rect 700 23280 734 23314
rect 768 23280 802 23314
rect 836 23280 870 23314
rect 904 23280 938 23314
rect 972 23280 1006 23314
rect 1040 23280 1074 23314
rect 1108 23280 1142 23314
rect 1176 23280 1210 23314
rect 1244 23280 1278 23314
rect 1312 23280 1346 23314
rect 1380 23280 1414 23314
rect 1448 23280 1482 23314
rect 1516 23280 1550 23314
rect 1584 23280 1682 23314
rect -1676 23201 -1642 23280
rect -1676 23133 -1642 23167
rect 1648 23201 1682 23280
rect -1676 23065 -1642 23099
rect -1676 22997 -1642 23031
rect -1676 22929 -1642 22963
rect -1676 22861 -1642 22895
rect -1676 22793 -1642 22827
rect -1676 22725 -1642 22759
rect -1676 22657 -1642 22691
rect -1676 22589 -1642 22623
rect -1676 22521 -1642 22555
rect -1676 22453 -1642 22487
rect -1676 22385 -1642 22419
rect -1676 22317 -1642 22351
rect -1676 22249 -1642 22283
rect -1676 22181 -1642 22215
rect -1676 22113 -1642 22147
rect 1648 23133 1682 23167
rect 1648 23065 1682 23099
rect 1648 22997 1682 23031
rect 1648 22929 1682 22963
rect 1648 22861 1682 22895
rect 1648 22793 1682 22827
rect 1648 22725 1682 22759
rect 1648 22657 1682 22691
rect 1648 22589 1682 22623
rect 1648 22521 1682 22555
rect 1648 22453 1682 22487
rect 1648 22385 1682 22419
rect 1648 22317 1682 22351
rect 1648 22249 1682 22283
rect 1648 22181 1682 22215
rect -1676 22000 -1642 22079
rect 1648 22113 1682 22147
rect 1648 22000 1682 22079
rect -1676 21966 -1578 22000
rect -1544 21966 -1510 22000
rect -1476 21966 -1442 22000
rect -1408 21966 -1374 22000
rect -1340 21966 -1306 22000
rect -1272 21966 -1238 22000
rect -1204 21966 -1170 22000
rect -1136 21966 -1102 22000
rect -1068 21966 -1034 22000
rect -1000 21966 -966 22000
rect -932 21966 -898 22000
rect -864 21966 -830 22000
rect -796 21966 -762 22000
rect -728 21966 -694 22000
rect -660 21966 -626 22000
rect -592 21966 -558 22000
rect -524 21966 -490 22000
rect -456 21966 -422 22000
rect -388 21966 -354 22000
rect -320 21966 -286 22000
rect -252 21966 -218 22000
rect -184 21966 -150 22000
rect -116 21966 -82 22000
rect -48 21966 -14 22000
rect 20 21966 54 22000
rect 88 21966 122 22000
rect 156 21966 190 22000
rect 224 21966 258 22000
rect 292 21966 326 22000
rect 360 21966 394 22000
rect 428 21966 462 22000
rect 496 21966 530 22000
rect 564 21966 598 22000
rect 632 21966 666 22000
rect 700 21966 734 22000
rect 768 21966 802 22000
rect 836 21966 870 22000
rect 904 21966 938 22000
rect 972 21966 1006 22000
rect 1040 21966 1074 22000
rect 1108 21966 1142 22000
rect 1176 21966 1210 22000
rect 1244 21966 1278 22000
rect 1312 21966 1346 22000
rect 1380 21966 1414 22000
rect 1448 21966 1482 22000
rect 1516 21966 1550 22000
rect 1584 21966 1682 22000
rect -1936 21760 -1818 21794
rect -1784 21760 -1750 21794
rect -1716 21760 -1682 21794
rect -1648 21760 -1614 21794
rect -1580 21760 -1546 21794
rect -1512 21760 -1478 21794
rect -1444 21760 -1410 21794
rect -1376 21760 -1342 21794
rect -1308 21760 -1274 21794
rect -1240 21760 -1206 21794
rect -1172 21760 -1138 21794
rect -1104 21760 -1070 21794
rect -1036 21760 -1002 21794
rect -968 21760 -934 21794
rect -900 21760 -866 21794
rect -832 21760 -798 21794
rect -764 21760 -730 21794
rect -696 21760 -662 21794
rect -628 21760 -594 21794
rect -560 21760 -526 21794
rect -492 21760 -458 21794
rect -424 21760 -390 21794
rect -356 21760 -322 21794
rect -288 21760 -254 21794
rect -220 21760 -186 21794
rect -152 21760 -118 21794
rect -84 21760 -50 21794
rect -16 21760 18 21794
rect 52 21760 86 21794
rect 120 21760 154 21794
rect 188 21760 222 21794
rect 256 21760 290 21794
rect 324 21760 358 21794
rect 392 21760 426 21794
rect 460 21760 494 21794
rect 528 21760 562 21794
rect 596 21760 630 21794
rect 664 21760 698 21794
rect 732 21760 766 21794
rect 800 21760 834 21794
rect 868 21760 902 21794
rect 936 21760 970 21794
rect 1004 21760 1038 21794
rect 1072 21760 1106 21794
rect 1140 21760 1174 21794
rect 1208 21760 1242 21794
rect 1276 21760 1310 21794
rect 1344 21760 1378 21794
rect 1412 21760 1446 21794
rect 1480 21760 1514 21794
rect 1548 21760 1582 21794
rect 1616 21760 1650 21794
rect 1684 21760 1718 21794
rect 1752 21760 1786 21794
rect 1820 21760 1938 21794
rect -1936 21681 -1902 21760
rect -1936 21613 -1902 21647
rect 1904 21681 1938 21760
rect -1936 21545 -1902 21579
rect -1936 21477 -1902 21511
rect -1936 21409 -1902 21443
rect -1936 21341 -1902 21375
rect -1936 21273 -1902 21307
rect -1936 21205 -1902 21239
rect -1936 21137 -1902 21171
rect -1936 21069 -1902 21103
rect -1936 21001 -1902 21035
rect -1936 20933 -1902 20967
rect -1936 20865 -1902 20899
rect -1936 20797 -1902 20831
rect -1936 20729 -1902 20763
rect -1936 20661 -1902 20695
rect -1936 20593 -1902 20627
rect 1904 21613 1938 21647
rect 1904 21545 1938 21579
rect 1904 21477 1938 21511
rect 1904 21409 1938 21443
rect 1904 21341 1938 21375
rect 1904 21273 1938 21307
rect 1904 21205 1938 21239
rect 1904 21137 1938 21171
rect 1904 21069 1938 21103
rect 1904 21001 1938 21035
rect 1904 20933 1938 20967
rect 1904 20865 1938 20899
rect 1904 20797 1938 20831
rect 1904 20729 1938 20763
rect 1904 20661 1938 20695
rect -1936 20480 -1902 20559
rect 1904 20593 1938 20627
rect 1904 20480 1938 20559
rect -1936 20446 -1818 20480
rect -1784 20446 -1750 20480
rect -1716 20446 -1682 20480
rect -1648 20446 -1614 20480
rect -1580 20446 -1546 20480
rect -1512 20446 -1478 20480
rect -1444 20446 -1410 20480
rect -1376 20446 -1342 20480
rect -1308 20446 -1274 20480
rect -1240 20446 -1206 20480
rect -1172 20446 -1138 20480
rect -1104 20446 -1070 20480
rect -1036 20446 -1002 20480
rect -968 20446 -934 20480
rect -900 20446 -866 20480
rect -832 20446 -798 20480
rect -764 20446 -730 20480
rect -696 20446 -662 20480
rect -628 20446 -594 20480
rect -560 20446 -526 20480
rect -492 20446 -458 20480
rect -424 20446 -390 20480
rect -356 20446 -322 20480
rect -288 20446 -254 20480
rect -220 20446 -186 20480
rect -152 20446 -118 20480
rect -84 20446 -50 20480
rect -16 20446 18 20480
rect 52 20446 86 20480
rect 120 20446 154 20480
rect 188 20446 222 20480
rect 256 20446 290 20480
rect 324 20446 358 20480
rect 392 20446 426 20480
rect 460 20446 494 20480
rect 528 20446 562 20480
rect 596 20446 630 20480
rect 664 20446 698 20480
rect 732 20446 766 20480
rect 800 20446 834 20480
rect 868 20446 902 20480
rect 936 20446 970 20480
rect 1004 20446 1038 20480
rect 1072 20446 1106 20480
rect 1140 20446 1174 20480
rect 1208 20446 1242 20480
rect 1276 20446 1310 20480
rect 1344 20446 1378 20480
rect 1412 20446 1446 20480
rect 1480 20446 1514 20480
rect 1548 20446 1582 20480
rect 1616 20446 1650 20480
rect 1684 20446 1718 20480
rect 1752 20446 1786 20480
rect 1820 20446 1938 20480
rect -1004 18132 -908 18166
rect 902 18132 998 18166
rect -1004 18070 -970 18132
rect 964 18070 998 18132
rect -1004 17680 -970 17742
rect 964 17680 998 17742
rect -1004 17646 -908 17680
rect 902 17646 998 17680
rect -784 17507 -688 17541
rect 686 17507 782 17541
rect -784 17445 -750 17507
rect 748 17445 782 17507
rect -784 17155 -750 17217
rect 748 17155 782 17217
rect -784 17121 -688 17155
rect 686 17121 782 17155
rect -3719 16982 -3623 17016
rect 3623 16982 3719 17016
rect -3719 16920 -3685 16982
rect 3685 16920 3719 16982
rect -3719 16530 -3685 16592
rect 3685 16530 3719 16592
rect -3719 16496 -3623 16530
rect 3623 16496 3719 16530
rect -3240 15220 -3120 15244
rect -3240 15076 -3120 15100
rect -3240 12220 -3120 12244
rect -3240 12076 -3120 12100
rect -3240 9220 -3120 9244
rect -3240 9076 -3120 9100
rect -3240 6220 -3120 6244
rect -3240 6076 -3120 6100
rect -3240 3220 -3120 3244
rect -3240 3076 -3120 3100
rect 3130 15220 3250 15244
rect 3130 15076 3250 15100
rect 3130 12220 3250 12244
rect 3130 12076 3250 12100
rect 3130 9220 3250 9244
rect 3130 9076 3250 9100
rect 3130 6220 3250 6244
rect 3130 6076 3250 6100
rect 3130 3220 3250 3244
rect 3130 3076 3250 3100
<< nsubdiff >>
rect -3286 31108 -3174 31142
rect -3140 31108 -3106 31142
rect -3072 31108 -3038 31142
rect -3004 31108 -2970 31142
rect -2936 31108 -2902 31142
rect -2868 31108 -2834 31142
rect -2800 31108 -2766 31142
rect -2732 31108 -2698 31142
rect -2664 31108 -2630 31142
rect -2596 31108 -2562 31142
rect -2528 31108 -2494 31142
rect -2460 31108 -2426 31142
rect -2392 31108 -2358 31142
rect -2324 31108 -2290 31142
rect -2256 31108 -2222 31142
rect -2188 31108 -2154 31142
rect -2120 31108 -2086 31142
rect -2052 31108 -2018 31142
rect -1984 31108 -1950 31142
rect -1916 31108 -1882 31142
rect -1848 31108 -1814 31142
rect -1780 31108 -1746 31142
rect -1712 31108 -1678 31142
rect -1644 31108 -1610 31142
rect -1576 31108 -1542 31142
rect -1508 31108 -1474 31142
rect -1440 31108 -1406 31142
rect -1372 31108 -1338 31142
rect -1304 31108 -1270 31142
rect -1236 31108 -1202 31142
rect -1168 31108 -1134 31142
rect -1100 31108 -1066 31142
rect -1032 31108 -998 31142
rect -964 31108 -930 31142
rect -896 31108 -862 31142
rect -828 31108 -794 31142
rect -760 31108 -726 31142
rect -692 31108 -658 31142
rect -624 31108 -590 31142
rect -556 31108 -522 31142
rect -488 31108 -454 31142
rect -420 31108 -386 31142
rect -352 31108 -318 31142
rect -284 31108 -250 31142
rect -216 31108 -182 31142
rect -148 31108 -114 31142
rect -80 31108 -46 31142
rect -12 31108 22 31142
rect 56 31108 90 31142
rect 124 31108 158 31142
rect 192 31108 226 31142
rect 260 31108 294 31142
rect 328 31108 362 31142
rect 396 31108 430 31142
rect 464 31108 498 31142
rect 532 31108 566 31142
rect 600 31108 634 31142
rect 668 31108 702 31142
rect 736 31108 770 31142
rect 804 31108 838 31142
rect 872 31108 906 31142
rect 940 31108 974 31142
rect 1008 31108 1042 31142
rect 1076 31108 1110 31142
rect 1144 31108 1178 31142
rect 1212 31108 1246 31142
rect 1280 31108 1314 31142
rect 1348 31108 1382 31142
rect 1416 31108 1450 31142
rect 1484 31108 1518 31142
rect 1552 31108 1586 31142
rect 1620 31108 1654 31142
rect 1688 31108 1722 31142
rect 1756 31108 1790 31142
rect 1824 31108 1858 31142
rect 1892 31108 1926 31142
rect 1960 31108 1994 31142
rect 2028 31108 2062 31142
rect 2096 31108 2130 31142
rect 2164 31108 2198 31142
rect 2232 31108 2266 31142
rect 2300 31108 2334 31142
rect 2368 31108 2402 31142
rect 2436 31108 2470 31142
rect 2504 31108 2538 31142
rect 2572 31108 2606 31142
rect 2640 31108 2674 31142
rect 2708 31108 2742 31142
rect 2776 31108 2810 31142
rect 2844 31108 2878 31142
rect 2912 31108 2946 31142
rect 2980 31108 3014 31142
rect 3048 31108 3082 31142
rect 3116 31108 3150 31142
rect 3184 31108 3296 31142
rect -3286 31020 -3252 31108
rect -3286 30952 -3252 30986
rect 3262 31020 3296 31108
rect -3286 30884 -3252 30918
rect -3286 30816 -3252 30850
rect -3286 30748 -3252 30782
rect -3286 30680 -3252 30714
rect -3286 30612 -3252 30646
rect -3286 30544 -3252 30578
rect -3286 30476 -3252 30510
rect -3286 30408 -3252 30442
rect -3286 30340 -3252 30374
rect -3286 30272 -3252 30306
rect -3286 30204 -3252 30238
rect -3286 30136 -3252 30170
rect -3286 30068 -3252 30102
rect -3286 30000 -3252 30034
rect -3286 29932 -3252 29966
rect 3262 30952 3296 30986
rect 3262 30884 3296 30918
rect 3262 30816 3296 30850
rect 3262 30748 3296 30782
rect 3262 30680 3296 30714
rect 3262 30612 3296 30646
rect 3262 30544 3296 30578
rect 3262 30476 3296 30510
rect 3262 30408 3296 30442
rect 3262 30340 3296 30374
rect 3262 30272 3296 30306
rect 3262 30204 3296 30238
rect 3262 30136 3296 30170
rect 3262 30068 3296 30102
rect 3262 30000 3296 30034
rect -3286 29810 -3252 29898
rect 3262 29932 3296 29966
rect 3262 29810 3296 29898
rect -3286 29776 -3174 29810
rect -3140 29776 -3106 29810
rect -3072 29776 -3038 29810
rect -3004 29776 -2970 29810
rect -2936 29776 -2902 29810
rect -2868 29776 -2834 29810
rect -2800 29776 -2766 29810
rect -2732 29776 -2698 29810
rect -2664 29776 -2630 29810
rect -2596 29776 -2562 29810
rect -2528 29776 -2494 29810
rect -2460 29776 -2426 29810
rect -2392 29776 -2358 29810
rect -2324 29776 -2290 29810
rect -2256 29776 -2222 29810
rect -2188 29776 -2154 29810
rect -2120 29776 -2086 29810
rect -2052 29776 -2018 29810
rect -1984 29776 -1950 29810
rect -1916 29776 -1882 29810
rect -1848 29776 -1814 29810
rect -1780 29776 -1746 29810
rect -1712 29776 -1678 29810
rect -1644 29776 -1610 29810
rect -1576 29776 -1542 29810
rect -1508 29776 -1474 29810
rect -1440 29776 -1406 29810
rect -1372 29776 -1338 29810
rect -1304 29776 -1270 29810
rect -1236 29776 -1202 29810
rect -1168 29776 -1134 29810
rect -1100 29776 -1066 29810
rect -1032 29776 -998 29810
rect -964 29776 -930 29810
rect -896 29776 -862 29810
rect -828 29776 -794 29810
rect -760 29776 -726 29810
rect -692 29776 -658 29810
rect -624 29776 -590 29810
rect -556 29776 -522 29810
rect -488 29776 -454 29810
rect -420 29776 -386 29810
rect -352 29776 -318 29810
rect -284 29776 -250 29810
rect -216 29776 -182 29810
rect -148 29776 -114 29810
rect -80 29776 -46 29810
rect -12 29776 22 29810
rect 56 29776 90 29810
rect 124 29776 158 29810
rect 192 29776 226 29810
rect 260 29776 294 29810
rect 328 29776 362 29810
rect 396 29776 430 29810
rect 464 29776 498 29810
rect 532 29776 566 29810
rect 600 29776 634 29810
rect 668 29776 702 29810
rect 736 29776 770 29810
rect 804 29776 838 29810
rect 872 29776 906 29810
rect 940 29776 974 29810
rect 1008 29776 1042 29810
rect 1076 29776 1110 29810
rect 1144 29776 1178 29810
rect 1212 29776 1246 29810
rect 1280 29776 1314 29810
rect 1348 29776 1382 29810
rect 1416 29776 1450 29810
rect 1484 29776 1518 29810
rect 1552 29776 1586 29810
rect 1620 29776 1654 29810
rect 1688 29776 1722 29810
rect 1756 29776 1790 29810
rect 1824 29776 1858 29810
rect 1892 29776 1926 29810
rect 1960 29776 1994 29810
rect 2028 29776 2062 29810
rect 2096 29776 2130 29810
rect 2164 29776 2198 29810
rect 2232 29776 2266 29810
rect 2300 29776 2334 29810
rect 2368 29776 2402 29810
rect 2436 29776 2470 29810
rect 2504 29776 2538 29810
rect 2572 29776 2606 29810
rect 2640 29776 2674 29810
rect 2708 29776 2742 29810
rect 2776 29776 2810 29810
rect 2844 29776 2878 29810
rect 2912 29776 2946 29810
rect 2980 29776 3014 29810
rect 3048 29776 3082 29810
rect 3116 29776 3150 29810
rect 3184 29776 3296 29810
rect -1786 29438 -1679 29472
rect -1645 29438 -1611 29472
rect -1577 29438 -1543 29472
rect -1509 29438 -1475 29472
rect -1441 29438 -1407 29472
rect -1373 29438 -1339 29472
rect -1305 29438 -1271 29472
rect -1237 29438 -1203 29472
rect -1169 29438 -1135 29472
rect -1101 29438 -1067 29472
rect -1033 29438 -999 29472
rect -965 29438 -931 29472
rect -897 29438 -863 29472
rect -829 29438 -795 29472
rect -761 29438 -727 29472
rect -693 29438 -659 29472
rect -625 29438 -591 29472
rect -557 29438 -523 29472
rect -489 29438 -455 29472
rect -421 29438 -387 29472
rect -353 29438 -319 29472
rect -285 29438 -251 29472
rect -217 29438 -183 29472
rect -149 29438 -115 29472
rect -81 29438 -47 29472
rect -13 29438 21 29472
rect 55 29438 89 29472
rect 123 29438 157 29472
rect 191 29438 225 29472
rect 259 29438 293 29472
rect 327 29438 361 29472
rect 395 29438 429 29472
rect 463 29438 497 29472
rect 531 29438 565 29472
rect 599 29438 633 29472
rect 667 29438 701 29472
rect 735 29438 769 29472
rect 803 29438 837 29472
rect 871 29438 905 29472
rect 939 29438 973 29472
rect 1007 29438 1041 29472
rect 1075 29438 1109 29472
rect 1143 29438 1177 29472
rect 1211 29438 1245 29472
rect 1279 29438 1313 29472
rect 1347 29438 1381 29472
rect 1415 29438 1449 29472
rect 1483 29438 1517 29472
rect 1551 29438 1585 29472
rect 1619 29438 1653 29472
rect 1687 29438 1794 29472
rect -1786 29350 -1752 29438
rect -1786 29282 -1752 29316
rect 1760 29350 1794 29438
rect -1786 29214 -1752 29248
rect -1786 29146 -1752 29180
rect -1786 29078 -1752 29112
rect -1786 29010 -1752 29044
rect -1786 28942 -1752 28976
rect -1786 28874 -1752 28908
rect -1786 28806 -1752 28840
rect -1786 28738 -1752 28772
rect -1786 28670 -1752 28704
rect -1786 28602 -1752 28636
rect -1786 28534 -1752 28568
rect -1786 28466 -1752 28500
rect -1786 28398 -1752 28432
rect -1786 28330 -1752 28364
rect -1786 28262 -1752 28296
rect 1760 29282 1794 29316
rect 1760 29214 1794 29248
rect 1760 29146 1794 29180
rect 1760 29078 1794 29112
rect 1760 29010 1794 29044
rect 1760 28942 1794 28976
rect 1760 28874 1794 28908
rect 1760 28806 1794 28840
rect 1760 28738 1794 28772
rect 1760 28670 1794 28704
rect 1760 28602 1794 28636
rect 1760 28534 1794 28568
rect 1760 28466 1794 28500
rect 1760 28398 1794 28432
rect 1760 28330 1794 28364
rect -1786 28140 -1752 28228
rect 1760 28262 1794 28296
rect 1760 28140 1794 28228
rect -1786 28106 -1679 28140
rect -1645 28106 -1611 28140
rect -1577 28106 -1543 28140
rect -1509 28106 -1475 28140
rect -1441 28106 -1407 28140
rect -1373 28106 -1339 28140
rect -1305 28106 -1271 28140
rect -1237 28106 -1203 28140
rect -1169 28106 -1135 28140
rect -1101 28106 -1067 28140
rect -1033 28106 -999 28140
rect -965 28106 -931 28140
rect -897 28106 -863 28140
rect -829 28106 -795 28140
rect -761 28106 -727 28140
rect -693 28106 -659 28140
rect -625 28106 -591 28140
rect -557 28106 -523 28140
rect -489 28106 -455 28140
rect -421 28106 -387 28140
rect -353 28106 -319 28140
rect -285 28106 -251 28140
rect -217 28106 -183 28140
rect -149 28106 -115 28140
rect -81 28106 -47 28140
rect -13 28106 21 28140
rect 55 28106 89 28140
rect 123 28106 157 28140
rect 191 28106 225 28140
rect 259 28106 293 28140
rect 327 28106 361 28140
rect 395 28106 429 28140
rect 463 28106 497 28140
rect 531 28106 565 28140
rect 599 28106 633 28140
rect 667 28106 701 28140
rect 735 28106 769 28140
rect 803 28106 837 28140
rect 871 28106 905 28140
rect 939 28106 973 28140
rect 1007 28106 1041 28140
rect 1075 28106 1109 28140
rect 1143 28106 1177 28140
rect 1211 28106 1245 28140
rect 1279 28106 1313 28140
rect 1347 28106 1381 28140
rect 1415 28106 1449 28140
rect 1483 28106 1517 28140
rect 1551 28106 1585 28140
rect 1619 28106 1653 28140
rect 1687 28106 1794 28140
rect -1786 27898 -1679 27932
rect -1645 27898 -1611 27932
rect -1577 27898 -1543 27932
rect -1509 27898 -1475 27932
rect -1441 27898 -1407 27932
rect -1373 27898 -1339 27932
rect -1305 27898 -1271 27932
rect -1237 27898 -1203 27932
rect -1169 27898 -1135 27932
rect -1101 27898 -1067 27932
rect -1033 27898 -999 27932
rect -965 27898 -931 27932
rect -897 27898 -863 27932
rect -829 27898 -795 27932
rect -761 27898 -727 27932
rect -693 27898 -659 27932
rect -625 27898 -591 27932
rect -557 27898 -523 27932
rect -489 27898 -455 27932
rect -421 27898 -387 27932
rect -353 27898 -319 27932
rect -285 27898 -251 27932
rect -217 27898 -183 27932
rect -149 27898 -115 27932
rect -81 27898 -47 27932
rect -13 27898 21 27932
rect 55 27898 89 27932
rect 123 27898 157 27932
rect 191 27898 225 27932
rect 259 27898 293 27932
rect 327 27898 361 27932
rect 395 27898 429 27932
rect 463 27898 497 27932
rect 531 27898 565 27932
rect 599 27898 633 27932
rect 667 27898 701 27932
rect 735 27898 769 27932
rect 803 27898 837 27932
rect 871 27898 905 27932
rect 939 27898 973 27932
rect 1007 27898 1041 27932
rect 1075 27898 1109 27932
rect 1143 27898 1177 27932
rect 1211 27898 1245 27932
rect 1279 27898 1313 27932
rect 1347 27898 1381 27932
rect 1415 27898 1449 27932
rect 1483 27898 1517 27932
rect 1551 27898 1585 27932
rect 1619 27898 1653 27932
rect 1687 27898 1794 27932
rect -1786 27810 -1752 27898
rect -1786 27742 -1752 27776
rect 1760 27810 1794 27898
rect -1786 27674 -1752 27708
rect -1786 27606 -1752 27640
rect -1786 27538 -1752 27572
rect -1786 27470 -1752 27504
rect -1786 27402 -1752 27436
rect -1786 27334 -1752 27368
rect -1786 27266 -1752 27300
rect -1786 27198 -1752 27232
rect -1786 27130 -1752 27164
rect -1786 27062 -1752 27096
rect -1786 26994 -1752 27028
rect -1786 26926 -1752 26960
rect -1786 26858 -1752 26892
rect -1786 26790 -1752 26824
rect -1786 26722 -1752 26756
rect 1760 27742 1794 27776
rect 1760 27674 1794 27708
rect 1760 27606 1794 27640
rect 1760 27538 1794 27572
rect 1760 27470 1794 27504
rect 1760 27402 1794 27436
rect 1760 27334 1794 27368
rect 1760 27266 1794 27300
rect 1760 27198 1794 27232
rect 1760 27130 1794 27164
rect 1760 27062 1794 27096
rect 1760 26994 1794 27028
rect 1760 26926 1794 26960
rect 1760 26858 1794 26892
rect 1760 26790 1794 26824
rect -1786 26600 -1752 26688
rect 1760 26722 1794 26756
rect 1760 26600 1794 26688
rect -1786 26566 -1679 26600
rect -1645 26566 -1611 26600
rect -1577 26566 -1543 26600
rect -1509 26566 -1475 26600
rect -1441 26566 -1407 26600
rect -1373 26566 -1339 26600
rect -1305 26566 -1271 26600
rect -1237 26566 -1203 26600
rect -1169 26566 -1135 26600
rect -1101 26566 -1067 26600
rect -1033 26566 -999 26600
rect -965 26566 -931 26600
rect -897 26566 -863 26600
rect -829 26566 -795 26600
rect -761 26566 -727 26600
rect -693 26566 -659 26600
rect -625 26566 -591 26600
rect -557 26566 -523 26600
rect -489 26566 -455 26600
rect -421 26566 -387 26600
rect -353 26566 -319 26600
rect -285 26566 -251 26600
rect -217 26566 -183 26600
rect -149 26566 -115 26600
rect -81 26566 -47 26600
rect -13 26566 21 26600
rect 55 26566 89 26600
rect 123 26566 157 26600
rect 191 26566 225 26600
rect 259 26566 293 26600
rect 327 26566 361 26600
rect 395 26566 429 26600
rect 463 26566 497 26600
rect 531 26566 565 26600
rect 599 26566 633 26600
rect 667 26566 701 26600
rect 735 26566 769 26600
rect 803 26566 837 26600
rect 871 26566 905 26600
rect 939 26566 973 26600
rect 1007 26566 1041 26600
rect 1075 26566 1109 26600
rect 1143 26566 1177 26600
rect 1211 26566 1245 26600
rect 1279 26566 1313 26600
rect 1347 26566 1381 26600
rect 1415 26566 1449 26600
rect 1483 26566 1517 26600
rect 1551 26566 1585 26600
rect 1619 26566 1653 26600
rect 1687 26566 1794 26600
rect -3774 19512 -3678 19546
rect 3676 19512 3772 19546
rect -3774 19450 -3740 19512
rect 3738 19450 3772 19512
rect -3774 19060 -3740 19122
rect 3738 19060 3772 19122
rect -3774 19026 -3678 19060
rect 3676 19026 3772 19060
rect -3774 18922 -3678 18956
rect 3676 18922 3772 18956
rect -3774 18860 -3740 18922
rect 3738 18860 3772 18922
rect -3774 18470 -3740 18532
rect 3738 18470 3772 18532
rect -3774 18436 -3678 18470
rect 3676 18436 3772 18470
<< psubdiffcont >>
rect -7168 32038 -4236 32072
rect -7264 30762 -7230 31976
rect -4174 30762 -4140 31976
rect 4261 32008 4295 32042
rect 4329 32008 4363 32042
rect 4397 32008 4431 32042
rect 4465 32008 4499 32042
rect 4533 32008 4567 32042
rect 4601 32008 4635 32042
rect 4669 32008 4703 32042
rect 4737 32008 4771 32042
rect 4805 32008 4839 32042
rect 4873 32008 4907 32042
rect 4941 32008 4975 32042
rect 5009 32008 5043 32042
rect 5077 32008 5111 32042
rect 5145 32008 5179 32042
rect 5213 32008 5247 32042
rect 5281 32008 5315 32042
rect 5349 32008 5383 32042
rect 5417 32008 5451 32042
rect 5485 32008 5519 32042
rect 5553 32008 5587 32042
rect 5621 32008 5655 32042
rect 5689 32008 5723 32042
rect 5757 32008 5791 32042
rect 5825 32008 5859 32042
rect 5893 32008 5927 32042
rect 5961 32008 5995 32042
rect 6029 32008 6063 32042
rect 6097 32008 6131 32042
rect 6165 32008 6199 32042
rect 6233 32008 6267 32042
rect 6301 32008 6335 32042
rect 6369 32008 6403 32042
rect 6437 32008 6471 32042
rect 6505 32008 6539 32042
rect 6573 32008 6607 32042
rect 6641 32008 6675 32042
rect 6709 32008 6743 32042
rect 6777 32008 6811 32042
rect 6845 32008 6879 32042
rect 6913 32008 6947 32042
rect 6981 32008 7015 32042
rect 7049 32008 7083 32042
rect 7117 32008 7151 32042
rect 4144 31900 4178 31934
rect 4144 31832 4178 31866
rect 4144 31764 4178 31798
rect 4144 31696 4178 31730
rect 4144 31628 4178 31662
rect 4144 31560 4178 31594
rect 4144 31492 4178 31526
rect 4144 31424 4178 31458
rect 4144 31356 4178 31390
rect 4144 31288 4178 31322
rect 4144 31220 4178 31254
rect 4144 31152 4178 31186
rect -7168 30666 -4236 30700
rect -7168 30538 -4236 30572
rect -7264 29262 -7230 30476
rect -4174 29262 -4140 30476
rect 4144 31084 4178 31118
rect 4144 31016 4178 31050
rect 4144 30948 4178 30982
rect 4144 30880 4178 30914
rect 4144 30812 4178 30846
rect 4144 30744 4178 30778
rect 7234 31900 7268 31934
rect 7234 31832 7268 31866
rect 7234 31764 7268 31798
rect 7234 31696 7268 31730
rect 7234 31628 7268 31662
rect 7234 31560 7268 31594
rect 7234 31492 7268 31526
rect 7234 31424 7268 31458
rect 7234 31356 7268 31390
rect 7234 31288 7268 31322
rect 7234 31220 7268 31254
rect 7234 31152 7268 31186
rect 7234 31084 7268 31118
rect 7234 31016 7268 31050
rect 7234 30948 7268 30982
rect 7234 30880 7268 30914
rect 7234 30812 7268 30846
rect 7234 30744 7268 30778
rect 4261 30636 4295 30670
rect 4329 30636 4363 30670
rect 4397 30636 4431 30670
rect 4465 30636 4499 30670
rect 4533 30636 4567 30670
rect 4601 30636 4635 30670
rect 4669 30636 4703 30670
rect 4737 30636 4771 30670
rect 4805 30636 4839 30670
rect 4873 30636 4907 30670
rect 4941 30636 4975 30670
rect 5009 30636 5043 30670
rect 5077 30636 5111 30670
rect 5145 30636 5179 30670
rect 5213 30636 5247 30670
rect 5281 30636 5315 30670
rect 5349 30636 5383 30670
rect 5417 30636 5451 30670
rect 5485 30636 5519 30670
rect 5553 30636 5587 30670
rect 5621 30636 5655 30670
rect 5689 30636 5723 30670
rect 5757 30636 5791 30670
rect 5825 30636 5859 30670
rect 5893 30636 5927 30670
rect 5961 30636 5995 30670
rect 6029 30636 6063 30670
rect 6097 30636 6131 30670
rect 6165 30636 6199 30670
rect 6233 30636 6267 30670
rect 6301 30636 6335 30670
rect 6369 30636 6403 30670
rect 6437 30636 6471 30670
rect 6505 30636 6539 30670
rect 6573 30636 6607 30670
rect 6641 30636 6675 30670
rect 6709 30636 6743 30670
rect 6777 30636 6811 30670
rect 6845 30636 6879 30670
rect 6913 30636 6947 30670
rect 6981 30636 7015 30670
rect 7049 30636 7083 30670
rect 7117 30636 7151 30670
rect 4261 30528 4295 30562
rect 4329 30528 4363 30562
rect 4397 30528 4431 30562
rect 4465 30528 4499 30562
rect 4533 30528 4567 30562
rect 4601 30528 4635 30562
rect 4669 30528 4703 30562
rect 4737 30528 4771 30562
rect 4805 30528 4839 30562
rect 4873 30528 4907 30562
rect 4941 30528 4975 30562
rect 5009 30528 5043 30562
rect 5077 30528 5111 30562
rect 5145 30528 5179 30562
rect 5213 30528 5247 30562
rect 5281 30528 5315 30562
rect 5349 30528 5383 30562
rect 5417 30528 5451 30562
rect 5485 30528 5519 30562
rect 5553 30528 5587 30562
rect 5621 30528 5655 30562
rect 5689 30528 5723 30562
rect 5757 30528 5791 30562
rect 5825 30528 5859 30562
rect 5893 30528 5927 30562
rect 5961 30528 5995 30562
rect 6029 30528 6063 30562
rect 6097 30528 6131 30562
rect 6165 30528 6199 30562
rect 6233 30528 6267 30562
rect 6301 30528 6335 30562
rect 6369 30528 6403 30562
rect 6437 30528 6471 30562
rect 6505 30528 6539 30562
rect 6573 30528 6607 30562
rect 6641 30528 6675 30562
rect 6709 30528 6743 30562
rect 6777 30528 6811 30562
rect 6845 30528 6879 30562
rect 6913 30528 6947 30562
rect 6981 30528 7015 30562
rect 7049 30528 7083 30562
rect 7117 30528 7151 30562
rect 4144 30420 4178 30454
rect 4144 30352 4178 30386
rect 4144 30284 4178 30318
rect 4144 30216 4178 30250
rect 4144 30148 4178 30182
rect 4144 30080 4178 30114
rect 4144 30012 4178 30046
rect 4144 29944 4178 29978
rect 4144 29876 4178 29910
rect 4144 29808 4178 29842
rect 4144 29740 4178 29774
rect 4144 29672 4178 29706
rect 4144 29604 4178 29638
rect 4144 29536 4178 29570
rect -7168 29166 -4236 29200
rect 4144 29468 4178 29502
rect 4144 29400 4178 29434
rect 4144 29332 4178 29366
rect 4144 29264 4178 29298
rect 7234 30420 7268 30454
rect 7234 30352 7268 30386
rect 7234 30284 7268 30318
rect 7234 30216 7268 30250
rect 7234 30148 7268 30182
rect 7234 30080 7268 30114
rect 7234 30012 7268 30046
rect 7234 29944 7268 29978
rect 7234 29876 7268 29910
rect 7234 29808 7268 29842
rect 7234 29740 7268 29774
rect 7234 29672 7268 29706
rect 7234 29604 7268 29638
rect 7234 29536 7268 29570
rect 7234 29468 7268 29502
rect 7234 29400 7268 29434
rect 7234 29332 7268 29366
rect 7234 29264 7268 29298
rect 4261 29156 4295 29190
rect 4329 29156 4363 29190
rect 4397 29156 4431 29190
rect 4465 29156 4499 29190
rect 4533 29156 4567 29190
rect 4601 29156 4635 29190
rect 4669 29156 4703 29190
rect 4737 29156 4771 29190
rect 4805 29156 4839 29190
rect 4873 29156 4907 29190
rect 4941 29156 4975 29190
rect 5009 29156 5043 29190
rect 5077 29156 5111 29190
rect 5145 29156 5179 29190
rect 5213 29156 5247 29190
rect 5281 29156 5315 29190
rect 5349 29156 5383 29190
rect 5417 29156 5451 29190
rect 5485 29156 5519 29190
rect 5553 29156 5587 29190
rect 5621 29156 5655 29190
rect 5689 29156 5723 29190
rect 5757 29156 5791 29190
rect 5825 29156 5859 29190
rect 5893 29156 5927 29190
rect 5961 29156 5995 29190
rect 6029 29156 6063 29190
rect 6097 29156 6131 29190
rect 6165 29156 6199 29190
rect 6233 29156 6267 29190
rect 6301 29156 6335 29190
rect 6369 29156 6403 29190
rect 6437 29156 6471 29190
rect 6505 29156 6539 29190
rect 6573 29156 6607 29190
rect 6641 29156 6675 29190
rect 6709 29156 6743 29190
rect 6777 29156 6811 29190
rect 6845 29156 6879 29190
rect 6913 29156 6947 29190
rect 6981 29156 7015 29190
rect 7049 29156 7083 29190
rect 7117 29156 7151 29190
rect -562 26321 -528 26355
rect -494 26321 -460 26355
rect -426 26321 -392 26355
rect -358 26321 -324 26355
rect -290 26321 -256 26355
rect -222 26321 -188 26355
rect -154 26321 -120 26355
rect -86 26321 -52 26355
rect -18 26321 16 26355
rect 50 26321 84 26355
rect 118 26321 152 26355
rect 186 26321 220 26355
rect 254 26321 288 26355
rect 322 26321 356 26355
rect 390 26321 424 26355
rect 458 26321 492 26355
rect 526 26321 560 26355
rect -685 26208 -651 26242
rect 649 26208 683 26242
rect -685 26140 -651 26174
rect -685 26072 -651 26106
rect -685 26004 -651 26038
rect -685 25936 -651 25970
rect -685 25868 -651 25902
rect -685 25800 -651 25834
rect -685 25732 -651 25766
rect -685 25664 -651 25698
rect -685 25596 -651 25630
rect -685 25528 -651 25562
rect -685 25460 -651 25494
rect -685 25392 -651 25426
rect -685 25324 -651 25358
rect -685 25256 -651 25290
rect -685 25188 -651 25222
rect 649 26140 683 26174
rect 649 26072 683 26106
rect 649 26004 683 26038
rect 649 25936 683 25970
rect 649 25868 683 25902
rect 649 25800 683 25834
rect 649 25732 683 25766
rect 649 25664 683 25698
rect 649 25596 683 25630
rect 649 25528 683 25562
rect 649 25460 683 25494
rect 649 25392 683 25426
rect 649 25324 683 25358
rect 649 25256 683 25290
rect 649 25188 683 25222
rect -685 25120 -651 25154
rect 649 25120 683 25154
rect -562 25007 -528 25041
rect -494 25007 -460 25041
rect -426 25007 -392 25041
rect -358 25007 -324 25041
rect -290 25007 -256 25041
rect -222 25007 -188 25041
rect -154 25007 -120 25041
rect -86 25007 -52 25041
rect -18 25007 16 25041
rect 50 25007 84 25041
rect 118 25007 152 25041
rect 186 25007 220 25041
rect 254 25007 288 25041
rect 322 25007 356 25041
rect 390 25007 424 25041
rect 458 25007 492 25041
rect 526 25007 560 25041
rect -562 24801 -528 24835
rect -494 24801 -460 24835
rect -426 24801 -392 24835
rect -358 24801 -324 24835
rect -290 24801 -256 24835
rect -222 24801 -188 24835
rect -154 24801 -120 24835
rect -86 24801 -52 24835
rect -18 24801 16 24835
rect 50 24801 84 24835
rect 118 24801 152 24835
rect 186 24801 220 24835
rect 254 24801 288 24835
rect 322 24801 356 24835
rect 390 24801 424 24835
rect 458 24801 492 24835
rect 526 24801 560 24835
rect -685 24688 -651 24722
rect 649 24688 683 24722
rect -685 24620 -651 24654
rect -685 24552 -651 24586
rect -685 24484 -651 24518
rect -685 24416 -651 24450
rect -685 24348 -651 24382
rect -685 24280 -651 24314
rect -685 24212 -651 24246
rect -685 24144 -651 24178
rect -685 24076 -651 24110
rect -685 24008 -651 24042
rect -685 23940 -651 23974
rect -685 23872 -651 23906
rect -685 23804 -651 23838
rect -685 23736 -651 23770
rect -685 23668 -651 23702
rect 649 24620 683 24654
rect 649 24552 683 24586
rect 649 24484 683 24518
rect 649 24416 683 24450
rect 649 24348 683 24382
rect 649 24280 683 24314
rect 649 24212 683 24246
rect 649 24144 683 24178
rect 649 24076 683 24110
rect 649 24008 683 24042
rect 649 23940 683 23974
rect 649 23872 683 23906
rect 649 23804 683 23838
rect 649 23736 683 23770
rect 649 23668 683 23702
rect -685 23600 -651 23634
rect 649 23600 683 23634
rect -562 23487 -528 23521
rect -494 23487 -460 23521
rect -426 23487 -392 23521
rect -358 23487 -324 23521
rect -290 23487 -256 23521
rect -222 23487 -188 23521
rect -154 23487 -120 23521
rect -86 23487 -52 23521
rect -18 23487 16 23521
rect 50 23487 84 23521
rect 118 23487 152 23521
rect 186 23487 220 23521
rect 254 23487 288 23521
rect 322 23487 356 23521
rect 390 23487 424 23521
rect 458 23487 492 23521
rect 526 23487 560 23521
rect -1578 23280 -1544 23314
rect -1510 23280 -1476 23314
rect -1442 23280 -1408 23314
rect -1374 23280 -1340 23314
rect -1306 23280 -1272 23314
rect -1238 23280 -1204 23314
rect -1170 23280 -1136 23314
rect -1102 23280 -1068 23314
rect -1034 23280 -1000 23314
rect -966 23280 -932 23314
rect -898 23280 -864 23314
rect -830 23280 -796 23314
rect -762 23280 -728 23314
rect -694 23280 -660 23314
rect -626 23280 -592 23314
rect -558 23280 -524 23314
rect -490 23280 -456 23314
rect -422 23280 -388 23314
rect -354 23280 -320 23314
rect -286 23280 -252 23314
rect -218 23280 -184 23314
rect -150 23280 -116 23314
rect -82 23280 -48 23314
rect -14 23280 20 23314
rect 54 23280 88 23314
rect 122 23280 156 23314
rect 190 23280 224 23314
rect 258 23280 292 23314
rect 326 23280 360 23314
rect 394 23280 428 23314
rect 462 23280 496 23314
rect 530 23280 564 23314
rect 598 23280 632 23314
rect 666 23280 700 23314
rect 734 23280 768 23314
rect 802 23280 836 23314
rect 870 23280 904 23314
rect 938 23280 972 23314
rect 1006 23280 1040 23314
rect 1074 23280 1108 23314
rect 1142 23280 1176 23314
rect 1210 23280 1244 23314
rect 1278 23280 1312 23314
rect 1346 23280 1380 23314
rect 1414 23280 1448 23314
rect 1482 23280 1516 23314
rect 1550 23280 1584 23314
rect -1676 23167 -1642 23201
rect 1648 23167 1682 23201
rect -1676 23099 -1642 23133
rect -1676 23031 -1642 23065
rect -1676 22963 -1642 22997
rect -1676 22895 -1642 22929
rect -1676 22827 -1642 22861
rect -1676 22759 -1642 22793
rect -1676 22691 -1642 22725
rect -1676 22623 -1642 22657
rect -1676 22555 -1642 22589
rect -1676 22487 -1642 22521
rect -1676 22419 -1642 22453
rect -1676 22351 -1642 22385
rect -1676 22283 -1642 22317
rect -1676 22215 -1642 22249
rect -1676 22147 -1642 22181
rect 1648 23099 1682 23133
rect 1648 23031 1682 23065
rect 1648 22963 1682 22997
rect 1648 22895 1682 22929
rect 1648 22827 1682 22861
rect 1648 22759 1682 22793
rect 1648 22691 1682 22725
rect 1648 22623 1682 22657
rect 1648 22555 1682 22589
rect 1648 22487 1682 22521
rect 1648 22419 1682 22453
rect 1648 22351 1682 22385
rect 1648 22283 1682 22317
rect 1648 22215 1682 22249
rect 1648 22147 1682 22181
rect -1676 22079 -1642 22113
rect 1648 22079 1682 22113
rect -1578 21966 -1544 22000
rect -1510 21966 -1476 22000
rect -1442 21966 -1408 22000
rect -1374 21966 -1340 22000
rect -1306 21966 -1272 22000
rect -1238 21966 -1204 22000
rect -1170 21966 -1136 22000
rect -1102 21966 -1068 22000
rect -1034 21966 -1000 22000
rect -966 21966 -932 22000
rect -898 21966 -864 22000
rect -830 21966 -796 22000
rect -762 21966 -728 22000
rect -694 21966 -660 22000
rect -626 21966 -592 22000
rect -558 21966 -524 22000
rect -490 21966 -456 22000
rect -422 21966 -388 22000
rect -354 21966 -320 22000
rect -286 21966 -252 22000
rect -218 21966 -184 22000
rect -150 21966 -116 22000
rect -82 21966 -48 22000
rect -14 21966 20 22000
rect 54 21966 88 22000
rect 122 21966 156 22000
rect 190 21966 224 22000
rect 258 21966 292 22000
rect 326 21966 360 22000
rect 394 21966 428 22000
rect 462 21966 496 22000
rect 530 21966 564 22000
rect 598 21966 632 22000
rect 666 21966 700 22000
rect 734 21966 768 22000
rect 802 21966 836 22000
rect 870 21966 904 22000
rect 938 21966 972 22000
rect 1006 21966 1040 22000
rect 1074 21966 1108 22000
rect 1142 21966 1176 22000
rect 1210 21966 1244 22000
rect 1278 21966 1312 22000
rect 1346 21966 1380 22000
rect 1414 21966 1448 22000
rect 1482 21966 1516 22000
rect 1550 21966 1584 22000
rect -1818 21760 -1784 21794
rect -1750 21760 -1716 21794
rect -1682 21760 -1648 21794
rect -1614 21760 -1580 21794
rect -1546 21760 -1512 21794
rect -1478 21760 -1444 21794
rect -1410 21760 -1376 21794
rect -1342 21760 -1308 21794
rect -1274 21760 -1240 21794
rect -1206 21760 -1172 21794
rect -1138 21760 -1104 21794
rect -1070 21760 -1036 21794
rect -1002 21760 -968 21794
rect -934 21760 -900 21794
rect -866 21760 -832 21794
rect -798 21760 -764 21794
rect -730 21760 -696 21794
rect -662 21760 -628 21794
rect -594 21760 -560 21794
rect -526 21760 -492 21794
rect -458 21760 -424 21794
rect -390 21760 -356 21794
rect -322 21760 -288 21794
rect -254 21760 -220 21794
rect -186 21760 -152 21794
rect -118 21760 -84 21794
rect -50 21760 -16 21794
rect 18 21760 52 21794
rect 86 21760 120 21794
rect 154 21760 188 21794
rect 222 21760 256 21794
rect 290 21760 324 21794
rect 358 21760 392 21794
rect 426 21760 460 21794
rect 494 21760 528 21794
rect 562 21760 596 21794
rect 630 21760 664 21794
rect 698 21760 732 21794
rect 766 21760 800 21794
rect 834 21760 868 21794
rect 902 21760 936 21794
rect 970 21760 1004 21794
rect 1038 21760 1072 21794
rect 1106 21760 1140 21794
rect 1174 21760 1208 21794
rect 1242 21760 1276 21794
rect 1310 21760 1344 21794
rect 1378 21760 1412 21794
rect 1446 21760 1480 21794
rect 1514 21760 1548 21794
rect 1582 21760 1616 21794
rect 1650 21760 1684 21794
rect 1718 21760 1752 21794
rect 1786 21760 1820 21794
rect -1936 21647 -1902 21681
rect 1904 21647 1938 21681
rect -1936 21579 -1902 21613
rect -1936 21511 -1902 21545
rect -1936 21443 -1902 21477
rect -1936 21375 -1902 21409
rect -1936 21307 -1902 21341
rect -1936 21239 -1902 21273
rect -1936 21171 -1902 21205
rect -1936 21103 -1902 21137
rect -1936 21035 -1902 21069
rect -1936 20967 -1902 21001
rect -1936 20899 -1902 20933
rect -1936 20831 -1902 20865
rect -1936 20763 -1902 20797
rect -1936 20695 -1902 20729
rect -1936 20627 -1902 20661
rect 1904 21579 1938 21613
rect 1904 21511 1938 21545
rect 1904 21443 1938 21477
rect 1904 21375 1938 21409
rect 1904 21307 1938 21341
rect 1904 21239 1938 21273
rect 1904 21171 1938 21205
rect 1904 21103 1938 21137
rect 1904 21035 1938 21069
rect 1904 20967 1938 21001
rect 1904 20899 1938 20933
rect 1904 20831 1938 20865
rect 1904 20763 1938 20797
rect 1904 20695 1938 20729
rect 1904 20627 1938 20661
rect -1936 20559 -1902 20593
rect 1904 20559 1938 20593
rect -1818 20446 -1784 20480
rect -1750 20446 -1716 20480
rect -1682 20446 -1648 20480
rect -1614 20446 -1580 20480
rect -1546 20446 -1512 20480
rect -1478 20446 -1444 20480
rect -1410 20446 -1376 20480
rect -1342 20446 -1308 20480
rect -1274 20446 -1240 20480
rect -1206 20446 -1172 20480
rect -1138 20446 -1104 20480
rect -1070 20446 -1036 20480
rect -1002 20446 -968 20480
rect -934 20446 -900 20480
rect -866 20446 -832 20480
rect -798 20446 -764 20480
rect -730 20446 -696 20480
rect -662 20446 -628 20480
rect -594 20446 -560 20480
rect -526 20446 -492 20480
rect -458 20446 -424 20480
rect -390 20446 -356 20480
rect -322 20446 -288 20480
rect -254 20446 -220 20480
rect -186 20446 -152 20480
rect -118 20446 -84 20480
rect -50 20446 -16 20480
rect 18 20446 52 20480
rect 86 20446 120 20480
rect 154 20446 188 20480
rect 222 20446 256 20480
rect 290 20446 324 20480
rect 358 20446 392 20480
rect 426 20446 460 20480
rect 494 20446 528 20480
rect 562 20446 596 20480
rect 630 20446 664 20480
rect 698 20446 732 20480
rect 766 20446 800 20480
rect 834 20446 868 20480
rect 902 20446 936 20480
rect 970 20446 1004 20480
rect 1038 20446 1072 20480
rect 1106 20446 1140 20480
rect 1174 20446 1208 20480
rect 1242 20446 1276 20480
rect 1310 20446 1344 20480
rect 1378 20446 1412 20480
rect 1446 20446 1480 20480
rect 1514 20446 1548 20480
rect 1582 20446 1616 20480
rect 1650 20446 1684 20480
rect 1718 20446 1752 20480
rect 1786 20446 1820 20480
rect -908 18132 902 18166
rect -1004 17742 -970 18070
rect 964 17742 998 18070
rect -908 17646 902 17680
rect -688 17507 686 17541
rect -784 17217 -750 17445
rect 748 17217 782 17445
rect -688 17121 686 17155
rect -3623 16982 3623 17016
rect -3719 16592 -3685 16920
rect 3685 16592 3719 16920
rect -3623 16496 3623 16530
rect -3240 15100 -3120 15220
rect -3240 12100 -3120 12220
rect -3240 9100 -3120 9220
rect -3240 6100 -3120 6220
rect -3240 3100 -3120 3220
rect 3130 15100 3250 15220
rect 3130 12100 3250 12220
rect 3130 9100 3250 9220
rect 3130 6100 3250 6220
rect 3130 3100 3250 3220
<< nsubdiffcont >>
rect -3174 31108 -3140 31142
rect -3106 31108 -3072 31142
rect -3038 31108 -3004 31142
rect -2970 31108 -2936 31142
rect -2902 31108 -2868 31142
rect -2834 31108 -2800 31142
rect -2766 31108 -2732 31142
rect -2698 31108 -2664 31142
rect -2630 31108 -2596 31142
rect -2562 31108 -2528 31142
rect -2494 31108 -2460 31142
rect -2426 31108 -2392 31142
rect -2358 31108 -2324 31142
rect -2290 31108 -2256 31142
rect -2222 31108 -2188 31142
rect -2154 31108 -2120 31142
rect -2086 31108 -2052 31142
rect -2018 31108 -1984 31142
rect -1950 31108 -1916 31142
rect -1882 31108 -1848 31142
rect -1814 31108 -1780 31142
rect -1746 31108 -1712 31142
rect -1678 31108 -1644 31142
rect -1610 31108 -1576 31142
rect -1542 31108 -1508 31142
rect -1474 31108 -1440 31142
rect -1406 31108 -1372 31142
rect -1338 31108 -1304 31142
rect -1270 31108 -1236 31142
rect -1202 31108 -1168 31142
rect -1134 31108 -1100 31142
rect -1066 31108 -1032 31142
rect -998 31108 -964 31142
rect -930 31108 -896 31142
rect -862 31108 -828 31142
rect -794 31108 -760 31142
rect -726 31108 -692 31142
rect -658 31108 -624 31142
rect -590 31108 -556 31142
rect -522 31108 -488 31142
rect -454 31108 -420 31142
rect -386 31108 -352 31142
rect -318 31108 -284 31142
rect -250 31108 -216 31142
rect -182 31108 -148 31142
rect -114 31108 -80 31142
rect -46 31108 -12 31142
rect 22 31108 56 31142
rect 90 31108 124 31142
rect 158 31108 192 31142
rect 226 31108 260 31142
rect 294 31108 328 31142
rect 362 31108 396 31142
rect 430 31108 464 31142
rect 498 31108 532 31142
rect 566 31108 600 31142
rect 634 31108 668 31142
rect 702 31108 736 31142
rect 770 31108 804 31142
rect 838 31108 872 31142
rect 906 31108 940 31142
rect 974 31108 1008 31142
rect 1042 31108 1076 31142
rect 1110 31108 1144 31142
rect 1178 31108 1212 31142
rect 1246 31108 1280 31142
rect 1314 31108 1348 31142
rect 1382 31108 1416 31142
rect 1450 31108 1484 31142
rect 1518 31108 1552 31142
rect 1586 31108 1620 31142
rect 1654 31108 1688 31142
rect 1722 31108 1756 31142
rect 1790 31108 1824 31142
rect 1858 31108 1892 31142
rect 1926 31108 1960 31142
rect 1994 31108 2028 31142
rect 2062 31108 2096 31142
rect 2130 31108 2164 31142
rect 2198 31108 2232 31142
rect 2266 31108 2300 31142
rect 2334 31108 2368 31142
rect 2402 31108 2436 31142
rect 2470 31108 2504 31142
rect 2538 31108 2572 31142
rect 2606 31108 2640 31142
rect 2674 31108 2708 31142
rect 2742 31108 2776 31142
rect 2810 31108 2844 31142
rect 2878 31108 2912 31142
rect 2946 31108 2980 31142
rect 3014 31108 3048 31142
rect 3082 31108 3116 31142
rect 3150 31108 3184 31142
rect -3286 30986 -3252 31020
rect 3262 30986 3296 31020
rect -3286 30918 -3252 30952
rect -3286 30850 -3252 30884
rect -3286 30782 -3252 30816
rect -3286 30714 -3252 30748
rect -3286 30646 -3252 30680
rect -3286 30578 -3252 30612
rect -3286 30510 -3252 30544
rect -3286 30442 -3252 30476
rect -3286 30374 -3252 30408
rect -3286 30306 -3252 30340
rect -3286 30238 -3252 30272
rect -3286 30170 -3252 30204
rect -3286 30102 -3252 30136
rect -3286 30034 -3252 30068
rect -3286 29966 -3252 30000
rect 3262 30918 3296 30952
rect 3262 30850 3296 30884
rect 3262 30782 3296 30816
rect 3262 30714 3296 30748
rect 3262 30646 3296 30680
rect 3262 30578 3296 30612
rect 3262 30510 3296 30544
rect 3262 30442 3296 30476
rect 3262 30374 3296 30408
rect 3262 30306 3296 30340
rect 3262 30238 3296 30272
rect 3262 30170 3296 30204
rect 3262 30102 3296 30136
rect 3262 30034 3296 30068
rect 3262 29966 3296 30000
rect -3286 29898 -3252 29932
rect 3262 29898 3296 29932
rect -3174 29776 -3140 29810
rect -3106 29776 -3072 29810
rect -3038 29776 -3004 29810
rect -2970 29776 -2936 29810
rect -2902 29776 -2868 29810
rect -2834 29776 -2800 29810
rect -2766 29776 -2732 29810
rect -2698 29776 -2664 29810
rect -2630 29776 -2596 29810
rect -2562 29776 -2528 29810
rect -2494 29776 -2460 29810
rect -2426 29776 -2392 29810
rect -2358 29776 -2324 29810
rect -2290 29776 -2256 29810
rect -2222 29776 -2188 29810
rect -2154 29776 -2120 29810
rect -2086 29776 -2052 29810
rect -2018 29776 -1984 29810
rect -1950 29776 -1916 29810
rect -1882 29776 -1848 29810
rect -1814 29776 -1780 29810
rect -1746 29776 -1712 29810
rect -1678 29776 -1644 29810
rect -1610 29776 -1576 29810
rect -1542 29776 -1508 29810
rect -1474 29776 -1440 29810
rect -1406 29776 -1372 29810
rect -1338 29776 -1304 29810
rect -1270 29776 -1236 29810
rect -1202 29776 -1168 29810
rect -1134 29776 -1100 29810
rect -1066 29776 -1032 29810
rect -998 29776 -964 29810
rect -930 29776 -896 29810
rect -862 29776 -828 29810
rect -794 29776 -760 29810
rect -726 29776 -692 29810
rect -658 29776 -624 29810
rect -590 29776 -556 29810
rect -522 29776 -488 29810
rect -454 29776 -420 29810
rect -386 29776 -352 29810
rect -318 29776 -284 29810
rect -250 29776 -216 29810
rect -182 29776 -148 29810
rect -114 29776 -80 29810
rect -46 29776 -12 29810
rect 22 29776 56 29810
rect 90 29776 124 29810
rect 158 29776 192 29810
rect 226 29776 260 29810
rect 294 29776 328 29810
rect 362 29776 396 29810
rect 430 29776 464 29810
rect 498 29776 532 29810
rect 566 29776 600 29810
rect 634 29776 668 29810
rect 702 29776 736 29810
rect 770 29776 804 29810
rect 838 29776 872 29810
rect 906 29776 940 29810
rect 974 29776 1008 29810
rect 1042 29776 1076 29810
rect 1110 29776 1144 29810
rect 1178 29776 1212 29810
rect 1246 29776 1280 29810
rect 1314 29776 1348 29810
rect 1382 29776 1416 29810
rect 1450 29776 1484 29810
rect 1518 29776 1552 29810
rect 1586 29776 1620 29810
rect 1654 29776 1688 29810
rect 1722 29776 1756 29810
rect 1790 29776 1824 29810
rect 1858 29776 1892 29810
rect 1926 29776 1960 29810
rect 1994 29776 2028 29810
rect 2062 29776 2096 29810
rect 2130 29776 2164 29810
rect 2198 29776 2232 29810
rect 2266 29776 2300 29810
rect 2334 29776 2368 29810
rect 2402 29776 2436 29810
rect 2470 29776 2504 29810
rect 2538 29776 2572 29810
rect 2606 29776 2640 29810
rect 2674 29776 2708 29810
rect 2742 29776 2776 29810
rect 2810 29776 2844 29810
rect 2878 29776 2912 29810
rect 2946 29776 2980 29810
rect 3014 29776 3048 29810
rect 3082 29776 3116 29810
rect 3150 29776 3184 29810
rect -1679 29438 -1645 29472
rect -1611 29438 -1577 29472
rect -1543 29438 -1509 29472
rect -1475 29438 -1441 29472
rect -1407 29438 -1373 29472
rect -1339 29438 -1305 29472
rect -1271 29438 -1237 29472
rect -1203 29438 -1169 29472
rect -1135 29438 -1101 29472
rect -1067 29438 -1033 29472
rect -999 29438 -965 29472
rect -931 29438 -897 29472
rect -863 29438 -829 29472
rect -795 29438 -761 29472
rect -727 29438 -693 29472
rect -659 29438 -625 29472
rect -591 29438 -557 29472
rect -523 29438 -489 29472
rect -455 29438 -421 29472
rect -387 29438 -353 29472
rect -319 29438 -285 29472
rect -251 29438 -217 29472
rect -183 29438 -149 29472
rect -115 29438 -81 29472
rect -47 29438 -13 29472
rect 21 29438 55 29472
rect 89 29438 123 29472
rect 157 29438 191 29472
rect 225 29438 259 29472
rect 293 29438 327 29472
rect 361 29438 395 29472
rect 429 29438 463 29472
rect 497 29438 531 29472
rect 565 29438 599 29472
rect 633 29438 667 29472
rect 701 29438 735 29472
rect 769 29438 803 29472
rect 837 29438 871 29472
rect 905 29438 939 29472
rect 973 29438 1007 29472
rect 1041 29438 1075 29472
rect 1109 29438 1143 29472
rect 1177 29438 1211 29472
rect 1245 29438 1279 29472
rect 1313 29438 1347 29472
rect 1381 29438 1415 29472
rect 1449 29438 1483 29472
rect 1517 29438 1551 29472
rect 1585 29438 1619 29472
rect 1653 29438 1687 29472
rect -1786 29316 -1752 29350
rect 1760 29316 1794 29350
rect -1786 29248 -1752 29282
rect -1786 29180 -1752 29214
rect -1786 29112 -1752 29146
rect -1786 29044 -1752 29078
rect -1786 28976 -1752 29010
rect -1786 28908 -1752 28942
rect -1786 28840 -1752 28874
rect -1786 28772 -1752 28806
rect -1786 28704 -1752 28738
rect -1786 28636 -1752 28670
rect -1786 28568 -1752 28602
rect -1786 28500 -1752 28534
rect -1786 28432 -1752 28466
rect -1786 28364 -1752 28398
rect -1786 28296 -1752 28330
rect 1760 29248 1794 29282
rect 1760 29180 1794 29214
rect 1760 29112 1794 29146
rect 1760 29044 1794 29078
rect 1760 28976 1794 29010
rect 1760 28908 1794 28942
rect 1760 28840 1794 28874
rect 1760 28772 1794 28806
rect 1760 28704 1794 28738
rect 1760 28636 1794 28670
rect 1760 28568 1794 28602
rect 1760 28500 1794 28534
rect 1760 28432 1794 28466
rect 1760 28364 1794 28398
rect 1760 28296 1794 28330
rect -1786 28228 -1752 28262
rect 1760 28228 1794 28262
rect -1679 28106 -1645 28140
rect -1611 28106 -1577 28140
rect -1543 28106 -1509 28140
rect -1475 28106 -1441 28140
rect -1407 28106 -1373 28140
rect -1339 28106 -1305 28140
rect -1271 28106 -1237 28140
rect -1203 28106 -1169 28140
rect -1135 28106 -1101 28140
rect -1067 28106 -1033 28140
rect -999 28106 -965 28140
rect -931 28106 -897 28140
rect -863 28106 -829 28140
rect -795 28106 -761 28140
rect -727 28106 -693 28140
rect -659 28106 -625 28140
rect -591 28106 -557 28140
rect -523 28106 -489 28140
rect -455 28106 -421 28140
rect -387 28106 -353 28140
rect -319 28106 -285 28140
rect -251 28106 -217 28140
rect -183 28106 -149 28140
rect -115 28106 -81 28140
rect -47 28106 -13 28140
rect 21 28106 55 28140
rect 89 28106 123 28140
rect 157 28106 191 28140
rect 225 28106 259 28140
rect 293 28106 327 28140
rect 361 28106 395 28140
rect 429 28106 463 28140
rect 497 28106 531 28140
rect 565 28106 599 28140
rect 633 28106 667 28140
rect 701 28106 735 28140
rect 769 28106 803 28140
rect 837 28106 871 28140
rect 905 28106 939 28140
rect 973 28106 1007 28140
rect 1041 28106 1075 28140
rect 1109 28106 1143 28140
rect 1177 28106 1211 28140
rect 1245 28106 1279 28140
rect 1313 28106 1347 28140
rect 1381 28106 1415 28140
rect 1449 28106 1483 28140
rect 1517 28106 1551 28140
rect 1585 28106 1619 28140
rect 1653 28106 1687 28140
rect -1679 27898 -1645 27932
rect -1611 27898 -1577 27932
rect -1543 27898 -1509 27932
rect -1475 27898 -1441 27932
rect -1407 27898 -1373 27932
rect -1339 27898 -1305 27932
rect -1271 27898 -1237 27932
rect -1203 27898 -1169 27932
rect -1135 27898 -1101 27932
rect -1067 27898 -1033 27932
rect -999 27898 -965 27932
rect -931 27898 -897 27932
rect -863 27898 -829 27932
rect -795 27898 -761 27932
rect -727 27898 -693 27932
rect -659 27898 -625 27932
rect -591 27898 -557 27932
rect -523 27898 -489 27932
rect -455 27898 -421 27932
rect -387 27898 -353 27932
rect -319 27898 -285 27932
rect -251 27898 -217 27932
rect -183 27898 -149 27932
rect -115 27898 -81 27932
rect -47 27898 -13 27932
rect 21 27898 55 27932
rect 89 27898 123 27932
rect 157 27898 191 27932
rect 225 27898 259 27932
rect 293 27898 327 27932
rect 361 27898 395 27932
rect 429 27898 463 27932
rect 497 27898 531 27932
rect 565 27898 599 27932
rect 633 27898 667 27932
rect 701 27898 735 27932
rect 769 27898 803 27932
rect 837 27898 871 27932
rect 905 27898 939 27932
rect 973 27898 1007 27932
rect 1041 27898 1075 27932
rect 1109 27898 1143 27932
rect 1177 27898 1211 27932
rect 1245 27898 1279 27932
rect 1313 27898 1347 27932
rect 1381 27898 1415 27932
rect 1449 27898 1483 27932
rect 1517 27898 1551 27932
rect 1585 27898 1619 27932
rect 1653 27898 1687 27932
rect -1786 27776 -1752 27810
rect 1760 27776 1794 27810
rect -1786 27708 -1752 27742
rect -1786 27640 -1752 27674
rect -1786 27572 -1752 27606
rect -1786 27504 -1752 27538
rect -1786 27436 -1752 27470
rect -1786 27368 -1752 27402
rect -1786 27300 -1752 27334
rect -1786 27232 -1752 27266
rect -1786 27164 -1752 27198
rect -1786 27096 -1752 27130
rect -1786 27028 -1752 27062
rect -1786 26960 -1752 26994
rect -1786 26892 -1752 26926
rect -1786 26824 -1752 26858
rect -1786 26756 -1752 26790
rect 1760 27708 1794 27742
rect 1760 27640 1794 27674
rect 1760 27572 1794 27606
rect 1760 27504 1794 27538
rect 1760 27436 1794 27470
rect 1760 27368 1794 27402
rect 1760 27300 1794 27334
rect 1760 27232 1794 27266
rect 1760 27164 1794 27198
rect 1760 27096 1794 27130
rect 1760 27028 1794 27062
rect 1760 26960 1794 26994
rect 1760 26892 1794 26926
rect 1760 26824 1794 26858
rect 1760 26756 1794 26790
rect -1786 26688 -1752 26722
rect 1760 26688 1794 26722
rect -1679 26566 -1645 26600
rect -1611 26566 -1577 26600
rect -1543 26566 -1509 26600
rect -1475 26566 -1441 26600
rect -1407 26566 -1373 26600
rect -1339 26566 -1305 26600
rect -1271 26566 -1237 26600
rect -1203 26566 -1169 26600
rect -1135 26566 -1101 26600
rect -1067 26566 -1033 26600
rect -999 26566 -965 26600
rect -931 26566 -897 26600
rect -863 26566 -829 26600
rect -795 26566 -761 26600
rect -727 26566 -693 26600
rect -659 26566 -625 26600
rect -591 26566 -557 26600
rect -523 26566 -489 26600
rect -455 26566 -421 26600
rect -387 26566 -353 26600
rect -319 26566 -285 26600
rect -251 26566 -217 26600
rect -183 26566 -149 26600
rect -115 26566 -81 26600
rect -47 26566 -13 26600
rect 21 26566 55 26600
rect 89 26566 123 26600
rect 157 26566 191 26600
rect 225 26566 259 26600
rect 293 26566 327 26600
rect 361 26566 395 26600
rect 429 26566 463 26600
rect 497 26566 531 26600
rect 565 26566 599 26600
rect 633 26566 667 26600
rect 701 26566 735 26600
rect 769 26566 803 26600
rect 837 26566 871 26600
rect 905 26566 939 26600
rect 973 26566 1007 26600
rect 1041 26566 1075 26600
rect 1109 26566 1143 26600
rect 1177 26566 1211 26600
rect 1245 26566 1279 26600
rect 1313 26566 1347 26600
rect 1381 26566 1415 26600
rect 1449 26566 1483 26600
rect 1517 26566 1551 26600
rect 1585 26566 1619 26600
rect 1653 26566 1687 26600
rect -3678 19512 3676 19546
rect -3774 19122 -3740 19450
rect 3738 19122 3772 19450
rect -3678 19026 3676 19060
rect -3678 18922 3676 18956
rect -3774 18532 -3740 18860
rect 3738 18532 3772 18860
rect -3678 18436 3676 18470
<< poly >>
rect -3126 31040 -3026 31056
rect -3126 31006 -3093 31040
rect -3059 31006 -3026 31040
rect -3126 30959 -3026 31006
rect -2968 31040 -2868 31056
rect -2968 31006 -2935 31040
rect -2901 31006 -2868 31040
rect -2968 30959 -2868 31006
rect -2810 31040 -2710 31056
rect -2810 31006 -2777 31040
rect -2743 31006 -2710 31040
rect -2810 30959 -2710 31006
rect -2652 31040 -2552 31056
rect -2652 31006 -2619 31040
rect -2585 31006 -2552 31040
rect -2652 30959 -2552 31006
rect -2494 31040 -2394 31056
rect -2494 31006 -2461 31040
rect -2427 31006 -2394 31040
rect -2494 30959 -2394 31006
rect -2336 31040 -2236 31056
rect -2336 31006 -2303 31040
rect -2269 31006 -2236 31040
rect -2336 30959 -2236 31006
rect -2178 31040 -2078 31056
rect -2178 31006 -2145 31040
rect -2111 31006 -2078 31040
rect -2178 30959 -2078 31006
rect -2020 31040 -1920 31056
rect -2020 31006 -1987 31040
rect -1953 31006 -1920 31040
rect -2020 30959 -1920 31006
rect -1862 31040 -1762 31056
rect -1862 31006 -1829 31040
rect -1795 31006 -1762 31040
rect -1862 30959 -1762 31006
rect -1704 31040 -1604 31056
rect -1704 31006 -1671 31040
rect -1637 31006 -1604 31040
rect -1704 30959 -1604 31006
rect -1546 31040 -1446 31056
rect -1546 31006 -1513 31040
rect -1479 31006 -1446 31040
rect -1546 30959 -1446 31006
rect -1388 31040 -1288 31056
rect -1388 31006 -1355 31040
rect -1321 31006 -1288 31040
rect -1388 30959 -1288 31006
rect -1230 31040 -1130 31056
rect -1230 31006 -1197 31040
rect -1163 31006 -1130 31040
rect -1230 30959 -1130 31006
rect -1072 31040 -972 31056
rect -1072 31006 -1039 31040
rect -1005 31006 -972 31040
rect -1072 30959 -972 31006
rect -914 31040 -814 31056
rect -914 31006 -881 31040
rect -847 31006 -814 31040
rect -914 30959 -814 31006
rect -756 31040 -656 31056
rect -756 31006 -723 31040
rect -689 31006 -656 31040
rect -756 30959 -656 31006
rect -598 31040 -498 31056
rect -598 31006 -565 31040
rect -531 31006 -498 31040
rect -598 30959 -498 31006
rect -440 31040 -340 31056
rect -440 31006 -407 31040
rect -373 31006 -340 31040
rect -440 30959 -340 31006
rect -282 31040 -182 31056
rect -282 31006 -249 31040
rect -215 31006 -182 31040
rect -282 30959 -182 31006
rect -124 31040 -24 31056
rect -124 31006 -91 31040
rect -57 31006 -24 31040
rect -124 30959 -24 31006
rect 34 31040 134 31056
rect 34 31006 67 31040
rect 101 31006 134 31040
rect 34 30959 134 31006
rect 192 31040 292 31056
rect 192 31006 225 31040
rect 259 31006 292 31040
rect 192 30959 292 31006
rect 350 31040 450 31056
rect 350 31006 383 31040
rect 417 31006 450 31040
rect 350 30959 450 31006
rect 508 31040 608 31056
rect 508 31006 541 31040
rect 575 31006 608 31040
rect 508 30959 608 31006
rect 666 31040 766 31056
rect 666 31006 699 31040
rect 733 31006 766 31040
rect 666 30959 766 31006
rect 824 31040 924 31056
rect 824 31006 857 31040
rect 891 31006 924 31040
rect 824 30959 924 31006
rect 982 31040 1082 31056
rect 982 31006 1015 31040
rect 1049 31006 1082 31040
rect 982 30959 1082 31006
rect 1140 31040 1240 31056
rect 1140 31006 1173 31040
rect 1207 31006 1240 31040
rect 1140 30959 1240 31006
rect 1298 31040 1398 31056
rect 1298 31006 1331 31040
rect 1365 31006 1398 31040
rect 1298 30959 1398 31006
rect 1456 31040 1556 31056
rect 1456 31006 1489 31040
rect 1523 31006 1556 31040
rect 1456 30959 1556 31006
rect 1614 31040 1714 31056
rect 1614 31006 1647 31040
rect 1681 31006 1714 31040
rect 1614 30959 1714 31006
rect 1772 31040 1872 31056
rect 1772 31006 1805 31040
rect 1839 31006 1872 31040
rect 1772 30959 1872 31006
rect 1930 31040 2030 31056
rect 1930 31006 1963 31040
rect 1997 31006 2030 31040
rect 1930 30959 2030 31006
rect 2088 31040 2188 31056
rect 2088 31006 2121 31040
rect 2155 31006 2188 31040
rect 2088 30959 2188 31006
rect 2246 31040 2346 31056
rect 2246 31006 2279 31040
rect 2313 31006 2346 31040
rect 2246 30959 2346 31006
rect 2404 31040 2504 31056
rect 2404 31006 2437 31040
rect 2471 31006 2504 31040
rect 2404 30959 2504 31006
rect 2562 31040 2662 31056
rect 2562 31006 2595 31040
rect 2629 31006 2662 31040
rect 2562 30959 2662 31006
rect 2720 31040 2820 31056
rect 2720 31006 2753 31040
rect 2787 31006 2820 31040
rect 2720 30959 2820 31006
rect 2878 31040 2978 31056
rect 2878 31006 2911 31040
rect 2945 31006 2978 31040
rect 2878 30959 2978 31006
rect 3036 31040 3136 31056
rect 3036 31006 3069 31040
rect 3103 31006 3136 31040
rect 3036 30959 3136 31006
rect -3126 29912 -3026 29959
rect -3126 29878 -3093 29912
rect -3059 29878 -3026 29912
rect -3126 29862 -3026 29878
rect -2968 29912 -2868 29959
rect -2968 29878 -2935 29912
rect -2901 29878 -2868 29912
rect -2968 29862 -2868 29878
rect -2810 29912 -2710 29959
rect -2810 29878 -2777 29912
rect -2743 29878 -2710 29912
rect -2810 29862 -2710 29878
rect -2652 29912 -2552 29959
rect -2652 29878 -2619 29912
rect -2585 29878 -2552 29912
rect -2652 29862 -2552 29878
rect -2494 29912 -2394 29959
rect -2494 29878 -2461 29912
rect -2427 29878 -2394 29912
rect -2494 29862 -2394 29878
rect -2336 29912 -2236 29959
rect -2336 29878 -2303 29912
rect -2269 29878 -2236 29912
rect -2336 29862 -2236 29878
rect -2178 29912 -2078 29959
rect -2178 29878 -2145 29912
rect -2111 29878 -2078 29912
rect -2178 29862 -2078 29878
rect -2020 29912 -1920 29959
rect -2020 29878 -1987 29912
rect -1953 29878 -1920 29912
rect -2020 29862 -1920 29878
rect -1862 29912 -1762 29959
rect -1862 29878 -1829 29912
rect -1795 29878 -1762 29912
rect -1862 29862 -1762 29878
rect -1704 29912 -1604 29959
rect -1704 29878 -1671 29912
rect -1637 29878 -1604 29912
rect -1704 29862 -1604 29878
rect -1546 29912 -1446 29959
rect -1546 29878 -1513 29912
rect -1479 29878 -1446 29912
rect -1546 29862 -1446 29878
rect -1388 29912 -1288 29959
rect -1388 29878 -1355 29912
rect -1321 29878 -1288 29912
rect -1388 29862 -1288 29878
rect -1230 29912 -1130 29959
rect -1230 29878 -1197 29912
rect -1163 29878 -1130 29912
rect -1230 29862 -1130 29878
rect -1072 29912 -972 29959
rect -1072 29878 -1039 29912
rect -1005 29878 -972 29912
rect -1072 29862 -972 29878
rect -914 29912 -814 29959
rect -914 29878 -881 29912
rect -847 29878 -814 29912
rect -914 29862 -814 29878
rect -756 29912 -656 29959
rect -756 29878 -723 29912
rect -689 29878 -656 29912
rect -756 29862 -656 29878
rect -598 29912 -498 29959
rect -598 29878 -565 29912
rect -531 29878 -498 29912
rect -598 29862 -498 29878
rect -440 29912 -340 29959
rect -440 29878 -407 29912
rect -373 29878 -340 29912
rect -440 29862 -340 29878
rect -282 29912 -182 29959
rect -282 29878 -249 29912
rect -215 29878 -182 29912
rect -282 29862 -182 29878
rect -124 29912 -24 29959
rect -124 29878 -91 29912
rect -57 29878 -24 29912
rect -124 29862 -24 29878
rect 34 29912 134 29959
rect 34 29878 67 29912
rect 101 29878 134 29912
rect 34 29862 134 29878
rect 192 29912 292 29959
rect 192 29878 225 29912
rect 259 29878 292 29912
rect 192 29862 292 29878
rect 350 29912 450 29959
rect 350 29878 383 29912
rect 417 29878 450 29912
rect 350 29862 450 29878
rect 508 29912 608 29959
rect 508 29878 541 29912
rect 575 29878 608 29912
rect 508 29862 608 29878
rect 666 29912 766 29959
rect 666 29878 699 29912
rect 733 29878 766 29912
rect 666 29862 766 29878
rect 824 29912 924 29959
rect 824 29878 857 29912
rect 891 29878 924 29912
rect 824 29862 924 29878
rect 982 29912 1082 29959
rect 982 29878 1015 29912
rect 1049 29878 1082 29912
rect 982 29862 1082 29878
rect 1140 29912 1240 29959
rect 1140 29878 1173 29912
rect 1207 29878 1240 29912
rect 1140 29862 1240 29878
rect 1298 29912 1398 29959
rect 1298 29878 1331 29912
rect 1365 29878 1398 29912
rect 1298 29862 1398 29878
rect 1456 29912 1556 29959
rect 1456 29878 1489 29912
rect 1523 29878 1556 29912
rect 1456 29862 1556 29878
rect 1614 29912 1714 29959
rect 1614 29878 1647 29912
rect 1681 29878 1714 29912
rect 1614 29862 1714 29878
rect 1772 29912 1872 29959
rect 1772 29878 1805 29912
rect 1839 29878 1872 29912
rect 1772 29862 1872 29878
rect 1930 29912 2030 29959
rect 1930 29878 1963 29912
rect 1997 29878 2030 29912
rect 1930 29862 2030 29878
rect 2088 29912 2188 29959
rect 2088 29878 2121 29912
rect 2155 29878 2188 29912
rect 2088 29862 2188 29878
rect 2246 29912 2346 29959
rect 2246 29878 2279 29912
rect 2313 29878 2346 29912
rect 2246 29862 2346 29878
rect 2404 29912 2504 29959
rect 2404 29878 2437 29912
rect 2471 29878 2504 29912
rect 2404 29862 2504 29878
rect 2562 29912 2662 29959
rect 2562 29878 2595 29912
rect 2629 29878 2662 29912
rect 2562 29862 2662 29878
rect 2720 29912 2820 29959
rect 2720 29878 2753 29912
rect 2787 29878 2820 29912
rect 2720 29862 2820 29878
rect 2878 29912 2978 29959
rect 2878 29878 2911 29912
rect 2945 29878 2978 29912
rect 2878 29862 2978 29878
rect 3036 29912 3136 29959
rect 3036 29878 3069 29912
rect 3103 29878 3136 29912
rect 3036 29862 3136 29878
rect -1626 29370 -1526 29386
rect -1626 29336 -1593 29370
rect -1559 29336 -1526 29370
rect -1626 29289 -1526 29336
rect -1468 29370 -1368 29386
rect -1468 29336 -1435 29370
rect -1401 29336 -1368 29370
rect -1468 29289 -1368 29336
rect -1310 29370 -1210 29386
rect -1310 29336 -1277 29370
rect -1243 29336 -1210 29370
rect -1310 29289 -1210 29336
rect -1152 29370 -1052 29386
rect -1152 29336 -1119 29370
rect -1085 29336 -1052 29370
rect -1152 29289 -1052 29336
rect -994 29370 -894 29386
rect -994 29336 -961 29370
rect -927 29336 -894 29370
rect -994 29289 -894 29336
rect -836 29370 -736 29386
rect -836 29336 -803 29370
rect -769 29336 -736 29370
rect -836 29289 -736 29336
rect -678 29370 -578 29386
rect -678 29336 -645 29370
rect -611 29336 -578 29370
rect -678 29289 -578 29336
rect -520 29370 -420 29386
rect -520 29336 -487 29370
rect -453 29336 -420 29370
rect -520 29289 -420 29336
rect -362 29370 -262 29386
rect -362 29336 -329 29370
rect -295 29336 -262 29370
rect -362 29289 -262 29336
rect -204 29370 -104 29386
rect -204 29336 -171 29370
rect -137 29336 -104 29370
rect -204 29289 -104 29336
rect -46 29370 54 29386
rect -46 29336 -13 29370
rect 21 29336 54 29370
rect -46 29289 54 29336
rect 112 29370 212 29386
rect 112 29336 145 29370
rect 179 29336 212 29370
rect 112 29289 212 29336
rect 270 29370 370 29386
rect 270 29336 303 29370
rect 337 29336 370 29370
rect 270 29289 370 29336
rect 428 29370 528 29386
rect 428 29336 461 29370
rect 495 29336 528 29370
rect 428 29289 528 29336
rect 586 29370 686 29386
rect 586 29336 619 29370
rect 653 29336 686 29370
rect 586 29289 686 29336
rect 744 29370 844 29386
rect 744 29336 777 29370
rect 811 29336 844 29370
rect 744 29289 844 29336
rect 902 29370 1002 29386
rect 902 29336 935 29370
rect 969 29336 1002 29370
rect 902 29289 1002 29336
rect 1060 29370 1160 29386
rect 1060 29336 1093 29370
rect 1127 29336 1160 29370
rect 1060 29289 1160 29336
rect 1218 29370 1318 29386
rect 1218 29336 1251 29370
rect 1285 29336 1318 29370
rect 1218 29289 1318 29336
rect 1376 29370 1476 29386
rect 1376 29336 1409 29370
rect 1443 29336 1476 29370
rect 1376 29289 1476 29336
rect 1534 29370 1634 29386
rect 1534 29336 1567 29370
rect 1601 29336 1634 29370
rect 1534 29289 1634 29336
rect -1626 28242 -1526 28289
rect -1626 28208 -1593 28242
rect -1559 28208 -1526 28242
rect -1626 28192 -1526 28208
rect -1468 28242 -1368 28289
rect -1468 28208 -1435 28242
rect -1401 28208 -1368 28242
rect -1468 28192 -1368 28208
rect -1310 28242 -1210 28289
rect -1310 28208 -1277 28242
rect -1243 28208 -1210 28242
rect -1310 28192 -1210 28208
rect -1152 28242 -1052 28289
rect -1152 28208 -1119 28242
rect -1085 28208 -1052 28242
rect -1152 28192 -1052 28208
rect -994 28242 -894 28289
rect -994 28208 -961 28242
rect -927 28208 -894 28242
rect -994 28192 -894 28208
rect -836 28242 -736 28289
rect -836 28208 -803 28242
rect -769 28208 -736 28242
rect -836 28192 -736 28208
rect -678 28242 -578 28289
rect -678 28208 -645 28242
rect -611 28208 -578 28242
rect -678 28192 -578 28208
rect -520 28242 -420 28289
rect -520 28208 -487 28242
rect -453 28208 -420 28242
rect -520 28192 -420 28208
rect -362 28242 -262 28289
rect -362 28208 -329 28242
rect -295 28208 -262 28242
rect -362 28192 -262 28208
rect -204 28242 -104 28289
rect -204 28208 -171 28242
rect -137 28208 -104 28242
rect -204 28192 -104 28208
rect -46 28242 54 28289
rect -46 28208 -13 28242
rect 21 28208 54 28242
rect -46 28192 54 28208
rect 112 28242 212 28289
rect 112 28208 145 28242
rect 179 28208 212 28242
rect 112 28192 212 28208
rect 270 28242 370 28289
rect 270 28208 303 28242
rect 337 28208 370 28242
rect 270 28192 370 28208
rect 428 28242 528 28289
rect 428 28208 461 28242
rect 495 28208 528 28242
rect 428 28192 528 28208
rect 586 28242 686 28289
rect 586 28208 619 28242
rect 653 28208 686 28242
rect 586 28192 686 28208
rect 744 28242 844 28289
rect 744 28208 777 28242
rect 811 28208 844 28242
rect 744 28192 844 28208
rect 902 28242 1002 28289
rect 902 28208 935 28242
rect 969 28208 1002 28242
rect 902 28192 1002 28208
rect 1060 28242 1160 28289
rect 1060 28208 1093 28242
rect 1127 28208 1160 28242
rect 1060 28192 1160 28208
rect 1218 28242 1318 28289
rect 1218 28208 1251 28242
rect 1285 28208 1318 28242
rect 1218 28192 1318 28208
rect 1376 28242 1476 28289
rect 1376 28208 1409 28242
rect 1443 28208 1476 28242
rect 1376 28192 1476 28208
rect 1534 28242 1634 28289
rect 1534 28208 1567 28242
rect 1601 28208 1634 28242
rect 1534 28192 1634 28208
rect -1626 27830 -1526 27846
rect -1626 27796 -1593 27830
rect -1559 27796 -1526 27830
rect -1626 27749 -1526 27796
rect -1468 27830 -1368 27846
rect -1468 27796 -1435 27830
rect -1401 27796 -1368 27830
rect -1468 27749 -1368 27796
rect -1310 27830 -1210 27846
rect -1310 27796 -1277 27830
rect -1243 27796 -1210 27830
rect -1310 27749 -1210 27796
rect -1152 27830 -1052 27846
rect -1152 27796 -1119 27830
rect -1085 27796 -1052 27830
rect -1152 27749 -1052 27796
rect -994 27830 -894 27846
rect -994 27796 -961 27830
rect -927 27796 -894 27830
rect -994 27749 -894 27796
rect -836 27830 -736 27846
rect -836 27796 -803 27830
rect -769 27796 -736 27830
rect -836 27749 -736 27796
rect -678 27830 -578 27846
rect -678 27796 -645 27830
rect -611 27796 -578 27830
rect -678 27749 -578 27796
rect -520 27830 -420 27846
rect -520 27796 -487 27830
rect -453 27796 -420 27830
rect -520 27749 -420 27796
rect -362 27830 -262 27846
rect -362 27796 -329 27830
rect -295 27796 -262 27830
rect -362 27749 -262 27796
rect -204 27830 -104 27846
rect -204 27796 -171 27830
rect -137 27796 -104 27830
rect -204 27749 -104 27796
rect -46 27830 54 27846
rect -46 27796 -13 27830
rect 21 27796 54 27830
rect -46 27749 54 27796
rect 112 27830 212 27846
rect 112 27796 145 27830
rect 179 27796 212 27830
rect 112 27749 212 27796
rect 270 27830 370 27846
rect 270 27796 303 27830
rect 337 27796 370 27830
rect 270 27749 370 27796
rect 428 27830 528 27846
rect 428 27796 461 27830
rect 495 27796 528 27830
rect 428 27749 528 27796
rect 586 27830 686 27846
rect 586 27796 619 27830
rect 653 27796 686 27830
rect 586 27749 686 27796
rect 744 27830 844 27846
rect 744 27796 777 27830
rect 811 27796 844 27830
rect 744 27749 844 27796
rect 902 27830 1002 27846
rect 902 27796 935 27830
rect 969 27796 1002 27830
rect 902 27749 1002 27796
rect 1060 27830 1160 27846
rect 1060 27796 1093 27830
rect 1127 27796 1160 27830
rect 1060 27749 1160 27796
rect 1218 27830 1318 27846
rect 1218 27796 1251 27830
rect 1285 27796 1318 27830
rect 1218 27749 1318 27796
rect 1376 27830 1476 27846
rect 1376 27796 1409 27830
rect 1443 27796 1476 27830
rect 1376 27749 1476 27796
rect 1534 27830 1634 27846
rect 1534 27796 1567 27830
rect 1601 27796 1634 27830
rect 1534 27749 1634 27796
rect -1626 26702 -1526 26749
rect -1626 26668 -1593 26702
rect -1559 26668 -1526 26702
rect -1626 26652 -1526 26668
rect -1468 26702 -1368 26749
rect -1468 26668 -1435 26702
rect -1401 26668 -1368 26702
rect -1468 26652 -1368 26668
rect -1310 26702 -1210 26749
rect -1310 26668 -1277 26702
rect -1243 26668 -1210 26702
rect -1310 26652 -1210 26668
rect -1152 26702 -1052 26749
rect -1152 26668 -1119 26702
rect -1085 26668 -1052 26702
rect -1152 26652 -1052 26668
rect -994 26702 -894 26749
rect -994 26668 -961 26702
rect -927 26668 -894 26702
rect -994 26652 -894 26668
rect -836 26702 -736 26749
rect -836 26668 -803 26702
rect -769 26668 -736 26702
rect -836 26652 -736 26668
rect -678 26702 -578 26749
rect -678 26668 -645 26702
rect -611 26668 -578 26702
rect -678 26652 -578 26668
rect -520 26702 -420 26749
rect -520 26668 -487 26702
rect -453 26668 -420 26702
rect -520 26652 -420 26668
rect -362 26702 -262 26749
rect -362 26668 -329 26702
rect -295 26668 -262 26702
rect -362 26652 -262 26668
rect -204 26702 -104 26749
rect -204 26668 -171 26702
rect -137 26668 -104 26702
rect -204 26652 -104 26668
rect -46 26702 54 26749
rect -46 26668 -13 26702
rect 21 26668 54 26702
rect -46 26652 54 26668
rect 112 26702 212 26749
rect 112 26668 145 26702
rect 179 26668 212 26702
rect 112 26652 212 26668
rect 270 26702 370 26749
rect 270 26668 303 26702
rect 337 26668 370 26702
rect 270 26652 370 26668
rect 428 26702 528 26749
rect 428 26668 461 26702
rect 495 26668 528 26702
rect 428 26652 528 26668
rect 586 26702 686 26749
rect 586 26668 619 26702
rect 653 26668 686 26702
rect 586 26652 686 26668
rect 744 26702 844 26749
rect 744 26668 777 26702
rect 811 26668 844 26702
rect 744 26652 844 26668
rect 902 26702 1002 26749
rect 902 26668 935 26702
rect 969 26668 1002 26702
rect 902 26652 1002 26668
rect 1060 26702 1160 26749
rect 1060 26668 1093 26702
rect 1127 26668 1160 26702
rect 1060 26652 1160 26668
rect 1218 26702 1318 26749
rect 1218 26668 1251 26702
rect 1285 26668 1318 26702
rect 1218 26652 1318 26668
rect 1376 26702 1476 26749
rect 1376 26668 1409 26702
rect 1443 26668 1476 26702
rect 1376 26652 1476 26668
rect 1534 26702 1634 26749
rect 1534 26668 1567 26702
rect 1601 26668 1634 26702
rect 1534 26652 1634 26668
rect -525 26253 -425 26269
rect -525 26219 -492 26253
rect -458 26219 -425 26253
rect -525 26181 -425 26219
rect -367 26253 -267 26269
rect -367 26219 -334 26253
rect -300 26219 -267 26253
rect -367 26181 -267 26219
rect -209 26253 -109 26269
rect -209 26219 -176 26253
rect -142 26219 -109 26253
rect -209 26181 -109 26219
rect -51 26253 49 26269
rect -51 26219 -18 26253
rect 16 26219 49 26253
rect -51 26181 49 26219
rect 107 26253 207 26269
rect 107 26219 140 26253
rect 174 26219 207 26253
rect 107 26181 207 26219
rect 265 26253 365 26269
rect 265 26219 298 26253
rect 332 26219 365 26253
rect 265 26181 365 26219
rect 423 26253 523 26269
rect 423 26219 456 26253
rect 490 26219 523 26253
rect 423 26181 523 26219
rect -525 25143 -425 25181
rect -525 25109 -492 25143
rect -458 25109 -425 25143
rect -525 25093 -425 25109
rect -367 25143 -267 25181
rect -367 25109 -334 25143
rect -300 25109 -267 25143
rect -367 25093 -267 25109
rect -209 25143 -109 25181
rect -209 25109 -176 25143
rect -142 25109 -109 25143
rect -209 25093 -109 25109
rect -51 25143 49 25181
rect -51 25109 -18 25143
rect 16 25109 49 25143
rect -51 25093 49 25109
rect 107 25143 207 25181
rect 107 25109 140 25143
rect 174 25109 207 25143
rect 107 25093 207 25109
rect 265 25143 365 25181
rect 265 25109 298 25143
rect 332 25109 365 25143
rect 265 25093 365 25109
rect 423 25143 523 25181
rect 423 25109 456 25143
rect 490 25109 523 25143
rect 423 25093 523 25109
rect -525 24733 -425 24749
rect -525 24699 -492 24733
rect -458 24699 -425 24733
rect -525 24661 -425 24699
rect -367 24733 -267 24749
rect -367 24699 -334 24733
rect -300 24699 -267 24733
rect -367 24661 -267 24699
rect -209 24733 -109 24749
rect -209 24699 -176 24733
rect -142 24699 -109 24733
rect -209 24661 -109 24699
rect -51 24733 49 24749
rect -51 24699 -18 24733
rect 16 24699 49 24733
rect -51 24661 49 24699
rect 107 24733 207 24749
rect 107 24699 140 24733
rect 174 24699 207 24733
rect 107 24661 207 24699
rect 265 24733 365 24749
rect 265 24699 298 24733
rect 332 24699 365 24733
rect 265 24661 365 24699
rect 423 24733 523 24749
rect 423 24699 456 24733
rect 490 24699 523 24733
rect 423 24661 523 24699
rect -525 23623 -425 23661
rect -525 23589 -492 23623
rect -458 23589 -425 23623
rect -525 23573 -425 23589
rect -367 23623 -267 23661
rect -367 23589 -334 23623
rect -300 23589 -267 23623
rect -367 23573 -267 23589
rect -209 23623 -109 23661
rect -209 23589 -176 23623
rect -142 23589 -109 23623
rect -209 23573 -109 23589
rect -51 23623 49 23661
rect -51 23589 -18 23623
rect 16 23589 49 23623
rect -51 23573 49 23589
rect 107 23623 207 23661
rect 107 23589 140 23623
rect 174 23589 207 23623
rect 107 23573 207 23589
rect 265 23623 365 23661
rect 265 23589 298 23623
rect 332 23589 365 23623
rect 265 23573 365 23589
rect 423 23623 523 23661
rect 423 23589 456 23623
rect 490 23589 523 23623
rect 423 23573 523 23589
rect -1516 23212 -1316 23228
rect -1516 23178 -1467 23212
rect -1433 23178 -1399 23212
rect -1365 23178 -1316 23212
rect -1516 23140 -1316 23178
rect -1258 23212 -1058 23228
rect -1258 23178 -1209 23212
rect -1175 23178 -1141 23212
rect -1107 23178 -1058 23212
rect -1258 23140 -1058 23178
rect -1000 23212 -800 23228
rect -1000 23178 -951 23212
rect -917 23178 -883 23212
rect -849 23178 -800 23212
rect -1000 23140 -800 23178
rect -742 23212 -542 23228
rect -742 23178 -693 23212
rect -659 23178 -625 23212
rect -591 23178 -542 23212
rect -742 23140 -542 23178
rect -484 23212 -284 23228
rect -484 23178 -435 23212
rect -401 23178 -367 23212
rect -333 23178 -284 23212
rect -484 23140 -284 23178
rect -226 23212 -26 23228
rect -226 23178 -177 23212
rect -143 23178 -109 23212
rect -75 23178 -26 23212
rect -226 23140 -26 23178
rect 32 23212 232 23228
rect 32 23178 81 23212
rect 115 23178 149 23212
rect 183 23178 232 23212
rect 32 23140 232 23178
rect 290 23212 490 23228
rect 290 23178 339 23212
rect 373 23178 407 23212
rect 441 23178 490 23212
rect 290 23140 490 23178
rect 548 23212 748 23228
rect 548 23178 597 23212
rect 631 23178 665 23212
rect 699 23178 748 23212
rect 548 23140 748 23178
rect 806 23212 1006 23228
rect 806 23178 855 23212
rect 889 23178 923 23212
rect 957 23178 1006 23212
rect 806 23140 1006 23178
rect 1064 23212 1264 23228
rect 1064 23178 1113 23212
rect 1147 23178 1181 23212
rect 1215 23178 1264 23212
rect 1064 23140 1264 23178
rect 1322 23212 1522 23228
rect 1322 23178 1371 23212
rect 1405 23178 1439 23212
rect 1473 23178 1522 23212
rect 1322 23140 1522 23178
rect -1516 22102 -1316 22140
rect -1516 22068 -1467 22102
rect -1433 22068 -1399 22102
rect -1365 22068 -1316 22102
rect -1516 22052 -1316 22068
rect -1258 22102 -1058 22140
rect -1258 22068 -1209 22102
rect -1175 22068 -1141 22102
rect -1107 22068 -1058 22102
rect -1258 22052 -1058 22068
rect -1000 22102 -800 22140
rect -1000 22068 -951 22102
rect -917 22068 -883 22102
rect -849 22068 -800 22102
rect -1000 22052 -800 22068
rect -742 22102 -542 22140
rect -742 22068 -693 22102
rect -659 22068 -625 22102
rect -591 22068 -542 22102
rect -742 22052 -542 22068
rect -484 22102 -284 22140
rect -484 22068 -435 22102
rect -401 22068 -367 22102
rect -333 22068 -284 22102
rect -484 22052 -284 22068
rect -226 22102 -26 22140
rect -226 22068 -177 22102
rect -143 22068 -109 22102
rect -75 22068 -26 22102
rect -226 22052 -26 22068
rect 32 22102 232 22140
rect 32 22068 81 22102
rect 115 22068 149 22102
rect 183 22068 232 22102
rect 32 22052 232 22068
rect 290 22102 490 22140
rect 290 22068 339 22102
rect 373 22068 407 22102
rect 441 22068 490 22102
rect 290 22052 490 22068
rect 548 22102 748 22140
rect 548 22068 597 22102
rect 631 22068 665 22102
rect 699 22068 748 22102
rect 548 22052 748 22068
rect 806 22102 1006 22140
rect 806 22068 855 22102
rect 889 22068 923 22102
rect 957 22068 1006 22102
rect 806 22052 1006 22068
rect 1064 22102 1264 22140
rect 1064 22068 1113 22102
rect 1147 22068 1181 22102
rect 1215 22068 1264 22102
rect 1064 22052 1264 22068
rect 1322 22102 1522 22140
rect 1322 22068 1371 22102
rect 1405 22068 1439 22102
rect 1473 22068 1522 22102
rect 1322 22052 1522 22068
rect -1776 21692 -1576 21708
rect -1776 21658 -1727 21692
rect -1693 21658 -1659 21692
rect -1625 21658 -1576 21692
rect -1776 21620 -1576 21658
rect -1518 21692 -1318 21708
rect -1518 21658 -1469 21692
rect -1435 21658 -1401 21692
rect -1367 21658 -1318 21692
rect -1518 21620 -1318 21658
rect -1260 21692 -1060 21708
rect -1260 21658 -1211 21692
rect -1177 21658 -1143 21692
rect -1109 21658 -1060 21692
rect -1260 21620 -1060 21658
rect -1002 21692 -802 21708
rect -1002 21658 -953 21692
rect -919 21658 -885 21692
rect -851 21658 -802 21692
rect -1002 21620 -802 21658
rect -744 21692 -544 21708
rect -744 21658 -695 21692
rect -661 21658 -627 21692
rect -593 21658 -544 21692
rect -744 21620 -544 21658
rect -486 21692 -286 21708
rect -486 21658 -437 21692
rect -403 21658 -369 21692
rect -335 21658 -286 21692
rect -486 21620 -286 21658
rect -228 21692 -28 21708
rect -228 21658 -179 21692
rect -145 21658 -111 21692
rect -77 21658 -28 21692
rect -228 21620 -28 21658
rect 30 21692 230 21708
rect 30 21658 79 21692
rect 113 21658 147 21692
rect 181 21658 230 21692
rect 30 21620 230 21658
rect 288 21692 488 21708
rect 288 21658 337 21692
rect 371 21658 405 21692
rect 439 21658 488 21692
rect 288 21620 488 21658
rect 546 21692 746 21708
rect 546 21658 595 21692
rect 629 21658 663 21692
rect 697 21658 746 21692
rect 546 21620 746 21658
rect 804 21692 1004 21708
rect 804 21658 853 21692
rect 887 21658 921 21692
rect 955 21658 1004 21692
rect 804 21620 1004 21658
rect 1062 21692 1262 21708
rect 1062 21658 1111 21692
rect 1145 21658 1179 21692
rect 1213 21658 1262 21692
rect 1062 21620 1262 21658
rect 1320 21692 1520 21708
rect 1320 21658 1369 21692
rect 1403 21658 1437 21692
rect 1471 21658 1520 21692
rect 1320 21620 1520 21658
rect 1578 21692 1778 21708
rect 1578 21658 1627 21692
rect 1661 21658 1695 21692
rect 1729 21658 1778 21692
rect 1578 21620 1778 21658
rect -1776 20582 -1576 20620
rect -1776 20548 -1727 20582
rect -1693 20548 -1659 20582
rect -1625 20548 -1576 20582
rect -1776 20532 -1576 20548
rect -1518 20582 -1318 20620
rect -1518 20548 -1469 20582
rect -1435 20548 -1401 20582
rect -1367 20548 -1318 20582
rect -1518 20532 -1318 20548
rect -1260 20582 -1060 20620
rect -1260 20548 -1211 20582
rect -1177 20548 -1143 20582
rect -1109 20548 -1060 20582
rect -1260 20532 -1060 20548
rect -1002 20582 -802 20620
rect -1002 20548 -953 20582
rect -919 20548 -885 20582
rect -851 20548 -802 20582
rect -1002 20532 -802 20548
rect -744 20582 -544 20620
rect -744 20548 -695 20582
rect -661 20548 -627 20582
rect -593 20548 -544 20582
rect -744 20532 -544 20548
rect -486 20582 -286 20620
rect -486 20548 -437 20582
rect -403 20548 -369 20582
rect -335 20548 -286 20582
rect -486 20532 -286 20548
rect -228 20582 -28 20620
rect -228 20548 -179 20582
rect -145 20548 -111 20582
rect -77 20548 -28 20582
rect -228 20532 -28 20548
rect 30 20582 230 20620
rect 30 20548 79 20582
rect 113 20548 147 20582
rect 181 20548 230 20582
rect 30 20532 230 20548
rect 288 20582 488 20620
rect 288 20548 337 20582
rect 371 20548 405 20582
rect 439 20548 488 20582
rect 288 20532 488 20548
rect 546 20582 746 20620
rect 546 20548 595 20582
rect 629 20548 663 20582
rect 697 20548 746 20582
rect 546 20532 746 20548
rect 804 20582 1004 20620
rect 804 20548 853 20582
rect 887 20548 921 20582
rect 955 20548 1004 20582
rect 804 20532 1004 20548
rect 1062 20582 1262 20620
rect 1062 20548 1111 20582
rect 1145 20548 1179 20582
rect 1213 20548 1262 20582
rect 1062 20532 1262 20548
rect 1320 20582 1520 20620
rect 1320 20548 1369 20582
rect 1403 20548 1437 20582
rect 1471 20548 1520 20582
rect 1320 20532 1520 20548
rect 1578 20582 1778 20620
rect 1578 20548 1627 20582
rect 1661 20548 1695 20582
rect 1729 20548 1778 20582
rect 1578 20532 1778 20548
rect -3688 19370 -3591 19386
rect -3688 19202 -3672 19370
rect -3638 19202 -3591 19370
rect -3688 19186 -3591 19202
rect -2591 19370 -2494 19386
rect -2591 19202 -2544 19370
rect -2510 19202 -2494 19370
rect -2591 19186 -2494 19202
rect -2452 19370 -2355 19386
rect -2452 19202 -2436 19370
rect -2402 19202 -2355 19370
rect -2452 19186 -2355 19202
rect -1355 19370 -1258 19386
rect -1355 19202 -1308 19370
rect -1274 19202 -1258 19370
rect -1355 19186 -1258 19202
rect -1216 19370 -1119 19386
rect -1216 19202 -1200 19370
rect -1166 19202 -1119 19370
rect -1216 19186 -1119 19202
rect -119 19370 -22 19386
rect -119 19202 -72 19370
rect -38 19202 -22 19370
rect -119 19186 -22 19202
rect 20 19370 117 19386
rect 20 19202 36 19370
rect 70 19202 117 19370
rect 20 19186 117 19202
rect 1117 19370 1214 19386
rect 1117 19202 1164 19370
rect 1198 19202 1214 19370
rect 1117 19186 1214 19202
rect 1256 19370 1353 19386
rect 1256 19202 1272 19370
rect 1306 19202 1353 19370
rect 1256 19186 1353 19202
rect 2353 19370 2450 19386
rect 2353 19202 2400 19370
rect 2434 19202 2450 19370
rect 2353 19186 2450 19202
rect 2492 19370 2589 19386
rect 2492 19202 2508 19370
rect 2542 19202 2589 19370
rect 2492 19186 2589 19202
rect 3589 19370 3686 19386
rect 3589 19202 3636 19370
rect 3670 19202 3686 19370
rect 3589 19186 3686 19202
rect -3688 18780 -3591 18796
rect -3688 18612 -3672 18780
rect -3638 18612 -3591 18780
rect -3688 18596 -3591 18612
rect -2591 18780 -2494 18796
rect -2591 18612 -2544 18780
rect -2510 18612 -2494 18780
rect -2591 18596 -2494 18612
rect -2452 18780 -2355 18796
rect -2452 18612 -2436 18780
rect -2402 18612 -2355 18780
rect -2452 18596 -2355 18612
rect -1355 18780 -1258 18796
rect -1355 18612 -1308 18780
rect -1274 18612 -1258 18780
rect -1355 18596 -1258 18612
rect -1216 18780 -1119 18796
rect -1216 18612 -1200 18780
rect -1166 18612 -1119 18780
rect -1216 18596 -1119 18612
rect -119 18780 -22 18796
rect -119 18612 -72 18780
rect -38 18612 -22 18780
rect -119 18596 -22 18612
rect 20 18780 117 18796
rect 20 18612 36 18780
rect 70 18612 117 18780
rect 20 18596 117 18612
rect 1117 18780 1214 18796
rect 1117 18612 1164 18780
rect 1198 18612 1214 18780
rect 1117 18596 1214 18612
rect 1256 18780 1353 18796
rect 1256 18612 1272 18780
rect 1306 18612 1353 18780
rect 1256 18596 1353 18612
rect 2353 18780 2450 18796
rect 2353 18612 2400 18780
rect 2434 18612 2450 18780
rect 2353 18596 2450 18612
rect 2492 18780 2589 18796
rect 2492 18612 2508 18780
rect 2542 18612 2589 18780
rect 2492 18596 2589 18612
rect 3589 18780 3686 18796
rect 3589 18612 3636 18780
rect 3670 18612 3686 18780
rect 3589 18596 3686 18612
rect -918 17990 -830 18006
rect -918 17822 -902 17990
rect -868 17822 -830 17990
rect -918 17806 -830 17822
rect -580 17990 -492 18006
rect -580 17822 -542 17990
rect -508 17822 -492 17990
rect -580 17806 -492 17822
rect -450 17990 -362 18006
rect -450 17822 -434 17990
rect -400 17822 -362 17990
rect -450 17806 -362 17822
rect -112 17990 -24 18006
rect -112 17822 -74 17990
rect -40 17822 -24 17990
rect -112 17806 -24 17822
rect 18 17990 106 18006
rect 18 17822 34 17990
rect 68 17822 106 17990
rect 18 17806 106 17822
rect 356 17990 444 18006
rect 356 17822 394 17990
rect 428 17822 444 17990
rect 356 17806 444 17822
rect 486 17990 574 18006
rect 486 17822 502 17990
rect 536 17822 574 17990
rect 486 17806 574 17822
rect 824 17990 912 18006
rect 824 17822 862 17990
rect 896 17822 912 17990
rect 824 17806 912 17822
rect -698 17365 -610 17381
rect -698 17297 -682 17365
rect -648 17297 -610 17365
rect -698 17281 -610 17297
rect -110 17365 -22 17381
rect -110 17297 -72 17365
rect -38 17297 -22 17365
rect -110 17281 -22 17297
rect 20 17365 108 17381
rect 20 17297 36 17365
rect 70 17297 108 17365
rect 20 17281 108 17297
rect 608 17365 696 17381
rect 608 17297 646 17365
rect 680 17297 696 17365
rect 608 17281 696 17297
rect -3633 16840 -3545 16856
rect -3633 16672 -3617 16840
rect -3583 16672 -3545 16840
rect -3633 16656 -3545 16672
rect -2545 16840 -2457 16856
rect -2545 16672 -2507 16840
rect -2473 16672 -2457 16840
rect -2545 16656 -2457 16672
rect -2415 16840 -2327 16856
rect -2415 16672 -2399 16840
rect -2365 16672 -2327 16840
rect -2415 16656 -2327 16672
rect -1327 16840 -1239 16856
rect -1327 16672 -1289 16840
rect -1255 16672 -1239 16840
rect -1327 16656 -1239 16672
rect -1197 16840 -1109 16856
rect -1197 16672 -1181 16840
rect -1147 16672 -1109 16840
rect -1197 16656 -1109 16672
rect -109 16840 -21 16856
rect -109 16672 -71 16840
rect -37 16672 -21 16840
rect -109 16656 -21 16672
rect 21 16840 109 16856
rect 21 16672 37 16840
rect 71 16672 109 16840
rect 21 16656 109 16672
rect 1109 16840 1197 16856
rect 1109 16672 1147 16840
rect 1181 16672 1197 16840
rect 1109 16656 1197 16672
rect 1239 16840 1327 16856
rect 1239 16672 1255 16840
rect 1289 16672 1327 16840
rect 1239 16656 1327 16672
rect 2327 16840 2415 16856
rect 2327 16672 2365 16840
rect 2399 16672 2415 16840
rect 2327 16656 2415 16672
rect 2457 16840 2545 16856
rect 2457 16672 2473 16840
rect 2507 16672 2545 16840
rect 2457 16656 2545 16672
rect 3545 16840 3633 16856
rect 3545 16672 3583 16840
rect 3617 16672 3633 16840
rect 3545 16656 3633 16672
<< polycont >>
rect -3093 31006 -3059 31040
rect -2935 31006 -2901 31040
rect -2777 31006 -2743 31040
rect -2619 31006 -2585 31040
rect -2461 31006 -2427 31040
rect -2303 31006 -2269 31040
rect -2145 31006 -2111 31040
rect -1987 31006 -1953 31040
rect -1829 31006 -1795 31040
rect -1671 31006 -1637 31040
rect -1513 31006 -1479 31040
rect -1355 31006 -1321 31040
rect -1197 31006 -1163 31040
rect -1039 31006 -1005 31040
rect -881 31006 -847 31040
rect -723 31006 -689 31040
rect -565 31006 -531 31040
rect -407 31006 -373 31040
rect -249 31006 -215 31040
rect -91 31006 -57 31040
rect 67 31006 101 31040
rect 225 31006 259 31040
rect 383 31006 417 31040
rect 541 31006 575 31040
rect 699 31006 733 31040
rect 857 31006 891 31040
rect 1015 31006 1049 31040
rect 1173 31006 1207 31040
rect 1331 31006 1365 31040
rect 1489 31006 1523 31040
rect 1647 31006 1681 31040
rect 1805 31006 1839 31040
rect 1963 31006 1997 31040
rect 2121 31006 2155 31040
rect 2279 31006 2313 31040
rect 2437 31006 2471 31040
rect 2595 31006 2629 31040
rect 2753 31006 2787 31040
rect 2911 31006 2945 31040
rect 3069 31006 3103 31040
rect -3093 29878 -3059 29912
rect -2935 29878 -2901 29912
rect -2777 29878 -2743 29912
rect -2619 29878 -2585 29912
rect -2461 29878 -2427 29912
rect -2303 29878 -2269 29912
rect -2145 29878 -2111 29912
rect -1987 29878 -1953 29912
rect -1829 29878 -1795 29912
rect -1671 29878 -1637 29912
rect -1513 29878 -1479 29912
rect -1355 29878 -1321 29912
rect -1197 29878 -1163 29912
rect -1039 29878 -1005 29912
rect -881 29878 -847 29912
rect -723 29878 -689 29912
rect -565 29878 -531 29912
rect -407 29878 -373 29912
rect -249 29878 -215 29912
rect -91 29878 -57 29912
rect 67 29878 101 29912
rect 225 29878 259 29912
rect 383 29878 417 29912
rect 541 29878 575 29912
rect 699 29878 733 29912
rect 857 29878 891 29912
rect 1015 29878 1049 29912
rect 1173 29878 1207 29912
rect 1331 29878 1365 29912
rect 1489 29878 1523 29912
rect 1647 29878 1681 29912
rect 1805 29878 1839 29912
rect 1963 29878 1997 29912
rect 2121 29878 2155 29912
rect 2279 29878 2313 29912
rect 2437 29878 2471 29912
rect 2595 29878 2629 29912
rect 2753 29878 2787 29912
rect 2911 29878 2945 29912
rect 3069 29878 3103 29912
rect -1593 29336 -1559 29370
rect -1435 29336 -1401 29370
rect -1277 29336 -1243 29370
rect -1119 29336 -1085 29370
rect -961 29336 -927 29370
rect -803 29336 -769 29370
rect -645 29336 -611 29370
rect -487 29336 -453 29370
rect -329 29336 -295 29370
rect -171 29336 -137 29370
rect -13 29336 21 29370
rect 145 29336 179 29370
rect 303 29336 337 29370
rect 461 29336 495 29370
rect 619 29336 653 29370
rect 777 29336 811 29370
rect 935 29336 969 29370
rect 1093 29336 1127 29370
rect 1251 29336 1285 29370
rect 1409 29336 1443 29370
rect 1567 29336 1601 29370
rect -1593 28208 -1559 28242
rect -1435 28208 -1401 28242
rect -1277 28208 -1243 28242
rect -1119 28208 -1085 28242
rect -961 28208 -927 28242
rect -803 28208 -769 28242
rect -645 28208 -611 28242
rect -487 28208 -453 28242
rect -329 28208 -295 28242
rect -171 28208 -137 28242
rect -13 28208 21 28242
rect 145 28208 179 28242
rect 303 28208 337 28242
rect 461 28208 495 28242
rect 619 28208 653 28242
rect 777 28208 811 28242
rect 935 28208 969 28242
rect 1093 28208 1127 28242
rect 1251 28208 1285 28242
rect 1409 28208 1443 28242
rect 1567 28208 1601 28242
rect -1593 27796 -1559 27830
rect -1435 27796 -1401 27830
rect -1277 27796 -1243 27830
rect -1119 27796 -1085 27830
rect -961 27796 -927 27830
rect -803 27796 -769 27830
rect -645 27796 -611 27830
rect -487 27796 -453 27830
rect -329 27796 -295 27830
rect -171 27796 -137 27830
rect -13 27796 21 27830
rect 145 27796 179 27830
rect 303 27796 337 27830
rect 461 27796 495 27830
rect 619 27796 653 27830
rect 777 27796 811 27830
rect 935 27796 969 27830
rect 1093 27796 1127 27830
rect 1251 27796 1285 27830
rect 1409 27796 1443 27830
rect 1567 27796 1601 27830
rect -1593 26668 -1559 26702
rect -1435 26668 -1401 26702
rect -1277 26668 -1243 26702
rect -1119 26668 -1085 26702
rect -961 26668 -927 26702
rect -803 26668 -769 26702
rect -645 26668 -611 26702
rect -487 26668 -453 26702
rect -329 26668 -295 26702
rect -171 26668 -137 26702
rect -13 26668 21 26702
rect 145 26668 179 26702
rect 303 26668 337 26702
rect 461 26668 495 26702
rect 619 26668 653 26702
rect 777 26668 811 26702
rect 935 26668 969 26702
rect 1093 26668 1127 26702
rect 1251 26668 1285 26702
rect 1409 26668 1443 26702
rect 1567 26668 1601 26702
rect -492 26219 -458 26253
rect -334 26219 -300 26253
rect -176 26219 -142 26253
rect -18 26219 16 26253
rect 140 26219 174 26253
rect 298 26219 332 26253
rect 456 26219 490 26253
rect -492 25109 -458 25143
rect -334 25109 -300 25143
rect -176 25109 -142 25143
rect -18 25109 16 25143
rect 140 25109 174 25143
rect 298 25109 332 25143
rect 456 25109 490 25143
rect -492 24699 -458 24733
rect -334 24699 -300 24733
rect -176 24699 -142 24733
rect -18 24699 16 24733
rect 140 24699 174 24733
rect 298 24699 332 24733
rect 456 24699 490 24733
rect -492 23589 -458 23623
rect -334 23589 -300 23623
rect -176 23589 -142 23623
rect -18 23589 16 23623
rect 140 23589 174 23623
rect 298 23589 332 23623
rect 456 23589 490 23623
rect -1467 23178 -1433 23212
rect -1399 23178 -1365 23212
rect -1209 23178 -1175 23212
rect -1141 23178 -1107 23212
rect -951 23178 -917 23212
rect -883 23178 -849 23212
rect -693 23178 -659 23212
rect -625 23178 -591 23212
rect -435 23178 -401 23212
rect -367 23178 -333 23212
rect -177 23178 -143 23212
rect -109 23178 -75 23212
rect 81 23178 115 23212
rect 149 23178 183 23212
rect 339 23178 373 23212
rect 407 23178 441 23212
rect 597 23178 631 23212
rect 665 23178 699 23212
rect 855 23178 889 23212
rect 923 23178 957 23212
rect 1113 23178 1147 23212
rect 1181 23178 1215 23212
rect 1371 23178 1405 23212
rect 1439 23178 1473 23212
rect -1467 22068 -1433 22102
rect -1399 22068 -1365 22102
rect -1209 22068 -1175 22102
rect -1141 22068 -1107 22102
rect -951 22068 -917 22102
rect -883 22068 -849 22102
rect -693 22068 -659 22102
rect -625 22068 -591 22102
rect -435 22068 -401 22102
rect -367 22068 -333 22102
rect -177 22068 -143 22102
rect -109 22068 -75 22102
rect 81 22068 115 22102
rect 149 22068 183 22102
rect 339 22068 373 22102
rect 407 22068 441 22102
rect 597 22068 631 22102
rect 665 22068 699 22102
rect 855 22068 889 22102
rect 923 22068 957 22102
rect 1113 22068 1147 22102
rect 1181 22068 1215 22102
rect 1371 22068 1405 22102
rect 1439 22068 1473 22102
rect -1727 21658 -1693 21692
rect -1659 21658 -1625 21692
rect -1469 21658 -1435 21692
rect -1401 21658 -1367 21692
rect -1211 21658 -1177 21692
rect -1143 21658 -1109 21692
rect -953 21658 -919 21692
rect -885 21658 -851 21692
rect -695 21658 -661 21692
rect -627 21658 -593 21692
rect -437 21658 -403 21692
rect -369 21658 -335 21692
rect -179 21658 -145 21692
rect -111 21658 -77 21692
rect 79 21658 113 21692
rect 147 21658 181 21692
rect 337 21658 371 21692
rect 405 21658 439 21692
rect 595 21658 629 21692
rect 663 21658 697 21692
rect 853 21658 887 21692
rect 921 21658 955 21692
rect 1111 21658 1145 21692
rect 1179 21658 1213 21692
rect 1369 21658 1403 21692
rect 1437 21658 1471 21692
rect 1627 21658 1661 21692
rect 1695 21658 1729 21692
rect -1727 20548 -1693 20582
rect -1659 20548 -1625 20582
rect -1469 20548 -1435 20582
rect -1401 20548 -1367 20582
rect -1211 20548 -1177 20582
rect -1143 20548 -1109 20582
rect -953 20548 -919 20582
rect -885 20548 -851 20582
rect -695 20548 -661 20582
rect -627 20548 -593 20582
rect -437 20548 -403 20582
rect -369 20548 -335 20582
rect -179 20548 -145 20582
rect -111 20548 -77 20582
rect 79 20548 113 20582
rect 147 20548 181 20582
rect 337 20548 371 20582
rect 405 20548 439 20582
rect 595 20548 629 20582
rect 663 20548 697 20582
rect 853 20548 887 20582
rect 921 20548 955 20582
rect 1111 20548 1145 20582
rect 1179 20548 1213 20582
rect 1369 20548 1403 20582
rect 1437 20548 1471 20582
rect 1627 20548 1661 20582
rect 1695 20548 1729 20582
rect -3672 19202 -3638 19370
rect -2544 19202 -2510 19370
rect -2436 19202 -2402 19370
rect -1308 19202 -1274 19370
rect -1200 19202 -1166 19370
rect -72 19202 -38 19370
rect 36 19202 70 19370
rect 1164 19202 1198 19370
rect 1272 19202 1306 19370
rect 2400 19202 2434 19370
rect 2508 19202 2542 19370
rect 3636 19202 3670 19370
rect -3672 18612 -3638 18780
rect -2544 18612 -2510 18780
rect -2436 18612 -2402 18780
rect -1308 18612 -1274 18780
rect -1200 18612 -1166 18780
rect -72 18612 -38 18780
rect 36 18612 70 18780
rect 1164 18612 1198 18780
rect 1272 18612 1306 18780
rect 2400 18612 2434 18780
rect 2508 18612 2542 18780
rect 3636 18612 3670 18780
rect -902 17822 -868 17990
rect -542 17822 -508 17990
rect -434 17822 -400 17990
rect -74 17822 -40 17990
rect 34 17822 68 17990
rect 394 17822 428 17990
rect 502 17822 536 17990
rect 862 17822 896 17990
rect -682 17297 -648 17365
rect -72 17297 -38 17365
rect 36 17297 70 17365
rect 646 17297 680 17365
rect -3617 16672 -3583 16840
rect -2507 16672 -2473 16840
rect -2399 16672 -2365 16840
rect -1289 16672 -1255 16840
rect -1181 16672 -1147 16840
rect -71 16672 -37 16840
rect 37 16672 71 16840
rect 1147 16672 1181 16840
rect 1255 16672 1289 16840
rect 2365 16672 2399 16840
rect 2473 16672 2507 16840
rect 3583 16672 3617 16840
<< xpolycontact >>
rect -7134 30796 -6702 31942
rect -4702 30796 -4270 31942
rect -7134 29296 -6702 30442
rect -4702 29296 -4270 30442
rect 4274 30766 4706 31912
rect 6706 30766 7138 31912
rect 4274 29286 4706 30432
rect 6706 29286 7138 30432
rect -2843 15732 -1697 16164
rect -2843 1500 -1697 1932
rect -1323 15732 -177 16164
rect -1323 1500 -177 1932
rect 187 15738 1333 16170
rect 187 1506 1333 1938
rect 1697 15738 2843 16170
rect 1697 1506 2843 1938
<< xpolyres >>
rect -6702 30796 -4702 31942
rect -6702 29296 -4702 30442
rect 4706 30766 6706 31912
rect 4706 29286 6706 30432
rect -2843 1932 -1697 15732
rect -1323 1932 -177 15732
rect 187 1938 1333 15738
rect 1697 1938 2843 15738
<< locali >>
rect -7264 32038 -7168 32072
rect -4236 32038 -4140 32072
rect -7264 31976 -7230 32038
rect -4174 31976 -4140 32038
rect -7264 30700 -7230 30762
rect 4144 32008 4261 32042
rect 4295 32008 4329 32042
rect 4363 32008 4397 32042
rect 4431 32008 4465 32042
rect 4499 32008 4533 32042
rect 4567 32008 4601 32042
rect 4635 32008 4669 32042
rect 4703 32008 4737 32042
rect 4771 32008 4805 32042
rect 4839 32008 4873 32042
rect 4907 32008 4941 32042
rect 4975 32008 5009 32042
rect 5043 32008 5077 32042
rect 5111 32008 5145 32042
rect 5179 32008 5213 32042
rect 5247 32008 5281 32042
rect 5315 32008 5349 32042
rect 5383 32008 5417 32042
rect 5451 32008 5485 32042
rect 5519 32008 5553 32042
rect 5587 32008 5621 32042
rect 5655 32008 5689 32042
rect 5723 32008 5757 32042
rect 5791 32008 5825 32042
rect 5859 32008 5893 32042
rect 5927 32008 5961 32042
rect 5995 32008 6029 32042
rect 6063 32008 6097 32042
rect 6131 32008 6165 32042
rect 6199 32008 6233 32042
rect 6267 32008 6301 32042
rect 6335 32008 6369 32042
rect 6403 32008 6437 32042
rect 6471 32008 6505 32042
rect 6539 32008 6573 32042
rect 6607 32008 6641 32042
rect 6675 32008 6709 32042
rect 6743 32008 6777 32042
rect 6811 32008 6845 32042
rect 6879 32008 6913 32042
rect 6947 32008 6981 32042
rect 7015 32008 7049 32042
rect 7083 32008 7117 32042
rect 7151 32008 7268 32042
rect 4144 31934 4178 32008
rect 7234 31934 7268 32008
rect 4144 31866 4178 31900
rect 4144 31798 4178 31832
rect 4144 31730 4178 31764
rect 4144 31662 4178 31696
rect 4144 31594 4178 31628
rect 4144 31526 4178 31560
rect 4144 31458 4178 31492
rect 4144 31390 4178 31424
rect 4144 31322 4178 31356
rect 4144 31254 4178 31288
rect 4144 31186 4178 31220
rect -4174 30700 -4140 30762
rect -7264 30666 -7168 30700
rect -4236 30666 -4140 30700
rect -3286 31108 -3174 31142
rect -3140 31108 -3106 31142
rect -3072 31108 -3038 31142
rect -3004 31108 -2970 31142
rect -2936 31108 -2902 31142
rect -2868 31108 -2834 31142
rect -2800 31108 -2766 31142
rect -2732 31108 -2698 31142
rect -2664 31108 -2630 31142
rect -2596 31108 -2562 31142
rect -2528 31108 -2494 31142
rect -2460 31108 -2426 31142
rect -2392 31108 -2358 31142
rect -2324 31108 -2290 31142
rect -2256 31108 -2222 31142
rect -2188 31108 -2154 31142
rect -2120 31108 -2086 31142
rect -2052 31108 -2018 31142
rect -1984 31108 -1950 31142
rect -1916 31108 -1882 31142
rect -1848 31108 -1814 31142
rect -1780 31108 -1746 31142
rect -1712 31108 -1678 31142
rect -1644 31108 -1610 31142
rect -1562 31108 -1542 31142
rect -1490 31108 -1474 31142
rect -1418 31108 -1406 31142
rect -1346 31108 -1338 31142
rect -1274 31108 -1270 31142
rect -1168 31108 -1164 31142
rect -1100 31108 -1092 31142
rect -1032 31108 -1020 31142
rect -964 31108 -948 31142
rect -896 31108 -876 31142
rect -828 31108 -804 31142
rect -760 31108 -732 31142
rect -692 31108 -660 31142
rect -624 31108 -590 31142
rect -554 31108 -522 31142
rect -482 31108 -454 31142
rect -410 31108 -386 31142
rect -338 31108 -318 31142
rect -266 31108 -250 31142
rect -194 31108 -182 31142
rect -122 31108 -114 31142
rect -50 31108 -46 31142
rect 56 31108 60 31142
rect 124 31108 132 31142
rect 192 31108 204 31142
rect 260 31108 276 31142
rect 328 31108 348 31142
rect 396 31108 420 31142
rect 464 31108 492 31142
rect 532 31108 564 31142
rect 600 31108 634 31142
rect 670 31108 702 31142
rect 742 31108 770 31142
rect 814 31108 838 31142
rect 886 31108 906 31142
rect 958 31108 974 31142
rect 1030 31108 1042 31142
rect 1102 31108 1110 31142
rect 1174 31108 1178 31142
rect 1280 31108 1284 31142
rect 1348 31108 1356 31142
rect 1416 31108 1428 31142
rect 1484 31108 1500 31142
rect 1552 31108 1572 31142
rect 1620 31108 1654 31142
rect 1688 31108 1722 31142
rect 1756 31108 1790 31142
rect 1824 31108 1858 31142
rect 1892 31108 1926 31142
rect 1960 31108 1994 31142
rect 2028 31108 2062 31142
rect 2096 31108 2130 31142
rect 2164 31108 2198 31142
rect 2232 31108 2266 31142
rect 2300 31108 2334 31142
rect 2368 31108 2402 31142
rect 2436 31108 2470 31142
rect 2504 31108 2538 31142
rect 2572 31108 2606 31142
rect 2640 31108 2674 31142
rect 2708 31108 2742 31142
rect 2776 31108 2810 31142
rect 2844 31108 2878 31142
rect 2912 31108 2946 31142
rect 2980 31108 3014 31142
rect 3048 31108 3082 31142
rect 3116 31108 3150 31142
rect 3184 31108 3296 31142
rect -3286 31020 -3252 31108
rect -3126 31006 -3093 31040
rect -3059 31006 -3026 31040
rect -2968 31006 -2935 31040
rect -2901 31006 -2868 31040
rect -2810 31006 -2777 31040
rect -2743 31006 -2710 31040
rect -2652 31006 -2619 31040
rect -2585 31006 -2552 31040
rect -2494 31006 -2461 31040
rect -2427 31006 -2394 31040
rect -2336 31006 -2303 31040
rect -2269 31006 -2236 31040
rect -2178 31006 -2145 31040
rect -2111 31006 -2078 31040
rect -2020 31006 -1987 31040
rect -1953 31006 -1920 31040
rect -1862 31006 -1829 31040
rect -1795 31006 -1762 31040
rect -1704 31006 -1671 31040
rect -1637 31006 -1604 31040
rect -1546 31006 -1513 31040
rect -1479 31006 -1446 31040
rect -1388 31006 -1355 31040
rect -1321 31006 -1288 31040
rect -1230 31006 -1197 31040
rect -1163 31006 -1130 31040
rect -1072 31006 -1039 31040
rect -1005 31006 -972 31040
rect -914 31006 -881 31040
rect -847 31006 -814 31040
rect -756 31006 -723 31040
rect -689 31006 -656 31040
rect -598 31006 -565 31040
rect -531 31006 -498 31040
rect -440 31006 -407 31040
rect -373 31006 -340 31040
rect -282 31006 -249 31040
rect -215 31006 -182 31040
rect -124 31006 -91 31040
rect -57 31006 -24 31040
rect 34 31006 67 31040
rect 101 31006 134 31040
rect 192 31006 225 31040
rect 259 31006 292 31040
rect 350 31006 383 31040
rect 417 31006 450 31040
rect 508 31006 541 31040
rect 575 31006 608 31040
rect 666 31006 699 31040
rect 733 31006 766 31040
rect 824 31006 857 31040
rect 891 31006 924 31040
rect 982 31006 1015 31040
rect 1049 31006 1082 31040
rect 1140 31006 1173 31040
rect 1207 31006 1240 31040
rect 1298 31006 1331 31040
rect 1365 31006 1398 31040
rect 1456 31006 1489 31040
rect 1523 31006 1556 31040
rect 1614 31006 1647 31040
rect 1681 31006 1714 31040
rect 1772 31006 1805 31040
rect 1839 31006 1872 31040
rect 1930 31006 1963 31040
rect 1997 31006 2030 31040
rect 2088 31006 2121 31040
rect 2155 31006 2188 31040
rect 2246 31006 2279 31040
rect 2313 31006 2346 31040
rect 2404 31006 2437 31040
rect 2471 31006 2504 31040
rect 2562 31006 2595 31040
rect 2629 31006 2662 31040
rect 2720 31006 2753 31040
rect 2787 31006 2820 31040
rect 2878 31006 2911 31040
rect 2945 31006 2978 31040
rect 3036 31006 3069 31040
rect 3103 31006 3136 31040
rect 3262 31020 3296 31108
rect -3286 30952 -3252 30986
rect -3286 30884 -3252 30918
rect -3286 30816 -3252 30850
rect -3286 30748 -3252 30782
rect -3286 30680 -3252 30714
rect -5750 30572 -5620 30666
rect -3286 30612 -3252 30646
rect -7264 30538 -7168 30572
rect -4236 30538 -4140 30572
rect -7264 30476 -7230 30538
rect -4174 30476 -4140 30538
rect -7264 29200 -7230 29262
rect -3286 30544 -3252 30578
rect -3286 30476 -3252 30510
rect -3286 30408 -3252 30442
rect -3286 30340 -3252 30374
rect -3286 30272 -3252 30306
rect -3286 30204 -3252 30238
rect -3286 30136 -3252 30170
rect -3286 30068 -3252 30102
rect -3286 30000 -3252 30034
rect -3286 29932 -3252 29966
rect -3172 30944 -3138 30963
rect -3172 30872 -3138 30884
rect -3172 30800 -3138 30816
rect -3172 30728 -3138 30748
rect -3172 30656 -3138 30680
rect -3172 30584 -3138 30612
rect -3172 30512 -3138 30544
rect -3172 30442 -3138 30476
rect -3172 30374 -3138 30406
rect -3172 30306 -3138 30334
rect -3172 30238 -3138 30262
rect -3172 30170 -3138 30190
rect -3172 30102 -3138 30118
rect -3172 30034 -3138 30046
rect -3172 29955 -3138 29974
rect -3014 30944 -2980 30963
rect -3014 30872 -2980 30884
rect -3014 30800 -2980 30816
rect -3014 30728 -2980 30748
rect -3014 30656 -2980 30680
rect -3014 30584 -2980 30612
rect -3014 30512 -2980 30544
rect -3014 30442 -2980 30476
rect -3014 30374 -2980 30406
rect -3014 30306 -2980 30334
rect -3014 30238 -2980 30262
rect -3014 30170 -2980 30190
rect -3014 30102 -2980 30118
rect -3014 30034 -2980 30046
rect -3014 29955 -2980 29974
rect -2856 30944 -2822 30963
rect -2856 30872 -2822 30884
rect -2856 30800 -2822 30816
rect -2856 30728 -2822 30748
rect -2856 30656 -2822 30680
rect -2856 30584 -2822 30612
rect -2856 30512 -2822 30544
rect -2856 30442 -2822 30476
rect -2856 30374 -2822 30406
rect -2856 30306 -2822 30334
rect -2856 30238 -2822 30262
rect -2856 30170 -2822 30190
rect -2856 30102 -2822 30118
rect -2856 30034 -2822 30046
rect -2856 29955 -2822 29974
rect -2698 30944 -2664 30963
rect -2698 30872 -2664 30884
rect -2698 30800 -2664 30816
rect -2698 30728 -2664 30748
rect -2698 30656 -2664 30680
rect -2698 30584 -2664 30612
rect -2698 30512 -2664 30544
rect -2698 30442 -2664 30476
rect -2698 30374 -2664 30406
rect -2698 30306 -2664 30334
rect -2698 30238 -2664 30262
rect -2698 30170 -2664 30190
rect -2698 30102 -2664 30118
rect -2698 30034 -2664 30046
rect -2698 29955 -2664 29974
rect -2540 30944 -2506 30963
rect -2540 30872 -2506 30884
rect -2540 30800 -2506 30816
rect -2540 30728 -2506 30748
rect -2540 30656 -2506 30680
rect -2540 30584 -2506 30612
rect -2540 30512 -2506 30544
rect -2540 30442 -2506 30476
rect -2540 30374 -2506 30406
rect -2540 30306 -2506 30334
rect -2540 30238 -2506 30262
rect -2540 30170 -2506 30190
rect -2540 30102 -2506 30118
rect -2540 30034 -2506 30046
rect -2540 29955 -2506 29974
rect -2382 30944 -2348 30963
rect -2382 30872 -2348 30884
rect -2382 30800 -2348 30816
rect -2382 30728 -2348 30748
rect -2382 30656 -2348 30680
rect -2382 30584 -2348 30612
rect -2382 30512 -2348 30544
rect -2382 30442 -2348 30476
rect -2382 30374 -2348 30406
rect -2382 30306 -2348 30334
rect -2382 30238 -2348 30262
rect -2382 30170 -2348 30190
rect -2382 30102 -2348 30118
rect -2382 30034 -2348 30046
rect -2382 29955 -2348 29974
rect -2224 30944 -2190 30963
rect -2224 30872 -2190 30884
rect -2224 30800 -2190 30816
rect -2224 30728 -2190 30748
rect -2224 30656 -2190 30680
rect -2224 30584 -2190 30612
rect -2224 30512 -2190 30544
rect -2224 30442 -2190 30476
rect -2224 30374 -2190 30406
rect -2224 30306 -2190 30334
rect -2224 30238 -2190 30262
rect -2224 30170 -2190 30190
rect -2224 30102 -2190 30118
rect -2224 30034 -2190 30046
rect -2224 29955 -2190 29974
rect -2066 30944 -2032 30963
rect -2066 30872 -2032 30884
rect -2066 30800 -2032 30816
rect -2066 30728 -2032 30748
rect -2066 30656 -2032 30680
rect -2066 30584 -2032 30612
rect -2066 30512 -2032 30544
rect -2066 30442 -2032 30476
rect -2066 30374 -2032 30406
rect -2066 30306 -2032 30334
rect -2066 30238 -2032 30262
rect -2066 30170 -2032 30190
rect -2066 30102 -2032 30118
rect -2066 30034 -2032 30046
rect -2066 29955 -2032 29974
rect -1908 30944 -1874 30963
rect -1908 30872 -1874 30884
rect -1908 30800 -1874 30816
rect -1908 30728 -1874 30748
rect -1908 30656 -1874 30680
rect -1908 30584 -1874 30612
rect -1908 30512 -1874 30544
rect -1908 30442 -1874 30476
rect -1908 30374 -1874 30406
rect -1908 30306 -1874 30334
rect -1908 30238 -1874 30262
rect -1908 30170 -1874 30190
rect -1908 30102 -1874 30118
rect -1908 30034 -1874 30046
rect -1908 29955 -1874 29974
rect -1750 30944 -1716 30963
rect -1750 30872 -1716 30884
rect -1750 30800 -1716 30816
rect -1750 30728 -1716 30748
rect -1750 30656 -1716 30680
rect -1750 30584 -1716 30612
rect -1750 30512 -1716 30544
rect -1750 30442 -1716 30476
rect -1750 30374 -1716 30406
rect -1750 30306 -1716 30334
rect -1750 30238 -1716 30262
rect -1750 30170 -1716 30190
rect -1750 30102 -1716 30118
rect -1750 30034 -1716 30046
rect -1750 29955 -1716 29974
rect -1592 30944 -1558 30963
rect -1592 30872 -1558 30884
rect -1592 30800 -1558 30816
rect -1592 30728 -1558 30748
rect -1592 30656 -1558 30680
rect -1592 30584 -1558 30612
rect -1592 30512 -1558 30544
rect -1592 30442 -1558 30476
rect -1592 30374 -1558 30406
rect -1592 30306 -1558 30334
rect -1592 30238 -1558 30262
rect -1592 30170 -1558 30190
rect -1592 30102 -1558 30118
rect -1592 30034 -1558 30046
rect -1592 29955 -1558 29974
rect -1434 30944 -1400 30963
rect -1434 30872 -1400 30884
rect -1434 30800 -1400 30816
rect -1434 30728 -1400 30748
rect -1434 30656 -1400 30680
rect -1434 30584 -1400 30612
rect -1434 30512 -1400 30544
rect -1434 30442 -1400 30476
rect -1434 30374 -1400 30406
rect -1434 30306 -1400 30334
rect -1434 30238 -1400 30262
rect -1434 30170 -1400 30190
rect -1434 30102 -1400 30118
rect -1434 30034 -1400 30046
rect -1434 29955 -1400 29974
rect -1276 30944 -1242 30963
rect -1276 30872 -1242 30884
rect -1276 30800 -1242 30816
rect -1276 30728 -1242 30748
rect -1276 30656 -1242 30680
rect -1276 30584 -1242 30612
rect -1276 30512 -1242 30544
rect -1276 30442 -1242 30476
rect -1276 30374 -1242 30406
rect -1276 30306 -1242 30334
rect -1276 30238 -1242 30262
rect -1276 30170 -1242 30190
rect -1276 30102 -1242 30118
rect -1276 30034 -1242 30046
rect -1276 29955 -1242 29974
rect -1118 30944 -1084 30963
rect -1118 30872 -1084 30884
rect -1118 30800 -1084 30816
rect -1118 30728 -1084 30748
rect -1118 30656 -1084 30680
rect -1118 30584 -1084 30612
rect -1118 30512 -1084 30544
rect -1118 30442 -1084 30476
rect -1118 30374 -1084 30406
rect -1118 30306 -1084 30334
rect -1118 30238 -1084 30262
rect -1118 30170 -1084 30190
rect -1118 30102 -1084 30118
rect -1118 30034 -1084 30046
rect -1118 29955 -1084 29974
rect -960 30944 -926 30963
rect -960 30872 -926 30884
rect -960 30800 -926 30816
rect -960 30728 -926 30748
rect -960 30656 -926 30680
rect -960 30584 -926 30612
rect -960 30512 -926 30544
rect -960 30442 -926 30476
rect -960 30374 -926 30406
rect -960 30306 -926 30334
rect -960 30238 -926 30262
rect -960 30170 -926 30190
rect -960 30102 -926 30118
rect -960 30034 -926 30046
rect -960 29955 -926 29974
rect -802 30944 -768 30963
rect -802 30872 -768 30884
rect -802 30800 -768 30816
rect -802 30728 -768 30748
rect -802 30656 -768 30680
rect -802 30584 -768 30612
rect -802 30512 -768 30544
rect -802 30442 -768 30476
rect -802 30374 -768 30406
rect -802 30306 -768 30334
rect -802 30238 -768 30262
rect -802 30170 -768 30190
rect -802 30102 -768 30118
rect -802 30034 -768 30046
rect -802 29955 -768 29974
rect -644 30944 -610 30963
rect -644 30872 -610 30884
rect -644 30800 -610 30816
rect -644 30728 -610 30748
rect -644 30656 -610 30680
rect -644 30584 -610 30612
rect -644 30512 -610 30544
rect -644 30442 -610 30476
rect -644 30374 -610 30406
rect -644 30306 -610 30334
rect -644 30238 -610 30262
rect -644 30170 -610 30190
rect -644 30102 -610 30118
rect -644 30034 -610 30046
rect -644 29955 -610 29974
rect -486 30944 -452 30963
rect -486 30872 -452 30884
rect -486 30800 -452 30816
rect -486 30728 -452 30748
rect -486 30656 -452 30680
rect -486 30584 -452 30612
rect -486 30512 -452 30544
rect -486 30442 -452 30476
rect -486 30374 -452 30406
rect -486 30306 -452 30334
rect -486 30238 -452 30262
rect -486 30170 -452 30190
rect -486 30102 -452 30118
rect -486 30034 -452 30046
rect -486 29955 -452 29974
rect -328 30944 -294 30963
rect -328 30872 -294 30884
rect -328 30800 -294 30816
rect -328 30728 -294 30748
rect -328 30656 -294 30680
rect -328 30584 -294 30612
rect -328 30512 -294 30544
rect -328 30442 -294 30476
rect -328 30374 -294 30406
rect -328 30306 -294 30334
rect -328 30238 -294 30262
rect -328 30170 -294 30190
rect -328 30102 -294 30118
rect -328 30034 -294 30046
rect -328 29955 -294 29974
rect -170 30944 -136 30963
rect -170 30872 -136 30884
rect -170 30800 -136 30816
rect -170 30728 -136 30748
rect -170 30656 -136 30680
rect -170 30584 -136 30612
rect -170 30512 -136 30544
rect -170 30442 -136 30476
rect -170 30374 -136 30406
rect -170 30306 -136 30334
rect -170 30238 -136 30262
rect -170 30170 -136 30190
rect -170 30102 -136 30118
rect -170 30034 -136 30046
rect -170 29955 -136 29974
rect -12 30944 22 30963
rect -12 30872 22 30884
rect -12 30800 22 30816
rect -12 30728 22 30748
rect -12 30656 22 30680
rect -12 30584 22 30612
rect -12 30512 22 30544
rect -12 30442 22 30476
rect -12 30374 22 30406
rect -12 30306 22 30334
rect -12 30238 22 30262
rect -12 30170 22 30190
rect -12 30102 22 30118
rect -12 30034 22 30046
rect -12 29955 22 29974
rect 146 30944 180 30963
rect 146 30872 180 30884
rect 146 30800 180 30816
rect 146 30728 180 30748
rect 146 30656 180 30680
rect 146 30584 180 30612
rect 146 30512 180 30544
rect 146 30442 180 30476
rect 146 30374 180 30406
rect 146 30306 180 30334
rect 146 30238 180 30262
rect 146 30170 180 30190
rect 146 30102 180 30118
rect 146 30034 180 30046
rect 146 29955 180 29974
rect 304 30944 338 30963
rect 304 30872 338 30884
rect 304 30800 338 30816
rect 304 30728 338 30748
rect 304 30656 338 30680
rect 304 30584 338 30612
rect 304 30512 338 30544
rect 304 30442 338 30476
rect 304 30374 338 30406
rect 304 30306 338 30334
rect 304 30238 338 30262
rect 304 30170 338 30190
rect 304 30102 338 30118
rect 304 30034 338 30046
rect 304 29955 338 29974
rect 462 30944 496 30963
rect 462 30872 496 30884
rect 462 30800 496 30816
rect 462 30728 496 30748
rect 462 30656 496 30680
rect 462 30584 496 30612
rect 462 30512 496 30544
rect 462 30442 496 30476
rect 462 30374 496 30406
rect 462 30306 496 30334
rect 462 30238 496 30262
rect 462 30170 496 30190
rect 462 30102 496 30118
rect 462 30034 496 30046
rect 462 29955 496 29974
rect 620 30944 654 30963
rect 620 30872 654 30884
rect 620 30800 654 30816
rect 620 30728 654 30748
rect 620 30656 654 30680
rect 620 30584 654 30612
rect 620 30512 654 30544
rect 620 30442 654 30476
rect 620 30374 654 30406
rect 620 30306 654 30334
rect 620 30238 654 30262
rect 620 30170 654 30190
rect 620 30102 654 30118
rect 620 30034 654 30046
rect 620 29955 654 29974
rect 778 30944 812 30963
rect 778 30872 812 30884
rect 778 30800 812 30816
rect 778 30728 812 30748
rect 778 30656 812 30680
rect 778 30584 812 30612
rect 778 30512 812 30544
rect 778 30442 812 30476
rect 778 30374 812 30406
rect 778 30306 812 30334
rect 778 30238 812 30262
rect 778 30170 812 30190
rect 778 30102 812 30118
rect 778 30034 812 30046
rect 778 29955 812 29974
rect 936 30944 970 30963
rect 936 30872 970 30884
rect 936 30800 970 30816
rect 936 30728 970 30748
rect 936 30656 970 30680
rect 936 30584 970 30612
rect 936 30512 970 30544
rect 936 30442 970 30476
rect 936 30374 970 30406
rect 936 30306 970 30334
rect 936 30238 970 30262
rect 936 30170 970 30190
rect 936 30102 970 30118
rect 936 30034 970 30046
rect 936 29955 970 29974
rect 1094 30944 1128 30963
rect 1094 30872 1128 30884
rect 1094 30800 1128 30816
rect 1094 30728 1128 30748
rect 1094 30656 1128 30680
rect 1094 30584 1128 30612
rect 1094 30512 1128 30544
rect 1094 30442 1128 30476
rect 1094 30374 1128 30406
rect 1094 30306 1128 30334
rect 1094 30238 1128 30262
rect 1094 30170 1128 30190
rect 1094 30102 1128 30118
rect 1094 30034 1128 30046
rect 1094 29955 1128 29974
rect 1252 30944 1286 30963
rect 1252 30872 1286 30884
rect 1252 30800 1286 30816
rect 1252 30728 1286 30748
rect 1252 30656 1286 30680
rect 1252 30584 1286 30612
rect 1252 30512 1286 30544
rect 1252 30442 1286 30476
rect 1252 30374 1286 30406
rect 1252 30306 1286 30334
rect 1252 30238 1286 30262
rect 1252 30170 1286 30190
rect 1252 30102 1286 30118
rect 1252 30034 1286 30046
rect 1252 29955 1286 29974
rect 1410 30944 1444 30963
rect 1410 30872 1444 30884
rect 1410 30800 1444 30816
rect 1410 30728 1444 30748
rect 1410 30656 1444 30680
rect 1410 30584 1444 30612
rect 1410 30512 1444 30544
rect 1410 30442 1444 30476
rect 1410 30374 1444 30406
rect 1410 30306 1444 30334
rect 1410 30238 1444 30262
rect 1410 30170 1444 30190
rect 1410 30102 1444 30118
rect 1410 30034 1444 30046
rect 1410 29955 1444 29974
rect 1568 30944 1602 30963
rect 1568 30872 1602 30884
rect 1568 30800 1602 30816
rect 1568 30728 1602 30748
rect 1568 30656 1602 30680
rect 1568 30584 1602 30612
rect 1568 30512 1602 30544
rect 1568 30442 1602 30476
rect 1568 30374 1602 30406
rect 1568 30306 1602 30334
rect 1568 30238 1602 30262
rect 1568 30170 1602 30190
rect 1568 30102 1602 30118
rect 1568 30034 1602 30046
rect 1568 29955 1602 29974
rect 1726 30944 1760 30963
rect 1726 30872 1760 30884
rect 1726 30800 1760 30816
rect 1726 30728 1760 30748
rect 1726 30656 1760 30680
rect 1726 30584 1760 30612
rect 1726 30512 1760 30544
rect 1726 30442 1760 30476
rect 1726 30374 1760 30406
rect 1726 30306 1760 30334
rect 1726 30238 1760 30262
rect 1726 30170 1760 30190
rect 1726 30102 1760 30118
rect 1726 30034 1760 30046
rect 1726 29955 1760 29974
rect 1884 30944 1918 30963
rect 1884 30872 1918 30884
rect 1884 30800 1918 30816
rect 1884 30728 1918 30748
rect 1884 30656 1918 30680
rect 1884 30584 1918 30612
rect 1884 30512 1918 30544
rect 1884 30442 1918 30476
rect 1884 30374 1918 30406
rect 1884 30306 1918 30334
rect 1884 30238 1918 30262
rect 1884 30170 1918 30190
rect 1884 30102 1918 30118
rect 1884 30034 1918 30046
rect 1884 29955 1918 29974
rect 2042 30944 2076 30963
rect 2042 30872 2076 30884
rect 2042 30800 2076 30816
rect 2042 30728 2076 30748
rect 2042 30656 2076 30680
rect 2042 30584 2076 30612
rect 2042 30512 2076 30544
rect 2042 30442 2076 30476
rect 2042 30374 2076 30406
rect 2042 30306 2076 30334
rect 2042 30238 2076 30262
rect 2042 30170 2076 30190
rect 2042 30102 2076 30118
rect 2042 30034 2076 30046
rect 2042 29955 2076 29974
rect 2200 30944 2234 30963
rect 2200 30872 2234 30884
rect 2200 30800 2234 30816
rect 2200 30728 2234 30748
rect 2200 30656 2234 30680
rect 2200 30584 2234 30612
rect 2200 30512 2234 30544
rect 2200 30442 2234 30476
rect 2200 30374 2234 30406
rect 2200 30306 2234 30334
rect 2200 30238 2234 30262
rect 2200 30170 2234 30190
rect 2200 30102 2234 30118
rect 2200 30034 2234 30046
rect 2200 29955 2234 29974
rect 2358 30944 2392 30963
rect 2358 30872 2392 30884
rect 2358 30800 2392 30816
rect 2358 30728 2392 30748
rect 2358 30656 2392 30680
rect 2358 30584 2392 30612
rect 2358 30512 2392 30544
rect 2358 30442 2392 30476
rect 2358 30374 2392 30406
rect 2358 30306 2392 30334
rect 2358 30238 2392 30262
rect 2358 30170 2392 30190
rect 2358 30102 2392 30118
rect 2358 30034 2392 30046
rect 2358 29955 2392 29974
rect 2516 30944 2550 30963
rect 2516 30872 2550 30884
rect 2516 30800 2550 30816
rect 2516 30728 2550 30748
rect 2516 30656 2550 30680
rect 2516 30584 2550 30612
rect 2516 30512 2550 30544
rect 2516 30442 2550 30476
rect 2516 30374 2550 30406
rect 2516 30306 2550 30334
rect 2516 30238 2550 30262
rect 2516 30170 2550 30190
rect 2516 30102 2550 30118
rect 2516 30034 2550 30046
rect 2516 29955 2550 29974
rect 2674 30944 2708 30963
rect 2674 30872 2708 30884
rect 2674 30800 2708 30816
rect 2674 30728 2708 30748
rect 2674 30656 2708 30680
rect 2674 30584 2708 30612
rect 2674 30512 2708 30544
rect 2674 30442 2708 30476
rect 2674 30374 2708 30406
rect 2674 30306 2708 30334
rect 2674 30238 2708 30262
rect 2674 30170 2708 30190
rect 2674 30102 2708 30118
rect 2674 30034 2708 30046
rect 2674 29955 2708 29974
rect 2832 30944 2866 30963
rect 2832 30872 2866 30884
rect 2832 30800 2866 30816
rect 2832 30728 2866 30748
rect 2832 30656 2866 30680
rect 2832 30584 2866 30612
rect 2832 30512 2866 30544
rect 2832 30442 2866 30476
rect 2832 30374 2866 30406
rect 2832 30306 2866 30334
rect 2832 30238 2866 30262
rect 2832 30170 2866 30190
rect 2832 30102 2866 30118
rect 2832 30034 2866 30046
rect 2832 29955 2866 29974
rect 2990 30944 3024 30963
rect 2990 30872 3024 30884
rect 2990 30800 3024 30816
rect 2990 30728 3024 30748
rect 2990 30656 3024 30680
rect 2990 30584 3024 30612
rect 2990 30512 3024 30544
rect 2990 30442 3024 30476
rect 2990 30374 3024 30406
rect 2990 30306 3024 30334
rect 2990 30238 3024 30262
rect 2990 30170 3024 30190
rect 2990 30102 3024 30118
rect 2990 30034 3024 30046
rect 2990 29955 3024 29974
rect 3148 30944 3182 30963
rect 3148 30872 3182 30884
rect 3148 30800 3182 30816
rect 3148 30728 3182 30748
rect 3148 30656 3182 30680
rect 3148 30584 3182 30612
rect 3148 30512 3182 30544
rect 3148 30442 3182 30476
rect 3148 30374 3182 30406
rect 3148 30306 3182 30334
rect 3148 30238 3182 30262
rect 3148 30170 3182 30190
rect 3148 30102 3182 30118
rect 3148 30034 3182 30046
rect 3148 29955 3182 29974
rect 3262 30952 3296 30986
rect 3262 30884 3296 30918
rect 3262 30816 3296 30850
rect 3262 30748 3296 30782
rect 3262 30680 3296 30714
rect 3262 30612 3296 30646
rect 4144 31118 4178 31152
rect 4144 31050 4178 31084
rect 4144 30982 4178 31016
rect 4144 30914 4178 30948
rect 4144 30846 4178 30880
rect 4144 30778 4178 30812
rect 7234 31866 7268 31900
rect 7234 31798 7268 31832
rect 7234 31730 7268 31764
rect 7234 31662 7268 31696
rect 7234 31594 7268 31628
rect 7234 31526 7268 31560
rect 7234 31458 7268 31492
rect 7234 31390 7268 31424
rect 7234 31322 7268 31356
rect 7234 31254 7268 31288
rect 7234 31186 7268 31220
rect 7234 31118 7268 31152
rect 7234 31050 7268 31084
rect 7234 30982 7268 31016
rect 7234 30914 7268 30948
rect 7234 30846 7268 30880
rect 7234 30778 7268 30812
rect 4144 30670 4178 30744
rect 7234 30670 7268 30744
rect 4144 30636 4261 30670
rect 4295 30636 4329 30670
rect 4363 30636 4397 30670
rect 4431 30636 4465 30670
rect 4499 30636 4533 30670
rect 4567 30636 4601 30670
rect 4635 30636 4669 30670
rect 4703 30636 4737 30670
rect 4771 30636 4805 30670
rect 4839 30636 4873 30670
rect 4907 30636 4941 30670
rect 4975 30636 5009 30670
rect 5043 30636 5077 30670
rect 5111 30636 5145 30670
rect 5179 30636 5213 30670
rect 5247 30636 5281 30670
rect 5315 30636 5349 30670
rect 5383 30636 5417 30670
rect 5451 30636 5485 30670
rect 5519 30636 5553 30670
rect 5587 30636 5621 30670
rect 5655 30636 5689 30670
rect 5723 30636 5757 30670
rect 5791 30636 5825 30670
rect 5859 30636 5893 30670
rect 5927 30636 5961 30670
rect 5995 30636 6029 30670
rect 6063 30636 6097 30670
rect 6131 30636 6165 30670
rect 6199 30636 6233 30670
rect 6267 30636 6301 30670
rect 6335 30636 6369 30670
rect 6403 30636 6437 30670
rect 6471 30636 6505 30670
rect 6539 30636 6573 30670
rect 6607 30636 6641 30670
rect 6675 30636 6709 30670
rect 6743 30636 6777 30670
rect 6811 30636 6845 30670
rect 6879 30636 6913 30670
rect 6947 30636 6981 30670
rect 7015 30636 7049 30670
rect 7083 30636 7117 30670
rect 7151 30636 7268 30670
rect 3262 30544 3296 30578
rect 5608 30562 5878 30636
rect 3262 30476 3296 30510
rect 3262 30408 3296 30442
rect 3262 30340 3296 30374
rect 3262 30272 3296 30306
rect 3262 30204 3296 30238
rect 3262 30136 3296 30170
rect 3262 30068 3296 30102
rect 3262 30000 3296 30034
rect 3262 29932 3296 29966
rect -3286 29810 -3252 29898
rect -3126 29878 -3093 29912
rect -3059 29878 -3026 29912
rect -2968 29878 -2935 29912
rect -2901 29878 -2868 29912
rect -2810 29878 -2777 29912
rect -2743 29878 -2710 29912
rect -2652 29878 -2619 29912
rect -2585 29878 -2552 29912
rect -2494 29878 -2461 29912
rect -2427 29878 -2394 29912
rect -2336 29878 -2303 29912
rect -2269 29878 -2236 29912
rect -2178 29878 -2145 29912
rect -2111 29878 -2078 29912
rect -2020 29878 -1987 29912
rect -1953 29878 -1920 29912
rect -1862 29878 -1829 29912
rect -1795 29878 -1762 29912
rect -1704 29878 -1671 29912
rect -1637 29878 -1604 29912
rect -1546 29878 -1513 29912
rect -1479 29878 -1446 29912
rect -1388 29878 -1355 29912
rect -1321 29878 -1288 29912
rect -1230 29878 -1197 29912
rect -1163 29878 -1130 29912
rect -1072 29878 -1039 29912
rect -1005 29878 -972 29912
rect -914 29878 -881 29912
rect -847 29878 -814 29912
rect -756 29878 -723 29912
rect -689 29878 -656 29912
rect -598 29878 -565 29912
rect -531 29878 -498 29912
rect -440 29878 -407 29912
rect -373 29878 -340 29912
rect -282 29878 -249 29912
rect -215 29878 -182 29912
rect -124 29878 -91 29912
rect -57 29878 -24 29912
rect 34 29878 67 29912
rect 101 29878 134 29912
rect 192 29878 225 29912
rect 259 29878 292 29912
rect 350 29878 383 29912
rect 417 29878 450 29912
rect 508 29878 541 29912
rect 575 29878 608 29912
rect 666 29878 699 29912
rect 733 29878 766 29912
rect 824 29878 857 29912
rect 891 29878 924 29912
rect 982 29878 1015 29912
rect 1049 29878 1082 29912
rect 1140 29878 1173 29912
rect 1207 29878 1240 29912
rect 1298 29878 1331 29912
rect 1365 29878 1398 29912
rect 1456 29878 1489 29912
rect 1523 29878 1556 29912
rect 1614 29878 1647 29912
rect 1681 29878 1714 29912
rect 1772 29878 1805 29912
rect 1839 29878 1872 29912
rect 1930 29878 1963 29912
rect 1997 29878 2030 29912
rect 2088 29878 2121 29912
rect 2155 29878 2188 29912
rect 2246 29878 2279 29912
rect 2313 29878 2346 29912
rect 2404 29878 2437 29912
rect 2471 29878 2504 29912
rect 2562 29878 2595 29912
rect 2629 29878 2662 29912
rect 2720 29878 2753 29912
rect 2787 29878 2820 29912
rect 2878 29878 2911 29912
rect 2945 29878 2978 29912
rect 3036 29878 3069 29912
rect 3103 29878 3136 29912
rect 3262 29810 3296 29898
rect -3286 29776 -3174 29810
rect -3140 29776 -3106 29810
rect -3072 29776 -3038 29810
rect -3004 29776 -2970 29810
rect -2936 29776 -2902 29810
rect -2868 29776 -2834 29810
rect -2800 29776 -2766 29810
rect -2732 29776 -2698 29810
rect -2664 29776 -2630 29810
rect -2596 29776 -2562 29810
rect -2528 29776 -2494 29810
rect -2460 29776 -2426 29810
rect -2392 29776 -2358 29810
rect -2324 29776 -2290 29810
rect -2256 29776 -2222 29810
rect -2188 29776 -2154 29810
rect -2120 29776 -2086 29810
rect -2052 29776 -2018 29810
rect -1984 29776 -1950 29810
rect -1916 29776 -1882 29810
rect -1848 29776 -1814 29810
rect -1780 29776 -1746 29810
rect -1712 29776 -1678 29810
rect -1644 29776 -1610 29810
rect -1562 29776 -1542 29810
rect -1490 29776 -1474 29810
rect -1418 29776 -1406 29810
rect -1346 29776 -1338 29810
rect -1274 29776 -1270 29810
rect -1168 29776 -1164 29810
rect -1100 29776 -1092 29810
rect -1032 29776 -1020 29810
rect -964 29776 -948 29810
rect -896 29776 -876 29810
rect -828 29776 -804 29810
rect -760 29776 -732 29810
rect -692 29776 -660 29810
rect -624 29776 -590 29810
rect -554 29776 -522 29810
rect -482 29776 -454 29810
rect -410 29776 -386 29810
rect -338 29776 -318 29810
rect -266 29776 -250 29810
rect -194 29776 -182 29810
rect -122 29776 -114 29810
rect -50 29776 -46 29810
rect 56 29776 60 29810
rect 124 29776 132 29810
rect 192 29776 204 29810
rect 260 29776 276 29810
rect 328 29776 348 29810
rect 396 29776 420 29810
rect 464 29776 492 29810
rect 532 29776 564 29810
rect 600 29776 634 29810
rect 670 29776 702 29810
rect 742 29776 770 29810
rect 814 29776 838 29810
rect 886 29776 906 29810
rect 958 29776 974 29810
rect 1030 29776 1042 29810
rect 1102 29776 1110 29810
rect 1174 29776 1178 29810
rect 1280 29776 1284 29810
rect 1348 29776 1356 29810
rect 1416 29776 1428 29810
rect 1484 29776 1500 29810
rect 1552 29776 1572 29810
rect 1620 29776 1654 29810
rect 1688 29776 1722 29810
rect 1756 29776 1790 29810
rect 1824 29776 1858 29810
rect 1892 29776 1926 29810
rect 1960 29776 1994 29810
rect 2028 29776 2062 29810
rect 2096 29776 2130 29810
rect 2164 29776 2198 29810
rect 2232 29776 2266 29810
rect 2300 29776 2334 29810
rect 2368 29776 2402 29810
rect 2436 29776 2470 29810
rect 2504 29776 2538 29810
rect 2572 29776 2606 29810
rect 2640 29776 2674 29810
rect 2708 29776 2742 29810
rect 2776 29776 2810 29810
rect 2844 29776 2878 29810
rect 2912 29776 2946 29810
rect 2980 29776 3014 29810
rect 3048 29776 3082 29810
rect 3116 29776 3150 29810
rect 3184 29776 3296 29810
rect 4144 30528 4261 30562
rect 4295 30528 4329 30562
rect 4363 30528 4397 30562
rect 4431 30528 4465 30562
rect 4499 30528 4533 30562
rect 4567 30528 4601 30562
rect 4635 30528 4669 30562
rect 4703 30528 4737 30562
rect 4771 30528 4805 30562
rect 4839 30528 4873 30562
rect 4907 30528 4941 30562
rect 4975 30528 5009 30562
rect 5043 30528 5077 30562
rect 5111 30528 5145 30562
rect 5179 30528 5213 30562
rect 5247 30528 5281 30562
rect 5315 30528 5349 30562
rect 5383 30528 5417 30562
rect 5451 30528 5485 30562
rect 5519 30528 5553 30562
rect 5587 30528 5621 30562
rect 5655 30528 5689 30562
rect 5723 30528 5757 30562
rect 5791 30528 5825 30562
rect 5859 30528 5893 30562
rect 5927 30528 5961 30562
rect 5995 30528 6029 30562
rect 6063 30528 6097 30562
rect 6131 30528 6165 30562
rect 6199 30528 6233 30562
rect 6267 30528 6301 30562
rect 6335 30528 6369 30562
rect 6403 30528 6437 30562
rect 6471 30528 6505 30562
rect 6539 30528 6573 30562
rect 6607 30528 6641 30562
rect 6675 30528 6709 30562
rect 6743 30528 6777 30562
rect 6811 30528 6845 30562
rect 6879 30528 6913 30562
rect 6947 30528 6981 30562
rect 7015 30528 7049 30562
rect 7083 30528 7117 30562
rect 7151 30528 7268 30562
rect 4144 30454 4178 30528
rect 7234 30454 7268 30528
rect 4144 30386 4178 30420
rect 4144 30318 4178 30352
rect 4144 30250 4178 30284
rect 4144 30182 4178 30216
rect 4144 30114 4178 30148
rect 4144 30046 4178 30080
rect 4144 29978 4178 30012
rect 4144 29910 4178 29944
rect 4144 29842 4178 29876
rect 4144 29774 4178 29808
rect 4144 29706 4178 29740
rect 4144 29638 4178 29672
rect 4144 29570 4178 29604
rect 4144 29502 4178 29536
rect -4174 29200 -4140 29262
rect -7264 29166 -7168 29200
rect -4236 29166 -4140 29200
rect -1786 29438 -1679 29472
rect -1645 29438 -1611 29472
rect -1577 29438 -1543 29472
rect -1509 29438 -1475 29472
rect -1441 29438 -1407 29472
rect -1373 29438 -1339 29472
rect -1305 29438 -1271 29472
rect -1237 29438 -1203 29472
rect -1169 29438 -1135 29472
rect -1101 29438 -1067 29472
rect -1033 29438 -999 29472
rect -965 29438 -931 29472
rect -897 29438 -863 29472
rect -807 29438 -795 29472
rect -735 29438 -727 29472
rect -663 29438 -659 29472
rect -557 29438 -553 29472
rect -489 29438 -481 29472
rect -421 29438 -409 29472
rect -353 29438 -337 29472
rect -285 29438 -265 29472
rect -217 29438 -193 29472
rect -149 29438 -121 29472
rect -81 29438 -49 29472
rect -13 29438 21 29472
rect 57 29438 89 29472
rect 129 29438 157 29472
rect 201 29438 225 29472
rect 273 29438 293 29472
rect 345 29438 361 29472
rect 417 29438 429 29472
rect 489 29438 497 29472
rect 561 29438 565 29472
rect 667 29438 671 29472
rect 735 29438 743 29472
rect 803 29438 815 29472
rect 871 29438 905 29472
rect 939 29438 973 29472
rect 1007 29438 1041 29472
rect 1075 29438 1109 29472
rect 1143 29438 1177 29472
rect 1211 29438 1245 29472
rect 1279 29438 1313 29472
rect 1347 29438 1381 29472
rect 1415 29438 1449 29472
rect 1483 29438 1517 29472
rect 1551 29438 1585 29472
rect 1619 29438 1653 29472
rect 1687 29438 1794 29472
rect -1786 29350 -1752 29438
rect -1626 29336 -1593 29370
rect -1559 29336 -1526 29370
rect -1468 29336 -1435 29370
rect -1401 29336 -1368 29370
rect -1310 29336 -1277 29370
rect -1243 29336 -1210 29370
rect -1152 29336 -1119 29370
rect -1085 29336 -1052 29370
rect -994 29336 -961 29370
rect -927 29336 -894 29370
rect -836 29336 -803 29370
rect -769 29336 -736 29370
rect -678 29336 -645 29370
rect -611 29336 -578 29370
rect -520 29336 -487 29370
rect -453 29336 -420 29370
rect -362 29336 -329 29370
rect -295 29336 -262 29370
rect -204 29336 -171 29370
rect -137 29336 -104 29370
rect -46 29336 -13 29370
rect 21 29336 54 29370
rect 112 29336 145 29370
rect 179 29336 212 29370
rect 270 29336 303 29370
rect 337 29336 370 29370
rect 428 29336 461 29370
rect 495 29336 528 29370
rect 586 29336 619 29370
rect 653 29336 686 29370
rect 744 29336 777 29370
rect 811 29336 844 29370
rect 902 29336 935 29370
rect 969 29336 1002 29370
rect 1060 29336 1093 29370
rect 1127 29336 1160 29370
rect 1218 29336 1251 29370
rect 1285 29336 1318 29370
rect 1376 29336 1409 29370
rect 1443 29336 1476 29370
rect 1534 29336 1567 29370
rect 1601 29336 1634 29370
rect 1760 29350 1794 29438
rect -1786 29282 -1752 29316
rect -1786 29214 -1752 29248
rect -1786 29146 -1752 29180
rect -1786 29078 -1752 29112
rect -1786 29010 -1752 29044
rect -1786 28942 -1752 28976
rect -1786 28874 -1752 28908
rect -1786 28806 -1752 28840
rect -1786 28738 -1752 28772
rect -1786 28670 -1752 28704
rect -1786 28602 -1752 28636
rect -1786 28534 -1752 28568
rect -1786 28466 -1752 28500
rect -1786 28398 -1752 28432
rect -1786 28330 -1752 28364
rect -1786 28262 -1752 28296
rect -1672 29274 -1638 29293
rect -1672 29202 -1638 29214
rect -1672 29130 -1638 29146
rect -1672 29058 -1638 29078
rect -1672 28986 -1638 29010
rect -1672 28914 -1638 28942
rect -1672 28842 -1638 28874
rect -1672 28772 -1638 28806
rect -1672 28704 -1638 28736
rect -1672 28636 -1638 28664
rect -1672 28568 -1638 28592
rect -1672 28500 -1638 28520
rect -1672 28432 -1638 28448
rect -1672 28364 -1638 28376
rect -1672 28285 -1638 28304
rect -1514 29274 -1480 29293
rect -1514 29202 -1480 29214
rect -1514 29130 -1480 29146
rect -1514 29058 -1480 29078
rect -1514 28986 -1480 29010
rect -1514 28914 -1480 28942
rect -1514 28842 -1480 28874
rect -1514 28772 -1480 28806
rect -1514 28704 -1480 28736
rect -1514 28636 -1480 28664
rect -1514 28568 -1480 28592
rect -1514 28500 -1480 28520
rect -1514 28432 -1480 28448
rect -1514 28364 -1480 28376
rect -1514 28285 -1480 28304
rect -1356 29274 -1322 29293
rect -1356 29202 -1322 29214
rect -1356 29130 -1322 29146
rect -1356 29058 -1322 29078
rect -1356 28986 -1322 29010
rect -1356 28914 -1322 28942
rect -1356 28842 -1322 28874
rect -1356 28772 -1322 28806
rect -1356 28704 -1322 28736
rect -1356 28636 -1322 28664
rect -1356 28568 -1322 28592
rect -1356 28500 -1322 28520
rect -1356 28432 -1322 28448
rect -1356 28364 -1322 28376
rect -1356 28285 -1322 28304
rect -1198 29274 -1164 29293
rect -1198 29202 -1164 29214
rect -1198 29130 -1164 29146
rect -1198 29058 -1164 29078
rect -1198 28986 -1164 29010
rect -1198 28914 -1164 28942
rect -1198 28842 -1164 28874
rect -1198 28772 -1164 28806
rect -1198 28704 -1164 28736
rect -1198 28636 -1164 28664
rect -1198 28568 -1164 28592
rect -1198 28500 -1164 28520
rect -1198 28432 -1164 28448
rect -1198 28364 -1164 28376
rect -1198 28285 -1164 28304
rect -1040 29274 -1006 29293
rect -1040 29202 -1006 29214
rect -1040 29130 -1006 29146
rect -1040 29058 -1006 29078
rect -1040 28986 -1006 29010
rect -1040 28914 -1006 28942
rect -1040 28842 -1006 28874
rect -1040 28772 -1006 28806
rect -1040 28704 -1006 28736
rect -1040 28636 -1006 28664
rect -1040 28568 -1006 28592
rect -1040 28500 -1006 28520
rect -1040 28432 -1006 28448
rect -1040 28364 -1006 28376
rect -1040 28285 -1006 28304
rect -882 29274 -848 29293
rect -882 29202 -848 29214
rect -882 29130 -848 29146
rect -882 29058 -848 29078
rect -882 28986 -848 29010
rect -882 28914 -848 28942
rect -882 28842 -848 28874
rect -882 28772 -848 28806
rect -882 28704 -848 28736
rect -882 28636 -848 28664
rect -882 28568 -848 28592
rect -882 28500 -848 28520
rect -882 28432 -848 28448
rect -882 28364 -848 28376
rect -882 28285 -848 28304
rect -724 29274 -690 29293
rect -724 29202 -690 29214
rect -724 29130 -690 29146
rect -724 29058 -690 29078
rect -724 28986 -690 29010
rect -724 28914 -690 28942
rect -724 28842 -690 28874
rect -724 28772 -690 28806
rect -724 28704 -690 28736
rect -724 28636 -690 28664
rect -724 28568 -690 28592
rect -724 28500 -690 28520
rect -724 28432 -690 28448
rect -724 28364 -690 28376
rect -724 28285 -690 28304
rect -566 29274 -532 29293
rect -566 29202 -532 29214
rect -566 29130 -532 29146
rect -566 29058 -532 29078
rect -566 28986 -532 29010
rect -566 28914 -532 28942
rect -566 28842 -532 28874
rect -566 28772 -532 28806
rect -566 28704 -532 28736
rect -566 28636 -532 28664
rect -566 28568 -532 28592
rect -566 28500 -532 28520
rect -566 28432 -532 28448
rect -566 28364 -532 28376
rect -566 28285 -532 28304
rect -408 29274 -374 29293
rect -408 29202 -374 29214
rect -408 29130 -374 29146
rect -408 29058 -374 29078
rect -408 28986 -374 29010
rect -408 28914 -374 28942
rect -408 28842 -374 28874
rect -408 28772 -374 28806
rect -408 28704 -374 28736
rect -408 28636 -374 28664
rect -408 28568 -374 28592
rect -408 28500 -374 28520
rect -408 28432 -374 28448
rect -408 28364 -374 28376
rect -408 28285 -374 28304
rect -250 29274 -216 29293
rect -250 29202 -216 29214
rect -250 29130 -216 29146
rect -250 29058 -216 29078
rect -250 28986 -216 29010
rect -250 28914 -216 28942
rect -250 28842 -216 28874
rect -250 28772 -216 28806
rect -250 28704 -216 28736
rect -250 28636 -216 28664
rect -250 28568 -216 28592
rect -250 28500 -216 28520
rect -250 28432 -216 28448
rect -250 28364 -216 28376
rect -250 28285 -216 28304
rect -92 29274 -58 29293
rect -92 29202 -58 29214
rect -92 29130 -58 29146
rect -92 29058 -58 29078
rect -92 28986 -58 29010
rect -92 28914 -58 28942
rect -92 28842 -58 28874
rect -92 28772 -58 28806
rect -92 28704 -58 28736
rect -92 28636 -58 28664
rect -92 28568 -58 28592
rect -92 28500 -58 28520
rect -92 28432 -58 28448
rect -92 28364 -58 28376
rect -92 28285 -58 28304
rect 66 29274 100 29293
rect 66 29202 100 29214
rect 66 29130 100 29146
rect 66 29058 100 29078
rect 66 28986 100 29010
rect 66 28914 100 28942
rect 66 28842 100 28874
rect 66 28772 100 28806
rect 66 28704 100 28736
rect 66 28636 100 28664
rect 66 28568 100 28592
rect 66 28500 100 28520
rect 66 28432 100 28448
rect 66 28364 100 28376
rect 66 28285 100 28304
rect 224 29274 258 29293
rect 224 29202 258 29214
rect 224 29130 258 29146
rect 224 29058 258 29078
rect 224 28986 258 29010
rect 224 28914 258 28942
rect 224 28842 258 28874
rect 224 28772 258 28806
rect 224 28704 258 28736
rect 224 28636 258 28664
rect 224 28568 258 28592
rect 224 28500 258 28520
rect 224 28432 258 28448
rect 224 28364 258 28376
rect 224 28285 258 28304
rect 382 29274 416 29293
rect 382 29202 416 29214
rect 382 29130 416 29146
rect 382 29058 416 29078
rect 382 28986 416 29010
rect 382 28914 416 28942
rect 382 28842 416 28874
rect 382 28772 416 28806
rect 382 28704 416 28736
rect 382 28636 416 28664
rect 382 28568 416 28592
rect 382 28500 416 28520
rect 382 28432 416 28448
rect 382 28364 416 28376
rect 382 28285 416 28304
rect 540 29274 574 29293
rect 540 29202 574 29214
rect 540 29130 574 29146
rect 540 29058 574 29078
rect 540 28986 574 29010
rect 540 28914 574 28942
rect 540 28842 574 28874
rect 540 28772 574 28806
rect 540 28704 574 28736
rect 540 28636 574 28664
rect 540 28568 574 28592
rect 540 28500 574 28520
rect 540 28432 574 28448
rect 540 28364 574 28376
rect 540 28285 574 28304
rect 698 29274 732 29293
rect 698 29202 732 29214
rect 698 29130 732 29146
rect 698 29058 732 29078
rect 698 28986 732 29010
rect 698 28914 732 28942
rect 698 28842 732 28874
rect 698 28772 732 28806
rect 698 28704 732 28736
rect 698 28636 732 28664
rect 698 28568 732 28592
rect 698 28500 732 28520
rect 698 28432 732 28448
rect 698 28364 732 28376
rect 698 28285 732 28304
rect 856 29274 890 29293
rect 856 29202 890 29214
rect 856 29130 890 29146
rect 856 29058 890 29078
rect 856 28986 890 29010
rect 856 28914 890 28942
rect 856 28842 890 28874
rect 856 28772 890 28806
rect 856 28704 890 28736
rect 856 28636 890 28664
rect 856 28568 890 28592
rect 856 28500 890 28520
rect 856 28432 890 28448
rect 856 28364 890 28376
rect 856 28285 890 28304
rect 1014 29274 1048 29293
rect 1014 29202 1048 29214
rect 1014 29130 1048 29146
rect 1014 29058 1048 29078
rect 1014 28986 1048 29010
rect 1014 28914 1048 28942
rect 1014 28842 1048 28874
rect 1014 28772 1048 28806
rect 1014 28704 1048 28736
rect 1014 28636 1048 28664
rect 1014 28568 1048 28592
rect 1014 28500 1048 28520
rect 1014 28432 1048 28448
rect 1014 28364 1048 28376
rect 1014 28285 1048 28304
rect 1172 29274 1206 29293
rect 1172 29202 1206 29214
rect 1172 29130 1206 29146
rect 1172 29058 1206 29078
rect 1172 28986 1206 29010
rect 1172 28914 1206 28942
rect 1172 28842 1206 28874
rect 1172 28772 1206 28806
rect 1172 28704 1206 28736
rect 1172 28636 1206 28664
rect 1172 28568 1206 28592
rect 1172 28500 1206 28520
rect 1172 28432 1206 28448
rect 1172 28364 1206 28376
rect 1172 28285 1206 28304
rect 1330 29274 1364 29293
rect 1330 29202 1364 29214
rect 1330 29130 1364 29146
rect 1330 29058 1364 29078
rect 1330 28986 1364 29010
rect 1330 28914 1364 28942
rect 1330 28842 1364 28874
rect 1330 28772 1364 28806
rect 1330 28704 1364 28736
rect 1330 28636 1364 28664
rect 1330 28568 1364 28592
rect 1330 28500 1364 28520
rect 1330 28432 1364 28448
rect 1330 28364 1364 28376
rect 1330 28285 1364 28304
rect 1488 29274 1522 29293
rect 1488 29202 1522 29214
rect 1488 29130 1522 29146
rect 1488 29058 1522 29078
rect 1488 28986 1522 29010
rect 1488 28914 1522 28942
rect 1488 28842 1522 28874
rect 1488 28772 1522 28806
rect 1488 28704 1522 28736
rect 1488 28636 1522 28664
rect 1488 28568 1522 28592
rect 1488 28500 1522 28520
rect 1488 28432 1522 28448
rect 1488 28364 1522 28376
rect 1488 28285 1522 28304
rect 1646 29274 1680 29293
rect 1646 29202 1680 29214
rect 1646 29130 1680 29146
rect 1646 29058 1680 29078
rect 1646 28986 1680 29010
rect 1646 28914 1680 28942
rect 1646 28842 1680 28874
rect 1646 28772 1680 28806
rect 1646 28704 1680 28736
rect 1646 28636 1680 28664
rect 1646 28568 1680 28592
rect 1646 28500 1680 28520
rect 1646 28432 1680 28448
rect 1646 28364 1680 28376
rect 1646 28285 1680 28304
rect 1760 29282 1794 29316
rect 1760 29214 1794 29248
rect 1760 29146 1794 29180
rect 4144 29434 4178 29468
rect 4144 29366 4178 29400
rect 4144 29298 4178 29332
rect 7234 30386 7268 30420
rect 7234 30318 7268 30352
rect 7234 30250 7268 30284
rect 7234 30182 7268 30216
rect 7234 30114 7268 30148
rect 7234 30046 7268 30080
rect 7234 29978 7268 30012
rect 7234 29910 7268 29944
rect 7234 29842 7268 29876
rect 7234 29774 7268 29808
rect 7234 29706 7268 29740
rect 7234 29638 7268 29672
rect 7234 29570 7268 29604
rect 7234 29502 7268 29536
rect 7234 29434 7268 29468
rect 7234 29366 7268 29400
rect 7234 29298 7268 29332
rect 4144 29190 4178 29264
rect 7234 29190 7268 29264
rect 4144 29156 4261 29190
rect 4295 29156 4329 29190
rect 4363 29156 4397 29190
rect 4431 29156 4465 29190
rect 4499 29156 4533 29190
rect 4567 29156 4601 29190
rect 4635 29156 4669 29190
rect 4703 29156 4737 29190
rect 4771 29156 4805 29190
rect 4839 29156 4873 29190
rect 4907 29156 4941 29190
rect 4975 29156 5009 29190
rect 5043 29156 5077 29190
rect 5111 29156 5145 29190
rect 5179 29156 5213 29190
rect 5247 29156 5281 29190
rect 5315 29156 5349 29190
rect 5383 29156 5417 29190
rect 5451 29180 5485 29190
rect 5519 29180 5553 29190
rect 5587 29180 5621 29190
rect 5655 29156 5689 29190
rect 5723 29156 5757 29190
rect 5791 29156 5825 29190
rect 5859 29156 5893 29190
rect 5927 29156 5961 29190
rect 5995 29156 6029 29190
rect 6063 29156 6097 29190
rect 6131 29180 6165 29190
rect 6199 29180 6233 29190
rect 6267 29180 6301 29190
rect 6298 29156 6301 29180
rect 6335 29156 6369 29190
rect 6403 29156 6437 29190
rect 6471 29156 6505 29190
rect 6539 29156 6573 29190
rect 6607 29156 6641 29190
rect 6675 29156 6709 29190
rect 6743 29156 6777 29190
rect 6811 29156 6845 29190
rect 6879 29156 6913 29190
rect 6947 29156 6981 29190
rect 7015 29156 7049 29190
rect 7083 29156 7117 29190
rect 7151 29156 7268 29190
rect 1760 29078 1794 29112
rect 1760 29010 1794 29044
rect 1760 28942 1794 28976
rect 1760 28874 1794 28908
rect 1760 28806 1794 28840
rect 1760 28738 1794 28772
rect 1760 28670 1794 28704
rect 1760 28602 1794 28636
rect 1760 28534 1794 28568
rect 1760 28466 1794 28500
rect 1760 28398 1794 28432
rect 1760 28330 1794 28364
rect 1760 28262 1794 28296
rect -1786 28140 -1752 28228
rect -1626 28208 -1593 28242
rect -1559 28208 -1526 28242
rect -1468 28208 -1435 28242
rect -1401 28208 -1368 28242
rect -1310 28208 -1277 28242
rect -1243 28208 -1210 28242
rect -1152 28208 -1119 28242
rect -1085 28208 -1052 28242
rect -994 28208 -961 28242
rect -927 28208 -894 28242
rect -836 28208 -803 28242
rect -769 28208 -736 28242
rect -678 28208 -645 28242
rect -611 28208 -578 28242
rect -520 28208 -487 28242
rect -453 28208 -420 28242
rect -362 28208 -329 28242
rect -295 28208 -262 28242
rect -204 28208 -171 28242
rect -137 28208 -104 28242
rect -46 28208 -13 28242
rect 21 28208 54 28242
rect 112 28208 145 28242
rect 179 28208 212 28242
rect 270 28208 303 28242
rect 337 28208 370 28242
rect 428 28208 461 28242
rect 495 28208 528 28242
rect 586 28208 619 28242
rect 653 28208 686 28242
rect 744 28208 777 28242
rect 811 28208 844 28242
rect 902 28208 935 28242
rect 969 28208 1002 28242
rect 1060 28208 1093 28242
rect 1127 28208 1160 28242
rect 1218 28208 1251 28242
rect 1285 28208 1318 28242
rect 1376 28208 1409 28242
rect 1443 28208 1476 28242
rect 1534 28208 1567 28242
rect 1601 28208 1634 28242
rect 1760 28140 1794 28228
rect -1786 28106 -1679 28140
rect -1645 28106 -1611 28140
rect -1577 28106 -1543 28140
rect -1509 28106 -1475 28140
rect -1441 28106 -1407 28140
rect -1373 28106 -1339 28140
rect -1305 28106 -1271 28140
rect -1237 28106 -1203 28140
rect -1169 28106 -1135 28140
rect -1101 28106 -1067 28140
rect -1033 28106 -999 28140
rect -965 28109 -931 28140
rect -897 28109 -863 28140
rect -829 28109 -795 28140
rect -761 28109 -727 28140
rect -693 28109 -659 28140
rect -625 28109 -591 28140
rect -557 28109 -523 28140
rect -489 28109 -455 28140
rect -458 28106 -455 28109
rect -421 28106 -387 28140
rect -353 28106 -319 28140
rect -285 28106 -251 28140
rect -217 28106 -183 28140
rect -149 28106 -115 28140
rect -81 28106 -47 28140
rect -13 28106 21 28140
rect 55 28106 89 28140
rect 123 28106 157 28140
rect 191 28106 225 28140
rect 259 28106 293 28140
rect 327 28106 361 28140
rect 395 28106 429 28140
rect 463 28109 497 28140
rect 531 28109 565 28140
rect 599 28109 633 28140
rect 667 28109 701 28140
rect 735 28109 769 28140
rect 803 28109 837 28140
rect 871 28109 905 28140
rect 939 28109 973 28140
rect 1007 28109 1041 28140
rect 463 28106 474 28109
rect 1012 28106 1041 28109
rect 1075 28106 1109 28140
rect 1143 28106 1177 28140
rect 1211 28106 1245 28140
rect 1279 28106 1313 28140
rect 1347 28106 1381 28140
rect 1415 28106 1449 28140
rect 1483 28106 1517 28140
rect 1551 28106 1585 28140
rect 1619 28106 1653 28140
rect 1687 28106 1794 28140
rect -1012 27932 -996 28106
rect -458 27932 -442 28106
rect 458 27932 474 28106
rect 1012 27932 1028 28106
rect -1786 27898 -1679 27932
rect -1645 27898 -1611 27932
rect -1577 27898 -1543 27932
rect -1509 27898 -1475 27932
rect -1441 27898 -1407 27932
rect -1373 27898 -1339 27932
rect -1305 27898 -1271 27932
rect -1237 27898 -1203 27932
rect -1169 27898 -1135 27932
rect -1101 27898 -1067 27932
rect -1033 27898 -999 27932
rect -458 27931 -455 27932
rect -965 27898 -931 27931
rect -897 27898 -863 27931
rect -829 27898 -795 27931
rect -761 27898 -727 27931
rect -693 27898 -659 27931
rect -625 27898 -591 27931
rect -557 27898 -523 27931
rect -489 27898 -455 27931
rect -421 27898 -387 27932
rect -353 27898 -319 27932
rect -285 27898 -251 27932
rect -217 27898 -183 27932
rect -149 27898 -115 27932
rect -81 27898 -47 27932
rect -13 27898 21 27932
rect 55 27898 89 27932
rect 123 27898 157 27932
rect 191 27898 225 27932
rect 259 27898 293 27932
rect 327 27898 361 27932
rect 395 27898 429 27932
rect 463 27931 474 27932
rect 1012 27931 1041 27932
rect 463 27898 497 27931
rect 531 27898 565 27931
rect 599 27898 633 27931
rect 667 27898 701 27931
rect 735 27898 769 27931
rect 803 27898 837 27931
rect 871 27898 905 27931
rect 939 27898 973 27931
rect 1007 27898 1041 27931
rect 1075 27898 1109 27932
rect 1143 27898 1177 27932
rect 1211 27898 1245 27932
rect 1279 27898 1313 27932
rect 1347 27898 1381 27932
rect 1415 27898 1449 27932
rect 1483 27898 1517 27932
rect 1551 27898 1585 27932
rect 1619 27898 1653 27932
rect 1687 27898 1794 27932
rect -1786 27810 -1752 27898
rect -1626 27796 -1593 27830
rect -1559 27796 -1526 27830
rect -1468 27796 -1435 27830
rect -1401 27796 -1368 27830
rect -1310 27796 -1277 27830
rect -1243 27796 -1210 27830
rect -1152 27796 -1119 27830
rect -1085 27796 -1052 27830
rect -994 27796 -961 27830
rect -927 27796 -894 27830
rect -836 27796 -803 27830
rect -769 27796 -736 27830
rect -678 27796 -645 27830
rect -611 27796 -578 27830
rect -520 27796 -487 27830
rect -453 27796 -420 27830
rect -362 27796 -329 27830
rect -295 27796 -262 27830
rect -204 27796 -171 27830
rect -137 27796 -104 27830
rect -46 27796 -13 27830
rect 21 27796 54 27830
rect 112 27796 145 27830
rect 179 27796 212 27830
rect 270 27796 303 27830
rect 337 27796 370 27830
rect 428 27796 461 27830
rect 495 27796 528 27830
rect 586 27796 619 27830
rect 653 27796 686 27830
rect 744 27796 777 27830
rect 811 27796 844 27830
rect 902 27796 935 27830
rect 969 27796 1002 27830
rect 1060 27796 1093 27830
rect 1127 27796 1160 27830
rect 1218 27796 1251 27830
rect 1285 27796 1318 27830
rect 1376 27796 1409 27830
rect 1443 27796 1476 27830
rect 1534 27796 1567 27830
rect 1601 27796 1634 27830
rect 1760 27810 1794 27898
rect -1786 27742 -1752 27776
rect -1786 27674 -1752 27708
rect -1786 27606 -1752 27640
rect -1786 27538 -1752 27572
rect -1786 27470 -1752 27504
rect -1786 27402 -1752 27436
rect -1786 27334 -1752 27368
rect -1786 27266 -1752 27300
rect -1786 27198 -1752 27232
rect -1786 27130 -1752 27164
rect -1786 27062 -1752 27096
rect -1786 26994 -1752 27028
rect -1786 26926 -1752 26960
rect -1786 26858 -1752 26892
rect -1786 26790 -1752 26824
rect -1786 26722 -1752 26756
rect -1672 27734 -1638 27753
rect -1672 27662 -1638 27674
rect -1672 27590 -1638 27606
rect -1672 27518 -1638 27538
rect -1672 27446 -1638 27470
rect -1672 27374 -1638 27402
rect -1672 27302 -1638 27334
rect -1672 27232 -1638 27266
rect -1672 27164 -1638 27196
rect -1672 27096 -1638 27124
rect -1672 27028 -1638 27052
rect -1672 26960 -1638 26980
rect -1672 26892 -1638 26908
rect -1672 26824 -1638 26836
rect -1672 26745 -1638 26764
rect -1514 27734 -1480 27753
rect -1514 27662 -1480 27674
rect -1514 27590 -1480 27606
rect -1514 27518 -1480 27538
rect -1514 27446 -1480 27470
rect -1514 27374 -1480 27402
rect -1514 27302 -1480 27334
rect -1514 27232 -1480 27266
rect -1514 27164 -1480 27196
rect -1514 27096 -1480 27124
rect -1514 27028 -1480 27052
rect -1514 26960 -1480 26980
rect -1514 26892 -1480 26908
rect -1514 26824 -1480 26836
rect -1514 26745 -1480 26764
rect -1356 27734 -1322 27753
rect -1356 27662 -1322 27674
rect -1356 27590 -1322 27606
rect -1356 27518 -1322 27538
rect -1356 27446 -1322 27470
rect -1356 27374 -1322 27402
rect -1356 27302 -1322 27334
rect -1356 27232 -1322 27266
rect -1356 27164 -1322 27196
rect -1356 27096 -1322 27124
rect -1356 27028 -1322 27052
rect -1356 26960 -1322 26980
rect -1356 26892 -1322 26908
rect -1356 26824 -1322 26836
rect -1356 26745 -1322 26764
rect -1198 27734 -1164 27753
rect -1198 27662 -1164 27674
rect -1198 27590 -1164 27606
rect -1198 27518 -1164 27538
rect -1198 27446 -1164 27470
rect -1198 27374 -1164 27402
rect -1198 27302 -1164 27334
rect -1198 27232 -1164 27266
rect -1198 27164 -1164 27196
rect -1198 27096 -1164 27124
rect -1198 27028 -1164 27052
rect -1198 26960 -1164 26980
rect -1198 26892 -1164 26908
rect -1198 26824 -1164 26836
rect -1198 26745 -1164 26764
rect -1040 27734 -1006 27753
rect -1040 27662 -1006 27674
rect -1040 27590 -1006 27606
rect -1040 27518 -1006 27538
rect -1040 27446 -1006 27470
rect -1040 27374 -1006 27402
rect -1040 27302 -1006 27334
rect -1040 27232 -1006 27266
rect -1040 27164 -1006 27196
rect -1040 27096 -1006 27124
rect -1040 27028 -1006 27052
rect -1040 26960 -1006 26980
rect -1040 26892 -1006 26908
rect -1040 26824 -1006 26836
rect -1040 26745 -1006 26764
rect -882 27734 -848 27753
rect -882 27662 -848 27674
rect -882 27590 -848 27606
rect -882 27518 -848 27538
rect -882 27446 -848 27470
rect -882 27374 -848 27402
rect -882 27302 -848 27334
rect -882 27232 -848 27266
rect -882 27164 -848 27196
rect -882 27096 -848 27124
rect -882 27028 -848 27052
rect -882 26960 -848 26980
rect -882 26892 -848 26908
rect -882 26824 -848 26836
rect -882 26745 -848 26764
rect -724 27734 -690 27753
rect -724 27662 -690 27674
rect -724 27590 -690 27606
rect -724 27518 -690 27538
rect -724 27446 -690 27470
rect -724 27374 -690 27402
rect -724 27302 -690 27334
rect -724 27232 -690 27266
rect -724 27164 -690 27196
rect -724 27096 -690 27124
rect -724 27028 -690 27052
rect -724 26960 -690 26980
rect -724 26892 -690 26908
rect -724 26824 -690 26836
rect -724 26745 -690 26764
rect -566 27734 -532 27753
rect -566 27662 -532 27674
rect -566 27590 -532 27606
rect -566 27518 -532 27538
rect -566 27446 -532 27470
rect -566 27374 -532 27402
rect -566 27302 -532 27334
rect -566 27232 -532 27266
rect -566 27164 -532 27196
rect -566 27096 -532 27124
rect -566 27028 -532 27052
rect -566 26960 -532 26980
rect -566 26892 -532 26908
rect -566 26824 -532 26836
rect -566 26745 -532 26764
rect -408 27734 -374 27753
rect -408 27662 -374 27674
rect -408 27590 -374 27606
rect -408 27518 -374 27538
rect -408 27446 -374 27470
rect -408 27374 -374 27402
rect -408 27302 -374 27334
rect -408 27232 -374 27266
rect -408 27164 -374 27196
rect -408 27096 -374 27124
rect -408 27028 -374 27052
rect -408 26960 -374 26980
rect -408 26892 -374 26908
rect -408 26824 -374 26836
rect -408 26745 -374 26764
rect -250 27734 -216 27753
rect -250 27662 -216 27674
rect -250 27590 -216 27606
rect -250 27518 -216 27538
rect -250 27446 -216 27470
rect -250 27374 -216 27402
rect -250 27302 -216 27334
rect -250 27232 -216 27266
rect -250 27164 -216 27196
rect -250 27096 -216 27124
rect -250 27028 -216 27052
rect -250 26960 -216 26980
rect -250 26892 -216 26908
rect -250 26824 -216 26836
rect -250 26745 -216 26764
rect -92 27734 -58 27753
rect -92 27662 -58 27674
rect -92 27590 -58 27606
rect -92 27518 -58 27538
rect -92 27446 -58 27470
rect -92 27374 -58 27402
rect -92 27302 -58 27334
rect -92 27232 -58 27266
rect -92 27164 -58 27196
rect -92 27096 -58 27124
rect -92 27028 -58 27052
rect -92 26960 -58 26980
rect -92 26892 -58 26908
rect -92 26824 -58 26836
rect -92 26745 -58 26764
rect 66 27734 100 27753
rect 66 27662 100 27674
rect 66 27590 100 27606
rect 66 27518 100 27538
rect 66 27446 100 27470
rect 66 27374 100 27402
rect 66 27302 100 27334
rect 66 27232 100 27266
rect 66 27164 100 27196
rect 66 27096 100 27124
rect 66 27028 100 27052
rect 66 26960 100 26980
rect 66 26892 100 26908
rect 66 26824 100 26836
rect 66 26745 100 26764
rect 224 27734 258 27753
rect 224 27662 258 27674
rect 224 27590 258 27606
rect 224 27518 258 27538
rect 224 27446 258 27470
rect 224 27374 258 27402
rect 224 27302 258 27334
rect 224 27232 258 27266
rect 224 27164 258 27196
rect 224 27096 258 27124
rect 224 27028 258 27052
rect 224 26960 258 26980
rect 224 26892 258 26908
rect 224 26824 258 26836
rect 224 26745 258 26764
rect 382 27734 416 27753
rect 382 27662 416 27674
rect 382 27590 416 27606
rect 382 27518 416 27538
rect 382 27446 416 27470
rect 382 27374 416 27402
rect 382 27302 416 27334
rect 382 27232 416 27266
rect 382 27164 416 27196
rect 382 27096 416 27124
rect 382 27028 416 27052
rect 382 26960 416 26980
rect 382 26892 416 26908
rect 382 26824 416 26836
rect 382 26745 416 26764
rect 540 27734 574 27753
rect 540 27662 574 27674
rect 540 27590 574 27606
rect 540 27518 574 27538
rect 540 27446 574 27470
rect 540 27374 574 27402
rect 540 27302 574 27334
rect 540 27232 574 27266
rect 540 27164 574 27196
rect 540 27096 574 27124
rect 540 27028 574 27052
rect 540 26960 574 26980
rect 540 26892 574 26908
rect 540 26824 574 26836
rect 540 26745 574 26764
rect 698 27734 732 27753
rect 698 27662 732 27674
rect 698 27590 732 27606
rect 698 27518 732 27538
rect 698 27446 732 27470
rect 698 27374 732 27402
rect 698 27302 732 27334
rect 698 27232 732 27266
rect 698 27164 732 27196
rect 698 27096 732 27124
rect 698 27028 732 27052
rect 698 26960 732 26980
rect 698 26892 732 26908
rect 698 26824 732 26836
rect 698 26745 732 26764
rect 856 27734 890 27753
rect 856 27662 890 27674
rect 856 27590 890 27606
rect 856 27518 890 27538
rect 856 27446 890 27470
rect 856 27374 890 27402
rect 856 27302 890 27334
rect 856 27232 890 27266
rect 856 27164 890 27196
rect 856 27096 890 27124
rect 856 27028 890 27052
rect 856 26960 890 26980
rect 856 26892 890 26908
rect 856 26824 890 26836
rect 856 26745 890 26764
rect 1014 27734 1048 27753
rect 1014 27662 1048 27674
rect 1014 27590 1048 27606
rect 1014 27518 1048 27538
rect 1014 27446 1048 27470
rect 1014 27374 1048 27402
rect 1014 27302 1048 27334
rect 1014 27232 1048 27266
rect 1014 27164 1048 27196
rect 1014 27096 1048 27124
rect 1014 27028 1048 27052
rect 1014 26960 1048 26980
rect 1014 26892 1048 26908
rect 1014 26824 1048 26836
rect 1014 26745 1048 26764
rect 1172 27734 1206 27753
rect 1172 27662 1206 27674
rect 1172 27590 1206 27606
rect 1172 27518 1206 27538
rect 1172 27446 1206 27470
rect 1172 27374 1206 27402
rect 1172 27302 1206 27334
rect 1172 27232 1206 27266
rect 1172 27164 1206 27196
rect 1172 27096 1206 27124
rect 1172 27028 1206 27052
rect 1172 26960 1206 26980
rect 1172 26892 1206 26908
rect 1172 26824 1206 26836
rect 1172 26745 1206 26764
rect 1330 27734 1364 27753
rect 1330 27662 1364 27674
rect 1330 27590 1364 27606
rect 1330 27518 1364 27538
rect 1330 27446 1364 27470
rect 1330 27374 1364 27402
rect 1330 27302 1364 27334
rect 1330 27232 1364 27266
rect 1330 27164 1364 27196
rect 1330 27096 1364 27124
rect 1330 27028 1364 27052
rect 1330 26960 1364 26980
rect 1330 26892 1364 26908
rect 1330 26824 1364 26836
rect 1330 26745 1364 26764
rect 1488 27734 1522 27753
rect 1488 27662 1522 27674
rect 1488 27590 1522 27606
rect 1488 27518 1522 27538
rect 1488 27446 1522 27470
rect 1488 27374 1522 27402
rect 1488 27302 1522 27334
rect 1488 27232 1522 27266
rect 1488 27164 1522 27196
rect 1488 27096 1522 27124
rect 1488 27028 1522 27052
rect 1488 26960 1522 26980
rect 1488 26892 1522 26908
rect 1488 26824 1522 26836
rect 1488 26745 1522 26764
rect 1646 27734 1680 27753
rect 1646 27662 1680 27674
rect 1646 27590 1680 27606
rect 1646 27518 1680 27538
rect 1646 27446 1680 27470
rect 1646 27374 1680 27402
rect 1646 27302 1680 27334
rect 1646 27232 1680 27266
rect 1646 27164 1680 27196
rect 1646 27096 1680 27124
rect 1646 27028 1680 27052
rect 1646 26960 1680 26980
rect 1646 26892 1680 26908
rect 1646 26824 1680 26836
rect 1646 26745 1680 26764
rect 1760 27742 1794 27776
rect 1760 27674 1794 27708
rect 1760 27606 1794 27640
rect 1760 27538 1794 27572
rect 1760 27470 1794 27504
rect 1760 27402 1794 27436
rect 1760 27334 1794 27368
rect 1760 27266 1794 27300
rect 1760 27198 1794 27232
rect 1760 27130 1794 27164
rect 1760 27062 1794 27096
rect 1760 26994 1794 27028
rect 1760 26926 1794 26960
rect 1760 26858 1794 26892
rect 1760 26790 1794 26824
rect 1760 26722 1794 26756
rect -1786 26600 -1752 26688
rect -1626 26668 -1593 26702
rect -1559 26668 -1526 26702
rect -1468 26668 -1435 26702
rect -1401 26668 -1368 26702
rect -1310 26668 -1277 26702
rect -1243 26668 -1210 26702
rect -1152 26668 -1119 26702
rect -1085 26668 -1052 26702
rect -994 26668 -961 26702
rect -927 26668 -894 26702
rect -836 26668 -803 26702
rect -769 26668 -736 26702
rect -678 26668 -645 26702
rect -611 26668 -578 26702
rect -520 26668 -487 26702
rect -453 26668 -420 26702
rect -362 26668 -329 26702
rect -295 26668 -262 26702
rect -204 26668 -171 26702
rect -137 26668 -104 26702
rect -46 26668 -13 26702
rect 21 26668 54 26702
rect 112 26668 145 26702
rect 179 26668 212 26702
rect 270 26668 303 26702
rect 337 26668 370 26702
rect 428 26668 461 26702
rect 495 26668 528 26702
rect 586 26668 619 26702
rect 653 26668 686 26702
rect 744 26668 777 26702
rect 811 26668 844 26702
rect 902 26668 935 26702
rect 969 26668 1002 26702
rect 1060 26668 1093 26702
rect 1127 26668 1160 26702
rect 1218 26668 1251 26702
rect 1285 26668 1318 26702
rect 1376 26668 1409 26702
rect 1443 26668 1476 26702
rect 1534 26668 1567 26702
rect 1601 26668 1634 26702
rect 1760 26600 1794 26688
rect -1786 26566 -1679 26600
rect -1645 26566 -1611 26600
rect -1577 26566 -1543 26600
rect -1509 26566 -1475 26600
rect -1441 26566 -1407 26600
rect -1373 26566 -1339 26600
rect -1305 26566 -1271 26600
rect -1237 26566 -1203 26600
rect -1169 26566 -1135 26600
rect -1101 26566 -1067 26600
rect -1033 26566 -999 26600
rect -965 26566 -931 26600
rect -897 26566 -863 26600
rect -829 26566 -795 26600
rect -761 26566 -727 26600
rect -693 26566 -659 26600
rect -625 26566 -591 26600
rect -557 26566 -523 26600
rect -489 26566 -455 26600
rect -421 26566 -387 26600
rect -353 26566 -319 26600
rect -285 26566 -251 26600
rect -217 26566 -183 26600
rect -149 26566 -115 26600
rect -81 26566 -47 26600
rect -13 26566 21 26600
rect 55 26566 89 26600
rect 123 26566 157 26600
rect 191 26566 225 26600
rect 259 26566 293 26600
rect 327 26566 361 26600
rect 395 26566 429 26600
rect 463 26566 497 26600
rect 531 26566 565 26600
rect 599 26566 633 26600
rect 667 26566 701 26600
rect 735 26566 769 26600
rect 803 26566 837 26600
rect 871 26566 905 26600
rect 939 26566 973 26600
rect 1007 26566 1041 26600
rect 1075 26566 1109 26600
rect 1143 26566 1177 26600
rect 1211 26566 1245 26600
rect 1279 26566 1313 26600
rect 1347 26566 1381 26600
rect 1415 26566 1449 26600
rect 1483 26566 1517 26600
rect 1551 26566 1585 26600
rect 1619 26566 1653 26600
rect 1687 26566 1794 26600
rect -685 26321 -562 26355
rect -528 26321 -494 26355
rect -460 26321 -426 26355
rect -392 26321 -358 26355
rect -324 26321 -306 26355
rect -256 26321 -234 26355
rect -188 26321 -162 26355
rect -120 26321 -90 26355
rect -52 26321 -18 26355
rect 16 26321 50 26355
rect 88 26321 118 26355
rect 160 26321 186 26355
rect 232 26321 254 26355
rect 304 26321 322 26355
rect 356 26321 390 26355
rect 424 26321 458 26355
rect 492 26321 526 26355
rect 560 26321 683 26355
rect -685 26242 -651 26321
rect -525 26219 -492 26253
rect -458 26219 -425 26253
rect -367 26219 -334 26253
rect -300 26219 -267 26253
rect -209 26219 -176 26253
rect -142 26219 -109 26253
rect -51 26219 -18 26253
rect 16 26219 49 26253
rect 107 26219 140 26253
rect 174 26219 207 26253
rect 265 26219 298 26253
rect 332 26219 365 26253
rect 423 26219 456 26253
rect 490 26219 523 26253
rect 649 26242 683 26321
rect -685 26174 -651 26208
rect -685 26106 -651 26140
rect -685 26038 -651 26072
rect -685 25970 -651 26004
rect -685 25902 -651 25936
rect -685 25834 -651 25868
rect -685 25766 -651 25800
rect -685 25698 -651 25732
rect -685 25630 -651 25664
rect -685 25562 -651 25596
rect -685 25494 -651 25528
rect -685 25426 -651 25460
rect -685 25358 -651 25392
rect -685 25290 -651 25324
rect -685 25222 -651 25256
rect -685 25154 -651 25188
rect -571 26166 -537 26185
rect -571 26094 -537 26106
rect -571 26022 -537 26038
rect -571 25950 -537 25970
rect -571 25878 -537 25902
rect -571 25806 -537 25834
rect -571 25734 -537 25766
rect -571 25664 -537 25698
rect -571 25596 -537 25628
rect -571 25528 -537 25556
rect -571 25460 -537 25484
rect -571 25392 -537 25412
rect -571 25324 -537 25340
rect -571 25256 -537 25268
rect -571 25177 -537 25196
rect -413 26166 -379 26185
rect -413 26094 -379 26106
rect -413 26022 -379 26038
rect -413 25950 -379 25970
rect -413 25878 -379 25902
rect -413 25806 -379 25834
rect -413 25734 -379 25766
rect -413 25664 -379 25698
rect -413 25596 -379 25628
rect -413 25528 -379 25556
rect -413 25460 -379 25484
rect -413 25392 -379 25412
rect -413 25324 -379 25340
rect -413 25256 -379 25268
rect -413 25177 -379 25196
rect -255 26166 -221 26185
rect -255 26094 -221 26106
rect -255 26022 -221 26038
rect -255 25950 -221 25970
rect -255 25878 -221 25902
rect -255 25806 -221 25834
rect -255 25734 -221 25766
rect -255 25664 -221 25698
rect -255 25596 -221 25628
rect -255 25528 -221 25556
rect -255 25460 -221 25484
rect -255 25392 -221 25412
rect -255 25324 -221 25340
rect -255 25256 -221 25268
rect -255 25177 -221 25196
rect -97 26166 -63 26185
rect -97 26094 -63 26106
rect -97 26022 -63 26038
rect -97 25950 -63 25970
rect -97 25878 -63 25902
rect -97 25806 -63 25834
rect -97 25734 -63 25766
rect -97 25664 -63 25698
rect -97 25596 -63 25628
rect -97 25528 -63 25556
rect -97 25460 -63 25484
rect -97 25392 -63 25412
rect -97 25324 -63 25340
rect -97 25256 -63 25268
rect -97 25177 -63 25196
rect 61 26166 95 26185
rect 61 26094 95 26106
rect 61 26022 95 26038
rect 61 25950 95 25970
rect 61 25878 95 25902
rect 61 25806 95 25834
rect 61 25734 95 25766
rect 61 25664 95 25698
rect 61 25596 95 25628
rect 61 25528 95 25556
rect 61 25460 95 25484
rect 61 25392 95 25412
rect 61 25324 95 25340
rect 61 25256 95 25268
rect 61 25177 95 25196
rect 219 26166 253 26185
rect 219 26094 253 26106
rect 219 26022 253 26038
rect 219 25950 253 25970
rect 219 25878 253 25902
rect 219 25806 253 25834
rect 219 25734 253 25766
rect 219 25664 253 25698
rect 219 25596 253 25628
rect 219 25528 253 25556
rect 219 25460 253 25484
rect 219 25392 253 25412
rect 219 25324 253 25340
rect 219 25256 253 25268
rect 219 25177 253 25196
rect 377 26166 411 26185
rect 377 26094 411 26106
rect 377 26022 411 26038
rect 377 25950 411 25970
rect 377 25878 411 25902
rect 377 25806 411 25834
rect 377 25734 411 25766
rect 377 25664 411 25698
rect 377 25596 411 25628
rect 377 25528 411 25556
rect 377 25460 411 25484
rect 377 25392 411 25412
rect 377 25324 411 25340
rect 377 25256 411 25268
rect 377 25177 411 25196
rect 535 26166 569 26185
rect 535 26094 569 26106
rect 535 26022 569 26038
rect 535 25950 569 25970
rect 535 25878 569 25902
rect 535 25806 569 25834
rect 535 25734 569 25766
rect 535 25664 569 25698
rect 535 25596 569 25628
rect 535 25528 569 25556
rect 535 25460 569 25484
rect 535 25392 569 25412
rect 535 25324 569 25340
rect 535 25256 569 25268
rect 535 25177 569 25196
rect 649 26174 683 26208
rect 649 26106 683 26140
rect 649 26038 683 26072
rect 649 25970 683 26004
rect 649 25902 683 25936
rect 649 25834 683 25868
rect 649 25766 683 25800
rect 649 25698 683 25732
rect 649 25630 683 25664
rect 649 25562 683 25596
rect 649 25494 683 25528
rect 649 25426 683 25460
rect 649 25358 683 25392
rect 649 25290 683 25324
rect 649 25222 683 25256
rect 649 25154 683 25188
rect -685 25041 -651 25120
rect -525 25109 -492 25143
rect -458 25109 -425 25143
rect -367 25109 -334 25143
rect -300 25109 -267 25143
rect -209 25109 -176 25143
rect -142 25109 -109 25143
rect -51 25109 -18 25143
rect 16 25109 49 25143
rect 107 25109 140 25143
rect 174 25109 207 25143
rect 265 25109 298 25143
rect 332 25109 365 25143
rect 423 25109 456 25143
rect 490 25109 523 25143
rect 649 25041 683 25120
rect -685 25007 -562 25041
rect -528 25007 -494 25041
rect -460 25007 -426 25041
rect -392 25007 -358 25041
rect -324 25007 -306 25041
rect -256 25007 -234 25041
rect -188 25007 -162 25041
rect -120 25007 -90 25041
rect -52 25007 -18 25041
rect 16 25007 50 25041
rect 88 25007 118 25041
rect 160 25007 186 25041
rect 232 25007 254 25041
rect 304 25007 322 25041
rect 356 25007 390 25041
rect 424 25007 458 25041
rect 492 25007 526 25041
rect 560 25007 683 25041
rect -685 24801 -562 24835
rect -528 24801 -494 24835
rect -460 24801 -426 24835
rect -392 24801 -358 24835
rect -324 24801 -306 24835
rect -256 24801 -234 24835
rect -188 24801 -162 24835
rect -120 24801 -90 24835
rect -52 24801 -18 24835
rect 16 24801 50 24835
rect 88 24801 118 24835
rect 160 24801 186 24835
rect 232 24801 254 24835
rect 304 24801 322 24835
rect 356 24801 390 24835
rect 424 24801 458 24835
rect 492 24801 526 24835
rect 560 24801 683 24835
rect -685 24722 -651 24801
rect -525 24699 -492 24733
rect -458 24699 -425 24733
rect -367 24699 -334 24733
rect -300 24699 -267 24733
rect -209 24699 -176 24733
rect -142 24699 -109 24733
rect -51 24699 -18 24733
rect 16 24699 49 24733
rect 107 24699 140 24733
rect 174 24699 207 24733
rect 265 24699 298 24733
rect 332 24699 365 24733
rect 423 24699 456 24733
rect 490 24699 523 24733
rect 649 24722 683 24801
rect -685 24654 -651 24688
rect -685 24586 -651 24620
rect -685 24518 -651 24552
rect -685 24450 -651 24484
rect -685 24382 -651 24416
rect -685 24314 -651 24348
rect -685 24246 -651 24280
rect -685 24178 -651 24212
rect -685 24110 -651 24144
rect -685 24042 -651 24076
rect -685 23974 -651 24008
rect -685 23906 -651 23940
rect -685 23838 -651 23872
rect -685 23770 -651 23804
rect -685 23702 -651 23736
rect -685 23634 -651 23668
rect -571 24646 -537 24665
rect -571 24574 -537 24586
rect -571 24502 -537 24518
rect -571 24430 -537 24450
rect -571 24358 -537 24382
rect -571 24286 -537 24314
rect -571 24214 -537 24246
rect -571 24144 -537 24178
rect -571 24076 -537 24108
rect -571 24008 -537 24036
rect -571 23940 -537 23964
rect -571 23872 -537 23892
rect -571 23804 -537 23820
rect -571 23736 -537 23748
rect -571 23657 -537 23676
rect -413 24646 -379 24665
rect -413 24574 -379 24586
rect -413 24502 -379 24518
rect -413 24430 -379 24450
rect -413 24358 -379 24382
rect -413 24286 -379 24314
rect -413 24214 -379 24246
rect -413 24144 -379 24178
rect -413 24076 -379 24108
rect -413 24008 -379 24036
rect -413 23940 -379 23964
rect -413 23872 -379 23892
rect -413 23804 -379 23820
rect -413 23736 -379 23748
rect -413 23657 -379 23676
rect -255 24646 -221 24665
rect -255 24574 -221 24586
rect -255 24502 -221 24518
rect -255 24430 -221 24450
rect -255 24358 -221 24382
rect -255 24286 -221 24314
rect -255 24214 -221 24246
rect -255 24144 -221 24178
rect -255 24076 -221 24108
rect -255 24008 -221 24036
rect -255 23940 -221 23964
rect -255 23872 -221 23892
rect -255 23804 -221 23820
rect -255 23736 -221 23748
rect -255 23657 -221 23676
rect -97 24646 -63 24665
rect -97 24574 -63 24586
rect -97 24502 -63 24518
rect -97 24430 -63 24450
rect -97 24358 -63 24382
rect -97 24286 -63 24314
rect -97 24214 -63 24246
rect -97 24144 -63 24178
rect -97 24076 -63 24108
rect -97 24008 -63 24036
rect -97 23940 -63 23964
rect -97 23872 -63 23892
rect -97 23804 -63 23820
rect -97 23736 -63 23748
rect -97 23657 -63 23676
rect 61 24646 95 24665
rect 61 24574 95 24586
rect 61 24502 95 24518
rect 61 24430 95 24450
rect 61 24358 95 24382
rect 61 24286 95 24314
rect 61 24214 95 24246
rect 61 24144 95 24178
rect 61 24076 95 24108
rect 61 24008 95 24036
rect 61 23940 95 23964
rect 61 23872 95 23892
rect 61 23804 95 23820
rect 61 23736 95 23748
rect 61 23657 95 23676
rect 219 24646 253 24665
rect 219 24574 253 24586
rect 219 24502 253 24518
rect 219 24430 253 24450
rect 219 24358 253 24382
rect 219 24286 253 24314
rect 219 24214 253 24246
rect 219 24144 253 24178
rect 219 24076 253 24108
rect 219 24008 253 24036
rect 219 23940 253 23964
rect 219 23872 253 23892
rect 219 23804 253 23820
rect 219 23736 253 23748
rect 219 23657 253 23676
rect 377 24646 411 24665
rect 377 24574 411 24586
rect 377 24502 411 24518
rect 377 24430 411 24450
rect 377 24358 411 24382
rect 377 24286 411 24314
rect 377 24214 411 24246
rect 377 24144 411 24178
rect 377 24076 411 24108
rect 377 24008 411 24036
rect 377 23940 411 23964
rect 377 23872 411 23892
rect 377 23804 411 23820
rect 377 23736 411 23748
rect 377 23657 411 23676
rect 535 24646 569 24665
rect 535 24574 569 24586
rect 535 24502 569 24518
rect 535 24430 569 24450
rect 535 24358 569 24382
rect 535 24286 569 24314
rect 535 24214 569 24246
rect 535 24144 569 24178
rect 535 24076 569 24108
rect 535 24008 569 24036
rect 535 23940 569 23964
rect 535 23872 569 23892
rect 535 23804 569 23820
rect 535 23736 569 23748
rect 535 23657 569 23676
rect 649 24654 683 24688
rect 649 24586 683 24620
rect 649 24518 683 24552
rect 649 24450 683 24484
rect 649 24382 683 24416
rect 649 24314 683 24348
rect 649 24246 683 24280
rect 649 24178 683 24212
rect 649 24110 683 24144
rect 649 24042 683 24076
rect 649 23974 683 24008
rect 649 23906 683 23940
rect 649 23838 683 23872
rect 649 23770 683 23804
rect 649 23702 683 23736
rect 649 23634 683 23668
rect -685 23521 -651 23600
rect -525 23589 -492 23623
rect -458 23589 -425 23623
rect -367 23589 -334 23623
rect -300 23589 -267 23623
rect -209 23589 -176 23623
rect -142 23589 -109 23623
rect -51 23589 -18 23623
rect 16 23589 49 23623
rect 107 23589 140 23623
rect 174 23589 207 23623
rect 265 23589 298 23623
rect 332 23589 365 23623
rect 423 23589 456 23623
rect 490 23589 523 23623
rect 649 23521 683 23600
rect -685 23487 -562 23521
rect -528 23487 -494 23521
rect -460 23487 -426 23521
rect -392 23487 -358 23521
rect -324 23487 -306 23521
rect -256 23487 -234 23521
rect -188 23487 -162 23521
rect -120 23487 -90 23521
rect -52 23487 -18 23521
rect 16 23487 50 23521
rect 88 23487 118 23521
rect 160 23487 186 23521
rect 232 23487 254 23521
rect 304 23487 322 23521
rect 356 23487 390 23521
rect 424 23487 458 23521
rect 492 23487 526 23521
rect 560 23487 683 23521
rect -1676 23280 -1578 23314
rect -1544 23280 -1510 23314
rect -1476 23280 -1442 23314
rect -1408 23280 -1374 23314
rect -1340 23280 -1306 23314
rect -1272 23280 -1238 23314
rect -1204 23280 -1170 23314
rect -1136 23280 -1102 23314
rect -1068 23280 -1034 23314
rect -1000 23280 -966 23314
rect -932 23280 -898 23314
rect -864 23280 -830 23314
rect -772 23280 -762 23314
rect -700 23280 -694 23314
rect -628 23280 -626 23314
rect -592 23280 -590 23314
rect -524 23280 -518 23314
rect -456 23280 -446 23314
rect -388 23280 -374 23314
rect -320 23280 -302 23314
rect -252 23280 -230 23314
rect -184 23280 -158 23314
rect -116 23280 -86 23314
rect -48 23280 -14 23314
rect 20 23280 54 23314
rect 92 23280 122 23314
rect 164 23280 190 23314
rect 236 23280 258 23314
rect 308 23280 326 23314
rect 380 23280 394 23314
rect 452 23280 462 23314
rect 524 23280 530 23314
rect 596 23280 598 23314
rect 632 23280 634 23314
rect 700 23280 706 23314
rect 768 23280 778 23314
rect 836 23280 870 23314
rect 904 23280 938 23314
rect 972 23280 1006 23314
rect 1040 23280 1074 23314
rect 1108 23280 1142 23314
rect 1176 23280 1210 23314
rect 1244 23280 1278 23314
rect 1312 23280 1346 23314
rect 1380 23280 1414 23314
rect 1448 23280 1482 23314
rect 1516 23280 1550 23314
rect 1584 23280 1682 23314
rect -1676 23201 -1642 23280
rect -1516 23178 -1469 23212
rect -1433 23178 -1399 23212
rect -1363 23178 -1316 23212
rect -1258 23178 -1211 23212
rect -1175 23178 -1141 23212
rect -1105 23178 -1058 23212
rect -1000 23178 -953 23212
rect -917 23178 -883 23212
rect -847 23178 -800 23212
rect -742 23178 -695 23212
rect -659 23178 -625 23212
rect -589 23178 -542 23212
rect -484 23178 -437 23212
rect -401 23178 -367 23212
rect -331 23178 -284 23212
rect -226 23178 -179 23212
rect -143 23178 -109 23212
rect -73 23178 -26 23212
rect 32 23178 79 23212
rect 115 23178 149 23212
rect 185 23178 232 23212
rect 290 23178 337 23212
rect 373 23178 407 23212
rect 443 23178 490 23212
rect 548 23178 595 23212
rect 631 23178 665 23212
rect 701 23178 748 23212
rect 806 23178 853 23212
rect 889 23178 923 23212
rect 959 23178 1006 23212
rect 1064 23178 1111 23212
rect 1147 23178 1181 23212
rect 1217 23178 1264 23212
rect 1322 23178 1369 23212
rect 1405 23178 1439 23212
rect 1475 23178 1522 23212
rect 1648 23201 1682 23280
rect -1676 23133 -1642 23167
rect -1676 23065 -1642 23099
rect -1676 22997 -1642 23031
rect -1676 22929 -1642 22963
rect -1676 22861 -1642 22895
rect -1676 22793 -1642 22827
rect -1676 22725 -1642 22759
rect -1676 22657 -1642 22691
rect -1676 22589 -1642 22623
rect -1676 22521 -1642 22555
rect -1676 22453 -1642 22487
rect -1676 22385 -1642 22419
rect -1676 22317 -1642 22351
rect -1676 22249 -1642 22283
rect -1676 22181 -1642 22215
rect -1676 22113 -1642 22147
rect -1562 23125 -1528 23144
rect -1562 23053 -1528 23065
rect -1562 22981 -1528 22997
rect -1562 22909 -1528 22929
rect -1562 22837 -1528 22861
rect -1562 22765 -1528 22793
rect -1562 22693 -1528 22725
rect -1562 22623 -1528 22657
rect -1562 22555 -1528 22587
rect -1562 22487 -1528 22515
rect -1562 22419 -1528 22443
rect -1562 22351 -1528 22371
rect -1562 22283 -1528 22299
rect -1562 22215 -1528 22227
rect -1562 22136 -1528 22155
rect -1304 23125 -1270 23144
rect -1304 23053 -1270 23065
rect -1304 22981 -1270 22997
rect -1304 22909 -1270 22929
rect -1304 22837 -1270 22861
rect -1304 22765 -1270 22793
rect -1304 22693 -1270 22725
rect -1304 22623 -1270 22657
rect -1304 22555 -1270 22587
rect -1304 22487 -1270 22515
rect -1304 22419 -1270 22443
rect -1304 22351 -1270 22371
rect -1304 22283 -1270 22299
rect -1304 22215 -1270 22227
rect -1304 22136 -1270 22155
rect -1046 23125 -1012 23144
rect -1046 23053 -1012 23065
rect -1046 22981 -1012 22997
rect -1046 22909 -1012 22929
rect -1046 22837 -1012 22861
rect -1046 22765 -1012 22793
rect -1046 22693 -1012 22725
rect -1046 22623 -1012 22657
rect -1046 22555 -1012 22587
rect -1046 22487 -1012 22515
rect -1046 22419 -1012 22443
rect -1046 22351 -1012 22371
rect -1046 22283 -1012 22299
rect -1046 22215 -1012 22227
rect -1046 22136 -1012 22155
rect -788 23125 -754 23144
rect -788 23053 -754 23065
rect -788 22981 -754 22997
rect -788 22909 -754 22929
rect -788 22837 -754 22861
rect -788 22765 -754 22793
rect -788 22693 -754 22725
rect -788 22623 -754 22657
rect -788 22555 -754 22587
rect -788 22487 -754 22515
rect -788 22419 -754 22443
rect -788 22351 -754 22371
rect -788 22283 -754 22299
rect -788 22215 -754 22227
rect -788 22136 -754 22155
rect -530 23125 -496 23144
rect -530 23053 -496 23065
rect -530 22981 -496 22997
rect -530 22909 -496 22929
rect -530 22837 -496 22861
rect -530 22765 -496 22793
rect -530 22693 -496 22725
rect -530 22623 -496 22657
rect -530 22555 -496 22587
rect -530 22487 -496 22515
rect -530 22419 -496 22443
rect -530 22351 -496 22371
rect -530 22283 -496 22299
rect -530 22215 -496 22227
rect -530 22136 -496 22155
rect -272 23125 -238 23144
rect -272 23053 -238 23065
rect -272 22981 -238 22997
rect -272 22909 -238 22929
rect -272 22837 -238 22861
rect -272 22765 -238 22793
rect -272 22693 -238 22725
rect -272 22623 -238 22657
rect -272 22555 -238 22587
rect -272 22487 -238 22515
rect -272 22419 -238 22443
rect -272 22351 -238 22371
rect -272 22283 -238 22299
rect -272 22215 -238 22227
rect -272 22136 -238 22155
rect -14 23125 20 23144
rect -14 23053 20 23065
rect -14 22981 20 22997
rect -14 22909 20 22929
rect -14 22837 20 22861
rect -14 22765 20 22793
rect -14 22693 20 22725
rect -14 22623 20 22657
rect -14 22555 20 22587
rect -14 22487 20 22515
rect -14 22419 20 22443
rect -14 22351 20 22371
rect -14 22283 20 22299
rect -14 22215 20 22227
rect -14 22136 20 22155
rect 244 23125 278 23144
rect 244 23053 278 23065
rect 244 22981 278 22997
rect 244 22909 278 22929
rect 244 22837 278 22861
rect 244 22765 278 22793
rect 244 22693 278 22725
rect 244 22623 278 22657
rect 244 22555 278 22587
rect 244 22487 278 22515
rect 244 22419 278 22443
rect 244 22351 278 22371
rect 244 22283 278 22299
rect 244 22215 278 22227
rect 244 22136 278 22155
rect 502 23125 536 23144
rect 502 23053 536 23065
rect 502 22981 536 22997
rect 502 22909 536 22929
rect 502 22837 536 22861
rect 502 22765 536 22793
rect 502 22693 536 22725
rect 502 22623 536 22657
rect 502 22555 536 22587
rect 502 22487 536 22515
rect 502 22419 536 22443
rect 502 22351 536 22371
rect 502 22283 536 22299
rect 502 22215 536 22227
rect 502 22136 536 22155
rect 760 23125 794 23144
rect 760 23053 794 23065
rect 760 22981 794 22997
rect 760 22909 794 22929
rect 760 22837 794 22861
rect 760 22765 794 22793
rect 760 22693 794 22725
rect 760 22623 794 22657
rect 760 22555 794 22587
rect 760 22487 794 22515
rect 760 22419 794 22443
rect 760 22351 794 22371
rect 760 22283 794 22299
rect 760 22215 794 22227
rect 760 22136 794 22155
rect 1018 23125 1052 23144
rect 1018 23053 1052 23065
rect 1018 22981 1052 22997
rect 1018 22909 1052 22929
rect 1018 22837 1052 22861
rect 1018 22765 1052 22793
rect 1018 22693 1052 22725
rect 1018 22623 1052 22657
rect 1018 22555 1052 22587
rect 1018 22487 1052 22515
rect 1018 22419 1052 22443
rect 1018 22351 1052 22371
rect 1018 22283 1052 22299
rect 1018 22215 1052 22227
rect 1018 22136 1052 22155
rect 1276 23125 1310 23144
rect 1276 23053 1310 23065
rect 1276 22981 1310 22997
rect 1276 22909 1310 22929
rect 1276 22837 1310 22861
rect 1276 22765 1310 22793
rect 1276 22693 1310 22725
rect 1276 22623 1310 22657
rect 1276 22555 1310 22587
rect 1276 22487 1310 22515
rect 1276 22419 1310 22443
rect 1276 22351 1310 22371
rect 1276 22283 1310 22299
rect 1276 22215 1310 22227
rect 1276 22136 1310 22155
rect 1534 23125 1568 23144
rect 1534 23053 1568 23065
rect 1534 22981 1568 22997
rect 1534 22909 1568 22929
rect 1534 22837 1568 22861
rect 1534 22765 1568 22793
rect 1534 22693 1568 22725
rect 1534 22623 1568 22657
rect 1534 22555 1568 22587
rect 1534 22487 1568 22515
rect 1534 22419 1568 22443
rect 1534 22351 1568 22371
rect 1534 22283 1568 22299
rect 1534 22215 1568 22227
rect 1534 22136 1568 22155
rect 1648 23133 1682 23167
rect 1648 23065 1682 23099
rect 1648 22997 1682 23031
rect 1648 22929 1682 22963
rect 1648 22861 1682 22895
rect 1648 22793 1682 22827
rect 1648 22725 1682 22759
rect 1648 22657 1682 22691
rect 1648 22589 1682 22623
rect 1648 22521 1682 22555
rect 1648 22453 1682 22487
rect 1648 22385 1682 22419
rect 1648 22317 1682 22351
rect 1648 22249 1682 22283
rect 1648 22181 1682 22215
rect 1648 22113 1682 22147
rect -1676 22000 -1642 22079
rect -1516 22068 -1469 22102
rect -1433 22068 -1399 22102
rect -1363 22068 -1316 22102
rect -1258 22068 -1211 22102
rect -1175 22068 -1141 22102
rect -1105 22068 -1058 22102
rect -1000 22068 -953 22102
rect -917 22068 -883 22102
rect -847 22068 -800 22102
rect -742 22068 -695 22102
rect -659 22068 -625 22102
rect -589 22068 -542 22102
rect -484 22068 -437 22102
rect -401 22068 -367 22102
rect -331 22068 -284 22102
rect -226 22068 -179 22102
rect -143 22068 -109 22102
rect -73 22068 -26 22102
rect 32 22068 79 22102
rect 115 22068 149 22102
rect 185 22068 232 22102
rect 290 22068 337 22102
rect 373 22068 407 22102
rect 443 22068 490 22102
rect 548 22068 595 22102
rect 631 22068 665 22102
rect 701 22068 748 22102
rect 806 22068 853 22102
rect 889 22068 923 22102
rect 959 22068 1006 22102
rect 1064 22068 1111 22102
rect 1147 22068 1181 22102
rect 1217 22068 1264 22102
rect 1322 22068 1369 22102
rect 1405 22068 1439 22102
rect 1475 22068 1522 22102
rect 1648 22000 1682 22079
rect -1676 21966 -1578 22000
rect -1544 21966 -1510 22000
rect -1476 21966 -1442 22000
rect -1408 21966 -1374 22000
rect -1340 21966 -1306 22000
rect -1272 21966 -1238 22000
rect -1204 21966 -1170 22000
rect -1136 21966 -1102 22000
rect -1068 21966 -1034 22000
rect -1000 21966 -966 22000
rect -932 21966 -898 22000
rect -864 21966 -830 22000
rect -772 21966 -762 22000
rect -700 21966 -694 22000
rect -628 21966 -626 22000
rect -592 21966 -590 22000
rect -524 21966 -518 22000
rect -456 21966 -446 22000
rect -388 21966 -374 22000
rect -320 21966 -302 22000
rect -252 21966 -230 22000
rect -184 21966 -158 22000
rect -116 21966 -86 22000
rect -48 21966 -14 22000
rect 20 21966 54 22000
rect 92 21966 122 22000
rect 164 21966 190 22000
rect 236 21966 258 22000
rect 308 21966 326 22000
rect 380 21966 394 22000
rect 452 21966 462 22000
rect 524 21966 530 22000
rect 596 21966 598 22000
rect 632 21966 634 22000
rect 700 21966 706 22000
rect 768 21966 778 22000
rect 836 21966 870 22000
rect 904 21966 938 22000
rect 972 21966 1006 22000
rect 1040 21966 1074 22000
rect 1108 21966 1142 22000
rect 1176 21966 1210 22000
rect 1244 21966 1278 22000
rect 1312 21966 1346 22000
rect 1380 21966 1414 22000
rect 1448 21966 1482 22000
rect 1516 21966 1550 22000
rect 1584 21966 1682 22000
rect -1936 21760 -1818 21794
rect -1784 21760 -1750 21794
rect -1716 21760 -1682 21794
rect -1648 21760 -1614 21794
rect -1580 21760 -1546 21794
rect -1512 21760 -1478 21794
rect -1444 21760 -1410 21794
rect -1376 21760 -1342 21794
rect -1308 21760 -1274 21794
rect -1240 21760 -1206 21794
rect -1172 21760 -1138 21794
rect -1104 21760 -1070 21794
rect -1036 21760 -1002 21794
rect -968 21760 -934 21794
rect -882 21760 -866 21794
rect -810 21760 -798 21794
rect -738 21760 -730 21794
rect -666 21760 -662 21794
rect -560 21760 -556 21794
rect -492 21760 -484 21794
rect -424 21760 -412 21794
rect -356 21760 -340 21794
rect -288 21760 -268 21794
rect -220 21760 -196 21794
rect -152 21760 -124 21794
rect -84 21760 -52 21794
rect -16 21760 18 21794
rect 54 21760 86 21794
rect 126 21760 154 21794
rect 198 21760 222 21794
rect 270 21760 290 21794
rect 342 21760 358 21794
rect 414 21760 426 21794
rect 486 21760 494 21794
rect 558 21760 562 21794
rect 664 21760 668 21794
rect 732 21760 740 21794
rect 800 21760 812 21794
rect 868 21760 884 21794
rect 936 21760 970 21794
rect 1004 21760 1038 21794
rect 1072 21760 1106 21794
rect 1140 21760 1174 21794
rect 1208 21760 1242 21794
rect 1276 21760 1310 21794
rect 1344 21760 1378 21794
rect 1412 21760 1446 21794
rect 1480 21760 1514 21794
rect 1548 21760 1582 21794
rect 1616 21760 1650 21794
rect 1684 21760 1718 21794
rect 1752 21760 1786 21794
rect 1820 21760 1938 21794
rect -1936 21681 -1902 21760
rect -1776 21658 -1729 21692
rect -1693 21658 -1659 21692
rect -1623 21658 -1576 21692
rect -1518 21658 -1471 21692
rect -1435 21658 -1401 21692
rect -1365 21658 -1318 21692
rect -1260 21658 -1213 21692
rect -1177 21658 -1143 21692
rect -1107 21658 -1060 21692
rect -1002 21658 -955 21692
rect -919 21658 -885 21692
rect -849 21658 -802 21692
rect -744 21658 -697 21692
rect -661 21658 -627 21692
rect -591 21658 -544 21692
rect -486 21658 -439 21692
rect -403 21658 -369 21692
rect -333 21658 -286 21692
rect -228 21658 -181 21692
rect -145 21658 -111 21692
rect -75 21658 -28 21692
rect 30 21658 77 21692
rect 113 21658 147 21692
rect 183 21658 230 21692
rect 288 21658 335 21692
rect 371 21658 405 21692
rect 441 21658 488 21692
rect 546 21658 593 21692
rect 629 21658 663 21692
rect 699 21658 746 21692
rect 804 21658 851 21692
rect 887 21658 921 21692
rect 957 21658 1004 21692
rect 1062 21658 1109 21692
rect 1145 21658 1179 21692
rect 1215 21658 1262 21692
rect 1320 21658 1367 21692
rect 1403 21658 1437 21692
rect 1473 21658 1520 21692
rect 1578 21658 1625 21692
rect 1661 21658 1695 21692
rect 1731 21658 1778 21692
rect 1904 21681 1938 21760
rect -1936 21613 -1902 21647
rect -1936 21545 -1902 21579
rect -1936 21477 -1902 21511
rect -1936 21409 -1902 21443
rect -1936 21341 -1902 21375
rect -1936 21273 -1902 21307
rect -1936 21205 -1902 21239
rect -1936 21137 -1902 21171
rect -1936 21069 -1902 21103
rect -1936 21001 -1902 21035
rect -1936 20933 -1902 20967
rect -1936 20865 -1902 20899
rect -1936 20797 -1902 20831
rect -1936 20729 -1902 20763
rect -1936 20661 -1902 20695
rect -1936 20593 -1902 20627
rect -1822 21605 -1788 21624
rect -1822 21533 -1788 21545
rect -1822 21461 -1788 21477
rect -1822 21389 -1788 21409
rect -1822 21317 -1788 21341
rect -1822 21245 -1788 21273
rect -1822 21173 -1788 21205
rect -1822 21103 -1788 21137
rect -1822 21035 -1788 21067
rect -1822 20967 -1788 20995
rect -1822 20899 -1788 20923
rect -1822 20831 -1788 20851
rect -1822 20763 -1788 20779
rect -1822 20695 -1788 20707
rect -1822 20616 -1788 20635
rect -1564 21605 -1530 21624
rect -1564 21533 -1530 21545
rect -1564 21461 -1530 21477
rect -1564 21389 -1530 21409
rect -1564 21317 -1530 21341
rect -1564 21245 -1530 21273
rect -1564 21173 -1530 21205
rect -1564 21103 -1530 21137
rect -1564 21035 -1530 21067
rect -1564 20967 -1530 20995
rect -1564 20899 -1530 20923
rect -1564 20831 -1530 20851
rect -1564 20763 -1530 20779
rect -1564 20695 -1530 20707
rect -1564 20616 -1530 20635
rect -1306 21605 -1272 21624
rect -1306 21533 -1272 21545
rect -1306 21461 -1272 21477
rect -1306 21389 -1272 21409
rect -1306 21317 -1272 21341
rect -1306 21245 -1272 21273
rect -1306 21173 -1272 21205
rect -1306 21103 -1272 21137
rect -1306 21035 -1272 21067
rect -1306 20967 -1272 20995
rect -1306 20899 -1272 20923
rect -1306 20831 -1272 20851
rect -1306 20763 -1272 20779
rect -1306 20695 -1272 20707
rect -1306 20616 -1272 20635
rect -1048 21605 -1014 21624
rect -1048 21533 -1014 21545
rect -1048 21461 -1014 21477
rect -1048 21389 -1014 21409
rect -1048 21317 -1014 21341
rect -1048 21245 -1014 21273
rect -1048 21173 -1014 21205
rect -1048 21103 -1014 21137
rect -1048 21035 -1014 21067
rect -1048 20967 -1014 20995
rect -1048 20899 -1014 20923
rect -1048 20831 -1014 20851
rect -1048 20763 -1014 20779
rect -1048 20695 -1014 20707
rect -1048 20616 -1014 20635
rect -790 21605 -756 21624
rect -790 21533 -756 21545
rect -790 21461 -756 21477
rect -790 21389 -756 21409
rect -790 21317 -756 21341
rect -790 21245 -756 21273
rect -790 21173 -756 21205
rect -790 21103 -756 21137
rect -790 21035 -756 21067
rect -790 20967 -756 20995
rect -790 20899 -756 20923
rect -790 20831 -756 20851
rect -790 20763 -756 20779
rect -790 20695 -756 20707
rect -790 20616 -756 20635
rect -532 21605 -498 21624
rect -532 21533 -498 21545
rect -532 21461 -498 21477
rect -532 21389 -498 21409
rect -532 21317 -498 21341
rect -532 21245 -498 21273
rect -532 21173 -498 21205
rect -532 21103 -498 21137
rect -532 21035 -498 21067
rect -532 20967 -498 20995
rect -532 20899 -498 20923
rect -532 20831 -498 20851
rect -532 20763 -498 20779
rect -532 20695 -498 20707
rect -532 20616 -498 20635
rect -274 21605 -240 21624
rect -274 21533 -240 21545
rect -274 21461 -240 21477
rect -274 21389 -240 21409
rect -274 21317 -240 21341
rect -274 21245 -240 21273
rect -274 21173 -240 21205
rect -274 21103 -240 21137
rect -274 21035 -240 21067
rect -274 20967 -240 20995
rect -274 20899 -240 20923
rect -274 20831 -240 20851
rect -274 20763 -240 20779
rect -274 20695 -240 20707
rect -274 20616 -240 20635
rect -16 21605 18 21624
rect -16 21533 18 21545
rect -16 21461 18 21477
rect -16 21389 18 21409
rect -16 21317 18 21341
rect -16 21245 18 21273
rect -16 21173 18 21205
rect -16 21103 18 21137
rect -16 21035 18 21067
rect -16 20967 18 20995
rect -16 20899 18 20923
rect -16 20831 18 20851
rect -16 20763 18 20779
rect -16 20695 18 20707
rect -16 20616 18 20635
rect 242 21605 276 21624
rect 242 21533 276 21545
rect 242 21461 276 21477
rect 242 21389 276 21409
rect 242 21317 276 21341
rect 242 21245 276 21273
rect 242 21173 276 21205
rect 242 21103 276 21137
rect 242 21035 276 21067
rect 242 20967 276 20995
rect 242 20899 276 20923
rect 242 20831 276 20851
rect 242 20763 276 20779
rect 242 20695 276 20707
rect 242 20616 276 20635
rect 500 21605 534 21624
rect 500 21533 534 21545
rect 500 21461 534 21477
rect 500 21389 534 21409
rect 500 21317 534 21341
rect 500 21245 534 21273
rect 500 21173 534 21205
rect 500 21103 534 21137
rect 500 21035 534 21067
rect 500 20967 534 20995
rect 500 20899 534 20923
rect 500 20831 534 20851
rect 500 20763 534 20779
rect 500 20695 534 20707
rect 500 20616 534 20635
rect 758 21605 792 21624
rect 758 21533 792 21545
rect 758 21461 792 21477
rect 758 21389 792 21409
rect 758 21317 792 21341
rect 758 21245 792 21273
rect 758 21173 792 21205
rect 758 21103 792 21137
rect 758 21035 792 21067
rect 758 20967 792 20995
rect 758 20899 792 20923
rect 758 20831 792 20851
rect 758 20763 792 20779
rect 758 20695 792 20707
rect 758 20616 792 20635
rect 1016 21605 1050 21624
rect 1016 21533 1050 21545
rect 1016 21461 1050 21477
rect 1016 21389 1050 21409
rect 1016 21317 1050 21341
rect 1016 21245 1050 21273
rect 1016 21173 1050 21205
rect 1016 21103 1050 21137
rect 1016 21035 1050 21067
rect 1016 20967 1050 20995
rect 1016 20899 1050 20923
rect 1016 20831 1050 20851
rect 1016 20763 1050 20779
rect 1016 20695 1050 20707
rect 1016 20616 1050 20635
rect 1274 21605 1308 21624
rect 1274 21533 1308 21545
rect 1274 21461 1308 21477
rect 1274 21389 1308 21409
rect 1274 21317 1308 21341
rect 1274 21245 1308 21273
rect 1274 21173 1308 21205
rect 1274 21103 1308 21137
rect 1274 21035 1308 21067
rect 1274 20967 1308 20995
rect 1274 20899 1308 20923
rect 1274 20831 1308 20851
rect 1274 20763 1308 20779
rect 1274 20695 1308 20707
rect 1274 20616 1308 20635
rect 1532 21605 1566 21624
rect 1532 21533 1566 21545
rect 1532 21461 1566 21477
rect 1532 21389 1566 21409
rect 1532 21317 1566 21341
rect 1532 21245 1566 21273
rect 1532 21173 1566 21205
rect 1532 21103 1566 21137
rect 1532 21035 1566 21067
rect 1532 20967 1566 20995
rect 1532 20899 1566 20923
rect 1532 20831 1566 20851
rect 1532 20763 1566 20779
rect 1532 20695 1566 20707
rect 1532 20616 1566 20635
rect 1790 21605 1824 21624
rect 1790 21533 1824 21545
rect 1790 21461 1824 21477
rect 1790 21389 1824 21409
rect 1790 21317 1824 21341
rect 1790 21245 1824 21273
rect 1790 21173 1824 21205
rect 1790 21103 1824 21137
rect 1790 21035 1824 21067
rect 1790 20967 1824 20995
rect 1790 20899 1824 20923
rect 1790 20831 1824 20851
rect 1790 20763 1824 20779
rect 1790 20695 1824 20707
rect 1790 20616 1824 20635
rect 1904 21613 1938 21647
rect 1904 21545 1938 21579
rect 1904 21477 1938 21511
rect 1904 21409 1938 21443
rect 1904 21341 1938 21375
rect 1904 21273 1938 21307
rect 1904 21205 1938 21239
rect 1904 21137 1938 21171
rect 1904 21069 1938 21103
rect 1904 21001 1938 21035
rect 1904 20933 1938 20967
rect 1904 20865 1938 20899
rect 1904 20797 1938 20831
rect 1904 20729 1938 20763
rect 1904 20661 1938 20695
rect 1904 20593 1938 20627
rect -1936 20480 -1902 20559
rect -1776 20548 -1729 20582
rect -1693 20548 -1659 20582
rect -1623 20548 -1576 20582
rect -1518 20548 -1471 20582
rect -1435 20548 -1401 20582
rect -1365 20548 -1318 20582
rect -1260 20548 -1213 20582
rect -1177 20548 -1143 20582
rect -1107 20548 -1060 20582
rect -1002 20548 -955 20582
rect -919 20548 -885 20582
rect -849 20548 -802 20582
rect -744 20548 -697 20582
rect -661 20548 -627 20582
rect -591 20548 -544 20582
rect -486 20548 -439 20582
rect -403 20548 -369 20582
rect -333 20548 -286 20582
rect -228 20548 -181 20582
rect -145 20548 -111 20582
rect -75 20548 -28 20582
rect 30 20548 77 20582
rect 113 20548 147 20582
rect 183 20548 230 20582
rect 288 20548 335 20582
rect 371 20548 405 20582
rect 441 20548 488 20582
rect 546 20548 593 20582
rect 629 20548 663 20582
rect 699 20548 746 20582
rect 804 20548 851 20582
rect 887 20548 921 20582
rect 957 20548 1004 20582
rect 1062 20548 1109 20582
rect 1145 20548 1179 20582
rect 1215 20548 1262 20582
rect 1320 20548 1367 20582
rect 1403 20548 1437 20582
rect 1473 20548 1520 20582
rect 1578 20548 1625 20582
rect 1661 20548 1695 20582
rect 1731 20548 1778 20582
rect 1904 20480 1938 20559
rect -1936 20446 -1818 20480
rect -1784 20446 -1750 20480
rect -1716 20446 -1682 20480
rect -1648 20446 -1614 20480
rect -1580 20446 -1546 20480
rect -1512 20446 -1478 20480
rect -1444 20446 -1410 20480
rect -1376 20446 -1342 20480
rect -1308 20446 -1274 20480
rect -1240 20446 -1206 20480
rect -1172 20446 -1138 20480
rect -1104 20446 -1070 20480
rect -1036 20446 -1002 20480
rect -968 20446 -934 20480
rect -882 20446 -866 20480
rect -810 20446 -798 20480
rect -738 20446 -730 20480
rect -666 20446 -662 20480
rect -560 20446 -556 20480
rect -492 20446 -484 20480
rect -424 20446 -412 20480
rect -356 20446 -340 20480
rect -288 20446 -268 20480
rect -220 20446 -196 20480
rect -152 20446 -124 20480
rect -84 20446 -52 20480
rect -16 20446 18 20480
rect 54 20446 86 20480
rect 126 20446 154 20480
rect 198 20446 222 20480
rect 270 20446 290 20480
rect 342 20446 358 20480
rect 414 20446 426 20480
rect 486 20446 494 20480
rect 558 20446 562 20480
rect 664 20446 668 20480
rect 732 20446 740 20480
rect 800 20446 812 20480
rect 868 20446 884 20480
rect 936 20446 970 20480
rect 1004 20446 1038 20480
rect 1072 20446 1106 20480
rect 1140 20446 1174 20480
rect 1208 20446 1242 20480
rect 1276 20446 1310 20480
rect 1344 20446 1378 20480
rect 1412 20446 1446 20480
rect 1480 20446 1514 20480
rect 1548 20446 1582 20480
rect 1616 20446 1650 20480
rect 1684 20446 1718 20480
rect 1752 20446 1786 20480
rect 1820 20446 1938 20480
rect -3774 19512 -3678 19546
rect 3676 19512 3772 19546
rect -3774 19450 -3740 19512
rect 3738 19450 3772 19512
rect -3595 19398 -3579 19432
rect -2603 19398 -2587 19432
rect -2359 19398 -2343 19432
rect -1367 19398 -1351 19432
rect -1123 19398 -1107 19432
rect -131 19398 -115 19432
rect 113 19398 129 19432
rect 1105 19398 1121 19432
rect 1349 19398 1365 19432
rect 2341 19398 2357 19432
rect 2585 19398 2601 19432
rect 3577 19398 3593 19432
rect -3672 19370 -3638 19386
rect -3672 19186 -3638 19202
rect -2544 19370 -2510 19386
rect -2544 19186 -2510 19202
rect -2436 19370 -2402 19386
rect -2436 19186 -2402 19202
rect -1308 19370 -1274 19386
rect -1308 19186 -1274 19202
rect -1200 19370 -1166 19386
rect -1200 19186 -1166 19202
rect -72 19370 -38 19386
rect -72 19186 -38 19202
rect 36 19370 70 19386
rect 36 19186 70 19202
rect 1164 19370 1198 19386
rect 1164 19186 1198 19202
rect 1272 19370 1306 19386
rect 1272 19186 1306 19202
rect 2400 19370 2434 19386
rect 2400 19186 2434 19202
rect 2508 19370 2542 19386
rect 2508 19186 2542 19202
rect 3636 19370 3670 19386
rect 3636 19186 3670 19202
rect -3595 19140 -3579 19174
rect -2603 19140 -2587 19174
rect -2359 19140 -2343 19174
rect -1367 19140 -1351 19174
rect -1123 19140 -1107 19174
rect -131 19140 -115 19174
rect 113 19140 129 19174
rect 1105 19140 1121 19174
rect 1349 19140 1365 19174
rect 2341 19140 2357 19174
rect 2585 19140 2601 19174
rect 3577 19140 3593 19174
rect -3774 19060 -3740 19122
rect 3738 19060 3772 19122
rect -3774 19026 -3678 19060
rect 3676 19026 3772 19060
rect -3774 18922 -3678 18956
rect 3676 18922 3772 18956
rect -3774 18860 -3740 18922
rect 3738 18860 3772 18922
rect -3595 18808 -3579 18842
rect -2603 18808 -2587 18842
rect -2359 18808 -2343 18842
rect -1367 18808 -1351 18842
rect -1123 18808 -1107 18842
rect -131 18808 -115 18842
rect 113 18808 129 18842
rect 1105 18808 1121 18842
rect 1349 18808 1365 18842
rect 2341 18808 2357 18842
rect 2585 18808 2601 18842
rect 3577 18808 3593 18842
rect -3672 18780 -3638 18796
rect -3672 18596 -3638 18612
rect -2544 18780 -2510 18796
rect -2544 18596 -2510 18612
rect -2436 18780 -2402 18796
rect -2436 18596 -2402 18612
rect -1308 18780 -1274 18796
rect -1308 18596 -1274 18612
rect -1200 18780 -1166 18796
rect -1200 18596 -1166 18612
rect -72 18780 -38 18796
rect -72 18596 -38 18612
rect 36 18780 70 18796
rect 36 18596 70 18612
rect 1164 18780 1198 18796
rect 1164 18596 1198 18612
rect 1272 18780 1306 18796
rect 1272 18596 1306 18612
rect 2400 18780 2434 18796
rect 2400 18596 2434 18612
rect 2508 18780 2542 18796
rect 2508 18596 2542 18612
rect 3636 18780 3670 18796
rect 3636 18596 3670 18612
rect -3595 18550 -3579 18584
rect -2603 18550 -2587 18584
rect -2359 18550 -2343 18584
rect -1367 18550 -1351 18584
rect -1123 18550 -1107 18584
rect -131 18550 -115 18584
rect 113 18550 129 18584
rect 1105 18550 1121 18584
rect 1349 18550 1365 18584
rect 2341 18550 2357 18584
rect 2585 18550 2601 18584
rect 3577 18550 3593 18584
rect -3774 18470 -3740 18532
rect 3738 18470 3772 18532
rect -3774 18436 -3678 18470
rect 3676 18436 3772 18470
rect -1004 18132 -908 18166
rect 902 18132 998 18166
rect -1004 18070 -970 18132
rect 964 18070 998 18132
rect -834 18018 -818 18052
rect -592 18018 -576 18052
rect -366 18018 -350 18052
rect -124 18018 -108 18052
rect 102 18018 118 18052
rect 344 18018 360 18052
rect 570 18018 586 18052
rect 812 18018 828 18052
rect -902 17990 -868 18006
rect -902 17806 -868 17822
rect -542 17990 -508 18006
rect -542 17806 -508 17822
rect -434 17990 -400 18006
rect -434 17806 -400 17822
rect -74 17990 -40 18006
rect -74 17806 -40 17822
rect 34 17990 68 18006
rect 34 17806 68 17822
rect 394 17990 428 18006
rect 394 17806 428 17822
rect 502 17990 536 18006
rect 502 17806 536 17822
rect 862 17990 896 18006
rect 862 17806 896 17822
rect -834 17760 -818 17794
rect -592 17760 -576 17794
rect -366 17760 -350 17794
rect -124 17760 -108 17794
rect 102 17760 118 17794
rect 344 17760 360 17794
rect 570 17760 586 17794
rect 812 17760 828 17794
rect -1004 17680 -970 17742
rect 964 17680 998 17742
rect -1004 17646 -908 17680
rect 902 17646 998 17680
rect -784 17507 -688 17530
rect 686 17507 782 17530
rect -784 17445 -750 17507
rect 748 17445 782 17507
rect -614 17393 -598 17427
rect -122 17393 -106 17427
rect 104 17393 120 17427
rect 596 17393 612 17427
rect -682 17365 -648 17381
rect -682 17281 -648 17297
rect -72 17365 -38 17381
rect -72 17281 -38 17297
rect 36 17365 70 17381
rect 36 17281 70 17297
rect 646 17365 680 17381
rect 646 17281 680 17297
rect -614 17235 -598 17269
rect -122 17235 -106 17269
rect 104 17235 120 17269
rect 596 17235 612 17269
rect -784 17155 -750 17217
rect 748 17155 782 17217
rect -784 17121 -688 17155
rect 686 17121 782 17155
rect -3719 16982 -3623 17016
rect 3623 16982 3719 17016
rect -3719 16920 -3685 16982
rect 3685 16920 3719 16982
rect -3549 16868 -3533 16902
rect -2557 16868 -2541 16902
rect -2331 16868 -2315 16902
rect -1339 16868 -1323 16902
rect -1113 16868 -1097 16902
rect -121 16868 -105 16902
rect 105 16868 121 16902
rect 1097 16868 1113 16902
rect 1323 16868 1339 16902
rect 2315 16868 2331 16902
rect 2541 16868 2557 16902
rect 3533 16868 3549 16902
rect -3617 16840 -3583 16856
rect -3617 16656 -3583 16672
rect -2507 16840 -2473 16856
rect -2507 16656 -2473 16672
rect -2399 16840 -2365 16856
rect -2399 16656 -2365 16672
rect -1289 16840 -1255 16856
rect -1289 16656 -1255 16672
rect -1181 16840 -1147 16856
rect -1181 16656 -1147 16672
rect -71 16840 -37 16856
rect -71 16656 -37 16672
rect 37 16840 71 16856
rect 37 16656 71 16672
rect 1147 16840 1181 16856
rect 1147 16656 1181 16672
rect 1255 16840 1289 16856
rect 1255 16656 1289 16672
rect 2365 16840 2399 16856
rect 2365 16656 2399 16672
rect 2473 16840 2507 16856
rect 2473 16656 2507 16672
rect 3583 16840 3617 16856
rect 3583 16656 3617 16672
rect -3549 16610 -3533 16644
rect -2557 16610 -2541 16644
rect -2331 16610 -2315 16644
rect -1339 16610 -1323 16644
rect -1113 16610 -1097 16644
rect -121 16610 -105 16644
rect 105 16610 121 16644
rect 1097 16610 1113 16644
rect 1323 16610 1339 16644
rect 2315 16610 2331 16644
rect 2541 16610 2557 16644
rect 3533 16610 3549 16644
rect -3719 16530 -3685 16592
rect 3685 16530 3719 16592
rect -3719 16496 -3623 16530
rect 3623 16496 3719 16530
rect -3240 15220 -3120 15236
rect -3240 15084 -3120 15100
rect 3130 15220 3250 15236
rect 3130 15084 3250 15100
rect -3240 12220 -3120 12236
rect -3240 12084 -3120 12100
rect 3130 12220 3250 12236
rect 3130 12084 3250 12100
rect -3240 9220 -3120 9236
rect -3240 9084 -3120 9100
rect 3130 9220 3250 9236
rect 3130 9084 3250 9100
rect -3240 6220 -3120 6236
rect -3240 6084 -3120 6100
rect 3130 6220 3250 6236
rect 3130 6084 3250 6100
rect -3240 3220 -3120 3236
rect -3240 3084 -3120 3100
rect 3130 3220 3250 3236
rect 3130 3084 3250 3100
<< viali >>
rect -7116 30812 -6719 31926
rect -4685 30812 -4288 31926
rect -1596 31108 -1576 31142
rect -1576 31108 -1562 31142
rect -1524 31108 -1508 31142
rect -1508 31108 -1490 31142
rect -1452 31108 -1440 31142
rect -1440 31108 -1418 31142
rect -1380 31108 -1372 31142
rect -1372 31108 -1346 31142
rect -1308 31108 -1304 31142
rect -1304 31108 -1274 31142
rect -1236 31108 -1202 31142
rect -1164 31108 -1134 31142
rect -1134 31108 -1130 31142
rect -1092 31108 -1066 31142
rect -1066 31108 -1058 31142
rect -1020 31108 -998 31142
rect -998 31108 -986 31142
rect -948 31108 -930 31142
rect -930 31108 -914 31142
rect -876 31108 -862 31142
rect -862 31108 -842 31142
rect -804 31108 -794 31142
rect -794 31108 -770 31142
rect -732 31108 -726 31142
rect -726 31108 -698 31142
rect -660 31108 -658 31142
rect -658 31108 -626 31142
rect -588 31108 -556 31142
rect -556 31108 -554 31142
rect -516 31108 -488 31142
rect -488 31108 -482 31142
rect -444 31108 -420 31142
rect -420 31108 -410 31142
rect -372 31108 -352 31142
rect -352 31108 -338 31142
rect -300 31108 -284 31142
rect -284 31108 -266 31142
rect -228 31108 -216 31142
rect -216 31108 -194 31142
rect -156 31108 -148 31142
rect -148 31108 -122 31142
rect -84 31108 -80 31142
rect -80 31108 -50 31142
rect -12 31108 22 31142
rect 60 31108 90 31142
rect 90 31108 94 31142
rect 132 31108 158 31142
rect 158 31108 166 31142
rect 204 31108 226 31142
rect 226 31108 238 31142
rect 276 31108 294 31142
rect 294 31108 310 31142
rect 348 31108 362 31142
rect 362 31108 382 31142
rect 420 31108 430 31142
rect 430 31108 454 31142
rect 492 31108 498 31142
rect 498 31108 526 31142
rect 564 31108 566 31142
rect 566 31108 598 31142
rect 636 31108 668 31142
rect 668 31108 670 31142
rect 708 31108 736 31142
rect 736 31108 742 31142
rect 780 31108 804 31142
rect 804 31108 814 31142
rect 852 31108 872 31142
rect 872 31108 886 31142
rect 924 31108 940 31142
rect 940 31108 958 31142
rect 996 31108 1008 31142
rect 1008 31108 1030 31142
rect 1068 31108 1076 31142
rect 1076 31108 1102 31142
rect 1140 31108 1144 31142
rect 1144 31108 1174 31142
rect 1212 31108 1246 31142
rect 1284 31108 1314 31142
rect 1314 31108 1318 31142
rect 1356 31108 1382 31142
rect 1382 31108 1390 31142
rect 1428 31108 1450 31142
rect 1450 31108 1462 31142
rect 1500 31108 1518 31142
rect 1518 31108 1534 31142
rect 1572 31108 1586 31142
rect 1586 31108 1606 31142
rect -3093 31006 -3059 31040
rect -2935 31006 -2901 31040
rect -2777 31006 -2743 31040
rect -2619 31006 -2585 31040
rect -2461 31006 -2427 31040
rect -2303 31006 -2269 31040
rect -2145 31006 -2111 31040
rect -1987 31006 -1953 31040
rect -1829 31006 -1795 31040
rect -1671 31006 -1637 31040
rect -1513 31006 -1479 31040
rect -1355 31006 -1321 31040
rect -1197 31006 -1163 31040
rect -1039 31006 -1005 31040
rect -881 31006 -847 31040
rect -723 31006 -689 31040
rect -565 31006 -531 31040
rect -407 31006 -373 31040
rect -249 31006 -215 31040
rect -91 31006 -57 31040
rect 67 31006 101 31040
rect 225 31006 259 31040
rect 383 31006 417 31040
rect 541 31006 575 31040
rect 699 31006 733 31040
rect 857 31006 891 31040
rect 1015 31006 1049 31040
rect 1173 31006 1207 31040
rect 1331 31006 1365 31040
rect 1489 31006 1523 31040
rect 1647 31006 1681 31040
rect 1805 31006 1839 31040
rect 1963 31006 1997 31040
rect 2121 31006 2155 31040
rect 2279 31006 2313 31040
rect 2437 31006 2471 31040
rect 2595 31006 2629 31040
rect 2753 31006 2787 31040
rect 2911 31006 2945 31040
rect 3069 31006 3103 31040
rect -7116 29312 -6719 30426
rect -4685 29312 -4288 30426
rect -3172 30918 -3138 30944
rect -3172 30910 -3138 30918
rect -3172 30850 -3138 30872
rect -3172 30838 -3138 30850
rect -3172 30782 -3138 30800
rect -3172 30766 -3138 30782
rect -3172 30714 -3138 30728
rect -3172 30694 -3138 30714
rect -3172 30646 -3138 30656
rect -3172 30622 -3138 30646
rect -3172 30578 -3138 30584
rect -3172 30550 -3138 30578
rect -3172 30510 -3138 30512
rect -3172 30478 -3138 30510
rect -3172 30408 -3138 30440
rect -3172 30406 -3138 30408
rect -3172 30340 -3138 30368
rect -3172 30334 -3138 30340
rect -3172 30272 -3138 30296
rect -3172 30262 -3138 30272
rect -3172 30204 -3138 30224
rect -3172 30190 -3138 30204
rect -3172 30136 -3138 30152
rect -3172 30118 -3138 30136
rect -3172 30068 -3138 30080
rect -3172 30046 -3138 30068
rect -3172 30000 -3138 30008
rect -3172 29974 -3138 30000
rect -3014 30918 -2980 30944
rect -3014 30910 -2980 30918
rect -3014 30850 -2980 30872
rect -3014 30838 -2980 30850
rect -3014 30782 -2980 30800
rect -3014 30766 -2980 30782
rect -3014 30714 -2980 30728
rect -3014 30694 -2980 30714
rect -3014 30646 -2980 30656
rect -3014 30622 -2980 30646
rect -3014 30578 -2980 30584
rect -3014 30550 -2980 30578
rect -3014 30510 -2980 30512
rect -3014 30478 -2980 30510
rect -3014 30408 -2980 30440
rect -3014 30406 -2980 30408
rect -3014 30340 -2980 30368
rect -3014 30334 -2980 30340
rect -3014 30272 -2980 30296
rect -3014 30262 -2980 30272
rect -3014 30204 -2980 30224
rect -3014 30190 -2980 30204
rect -3014 30136 -2980 30152
rect -3014 30118 -2980 30136
rect -3014 30068 -2980 30080
rect -3014 30046 -2980 30068
rect -3014 30000 -2980 30008
rect -3014 29974 -2980 30000
rect -2856 30918 -2822 30944
rect -2856 30910 -2822 30918
rect -2856 30850 -2822 30872
rect -2856 30838 -2822 30850
rect -2856 30782 -2822 30800
rect -2856 30766 -2822 30782
rect -2856 30714 -2822 30728
rect -2856 30694 -2822 30714
rect -2856 30646 -2822 30656
rect -2856 30622 -2822 30646
rect -2856 30578 -2822 30584
rect -2856 30550 -2822 30578
rect -2856 30510 -2822 30512
rect -2856 30478 -2822 30510
rect -2856 30408 -2822 30440
rect -2856 30406 -2822 30408
rect -2856 30340 -2822 30368
rect -2856 30334 -2822 30340
rect -2856 30272 -2822 30296
rect -2856 30262 -2822 30272
rect -2856 30204 -2822 30224
rect -2856 30190 -2822 30204
rect -2856 30136 -2822 30152
rect -2856 30118 -2822 30136
rect -2856 30068 -2822 30080
rect -2856 30046 -2822 30068
rect -2856 30000 -2822 30008
rect -2856 29974 -2822 30000
rect -2698 30918 -2664 30944
rect -2698 30910 -2664 30918
rect -2698 30850 -2664 30872
rect -2698 30838 -2664 30850
rect -2698 30782 -2664 30800
rect -2698 30766 -2664 30782
rect -2698 30714 -2664 30728
rect -2698 30694 -2664 30714
rect -2698 30646 -2664 30656
rect -2698 30622 -2664 30646
rect -2698 30578 -2664 30584
rect -2698 30550 -2664 30578
rect -2698 30510 -2664 30512
rect -2698 30478 -2664 30510
rect -2698 30408 -2664 30440
rect -2698 30406 -2664 30408
rect -2698 30340 -2664 30368
rect -2698 30334 -2664 30340
rect -2698 30272 -2664 30296
rect -2698 30262 -2664 30272
rect -2698 30204 -2664 30224
rect -2698 30190 -2664 30204
rect -2698 30136 -2664 30152
rect -2698 30118 -2664 30136
rect -2698 30068 -2664 30080
rect -2698 30046 -2664 30068
rect -2698 30000 -2664 30008
rect -2698 29974 -2664 30000
rect -2540 30918 -2506 30944
rect -2540 30910 -2506 30918
rect -2540 30850 -2506 30872
rect -2540 30838 -2506 30850
rect -2540 30782 -2506 30800
rect -2540 30766 -2506 30782
rect -2540 30714 -2506 30728
rect -2540 30694 -2506 30714
rect -2540 30646 -2506 30656
rect -2540 30622 -2506 30646
rect -2540 30578 -2506 30584
rect -2540 30550 -2506 30578
rect -2540 30510 -2506 30512
rect -2540 30478 -2506 30510
rect -2540 30408 -2506 30440
rect -2540 30406 -2506 30408
rect -2540 30340 -2506 30368
rect -2540 30334 -2506 30340
rect -2540 30272 -2506 30296
rect -2540 30262 -2506 30272
rect -2540 30204 -2506 30224
rect -2540 30190 -2506 30204
rect -2540 30136 -2506 30152
rect -2540 30118 -2506 30136
rect -2540 30068 -2506 30080
rect -2540 30046 -2506 30068
rect -2540 30000 -2506 30008
rect -2540 29974 -2506 30000
rect -2382 30918 -2348 30944
rect -2382 30910 -2348 30918
rect -2382 30850 -2348 30872
rect -2382 30838 -2348 30850
rect -2382 30782 -2348 30800
rect -2382 30766 -2348 30782
rect -2382 30714 -2348 30728
rect -2382 30694 -2348 30714
rect -2382 30646 -2348 30656
rect -2382 30622 -2348 30646
rect -2382 30578 -2348 30584
rect -2382 30550 -2348 30578
rect -2382 30510 -2348 30512
rect -2382 30478 -2348 30510
rect -2382 30408 -2348 30440
rect -2382 30406 -2348 30408
rect -2382 30340 -2348 30368
rect -2382 30334 -2348 30340
rect -2382 30272 -2348 30296
rect -2382 30262 -2348 30272
rect -2382 30204 -2348 30224
rect -2382 30190 -2348 30204
rect -2382 30136 -2348 30152
rect -2382 30118 -2348 30136
rect -2382 30068 -2348 30080
rect -2382 30046 -2348 30068
rect -2382 30000 -2348 30008
rect -2382 29974 -2348 30000
rect -2224 30918 -2190 30944
rect -2224 30910 -2190 30918
rect -2224 30850 -2190 30872
rect -2224 30838 -2190 30850
rect -2224 30782 -2190 30800
rect -2224 30766 -2190 30782
rect -2224 30714 -2190 30728
rect -2224 30694 -2190 30714
rect -2224 30646 -2190 30656
rect -2224 30622 -2190 30646
rect -2224 30578 -2190 30584
rect -2224 30550 -2190 30578
rect -2224 30510 -2190 30512
rect -2224 30478 -2190 30510
rect -2224 30408 -2190 30440
rect -2224 30406 -2190 30408
rect -2224 30340 -2190 30368
rect -2224 30334 -2190 30340
rect -2224 30272 -2190 30296
rect -2224 30262 -2190 30272
rect -2224 30204 -2190 30224
rect -2224 30190 -2190 30204
rect -2224 30136 -2190 30152
rect -2224 30118 -2190 30136
rect -2224 30068 -2190 30080
rect -2224 30046 -2190 30068
rect -2224 30000 -2190 30008
rect -2224 29974 -2190 30000
rect -2066 30918 -2032 30944
rect -2066 30910 -2032 30918
rect -2066 30850 -2032 30872
rect -2066 30838 -2032 30850
rect -2066 30782 -2032 30800
rect -2066 30766 -2032 30782
rect -2066 30714 -2032 30728
rect -2066 30694 -2032 30714
rect -2066 30646 -2032 30656
rect -2066 30622 -2032 30646
rect -2066 30578 -2032 30584
rect -2066 30550 -2032 30578
rect -2066 30510 -2032 30512
rect -2066 30478 -2032 30510
rect -2066 30408 -2032 30440
rect -2066 30406 -2032 30408
rect -2066 30340 -2032 30368
rect -2066 30334 -2032 30340
rect -2066 30272 -2032 30296
rect -2066 30262 -2032 30272
rect -2066 30204 -2032 30224
rect -2066 30190 -2032 30204
rect -2066 30136 -2032 30152
rect -2066 30118 -2032 30136
rect -2066 30068 -2032 30080
rect -2066 30046 -2032 30068
rect -2066 30000 -2032 30008
rect -2066 29974 -2032 30000
rect -1908 30918 -1874 30944
rect -1908 30910 -1874 30918
rect -1908 30850 -1874 30872
rect -1908 30838 -1874 30850
rect -1908 30782 -1874 30800
rect -1908 30766 -1874 30782
rect -1908 30714 -1874 30728
rect -1908 30694 -1874 30714
rect -1908 30646 -1874 30656
rect -1908 30622 -1874 30646
rect -1908 30578 -1874 30584
rect -1908 30550 -1874 30578
rect -1908 30510 -1874 30512
rect -1908 30478 -1874 30510
rect -1908 30408 -1874 30440
rect -1908 30406 -1874 30408
rect -1908 30340 -1874 30368
rect -1908 30334 -1874 30340
rect -1908 30272 -1874 30296
rect -1908 30262 -1874 30272
rect -1908 30204 -1874 30224
rect -1908 30190 -1874 30204
rect -1908 30136 -1874 30152
rect -1908 30118 -1874 30136
rect -1908 30068 -1874 30080
rect -1908 30046 -1874 30068
rect -1908 30000 -1874 30008
rect -1908 29974 -1874 30000
rect -1750 30918 -1716 30944
rect -1750 30910 -1716 30918
rect -1750 30850 -1716 30872
rect -1750 30838 -1716 30850
rect -1750 30782 -1716 30800
rect -1750 30766 -1716 30782
rect -1750 30714 -1716 30728
rect -1750 30694 -1716 30714
rect -1750 30646 -1716 30656
rect -1750 30622 -1716 30646
rect -1750 30578 -1716 30584
rect -1750 30550 -1716 30578
rect -1750 30510 -1716 30512
rect -1750 30478 -1716 30510
rect -1750 30408 -1716 30440
rect -1750 30406 -1716 30408
rect -1750 30340 -1716 30368
rect -1750 30334 -1716 30340
rect -1750 30272 -1716 30296
rect -1750 30262 -1716 30272
rect -1750 30204 -1716 30224
rect -1750 30190 -1716 30204
rect -1750 30136 -1716 30152
rect -1750 30118 -1716 30136
rect -1750 30068 -1716 30080
rect -1750 30046 -1716 30068
rect -1750 30000 -1716 30008
rect -1750 29974 -1716 30000
rect -1592 30918 -1558 30944
rect -1592 30910 -1558 30918
rect -1592 30850 -1558 30872
rect -1592 30838 -1558 30850
rect -1592 30782 -1558 30800
rect -1592 30766 -1558 30782
rect -1592 30714 -1558 30728
rect -1592 30694 -1558 30714
rect -1592 30646 -1558 30656
rect -1592 30622 -1558 30646
rect -1592 30578 -1558 30584
rect -1592 30550 -1558 30578
rect -1592 30510 -1558 30512
rect -1592 30478 -1558 30510
rect -1592 30408 -1558 30440
rect -1592 30406 -1558 30408
rect -1592 30340 -1558 30368
rect -1592 30334 -1558 30340
rect -1592 30272 -1558 30296
rect -1592 30262 -1558 30272
rect -1592 30204 -1558 30224
rect -1592 30190 -1558 30204
rect -1592 30136 -1558 30152
rect -1592 30118 -1558 30136
rect -1592 30068 -1558 30080
rect -1592 30046 -1558 30068
rect -1592 30000 -1558 30008
rect -1592 29974 -1558 30000
rect -1434 30918 -1400 30944
rect -1434 30910 -1400 30918
rect -1434 30850 -1400 30872
rect -1434 30838 -1400 30850
rect -1434 30782 -1400 30800
rect -1434 30766 -1400 30782
rect -1434 30714 -1400 30728
rect -1434 30694 -1400 30714
rect -1434 30646 -1400 30656
rect -1434 30622 -1400 30646
rect -1434 30578 -1400 30584
rect -1434 30550 -1400 30578
rect -1434 30510 -1400 30512
rect -1434 30478 -1400 30510
rect -1434 30408 -1400 30440
rect -1434 30406 -1400 30408
rect -1434 30340 -1400 30368
rect -1434 30334 -1400 30340
rect -1434 30272 -1400 30296
rect -1434 30262 -1400 30272
rect -1434 30204 -1400 30224
rect -1434 30190 -1400 30204
rect -1434 30136 -1400 30152
rect -1434 30118 -1400 30136
rect -1434 30068 -1400 30080
rect -1434 30046 -1400 30068
rect -1434 30000 -1400 30008
rect -1434 29974 -1400 30000
rect -1276 30918 -1242 30944
rect -1276 30910 -1242 30918
rect -1276 30850 -1242 30872
rect -1276 30838 -1242 30850
rect -1276 30782 -1242 30800
rect -1276 30766 -1242 30782
rect -1276 30714 -1242 30728
rect -1276 30694 -1242 30714
rect -1276 30646 -1242 30656
rect -1276 30622 -1242 30646
rect -1276 30578 -1242 30584
rect -1276 30550 -1242 30578
rect -1276 30510 -1242 30512
rect -1276 30478 -1242 30510
rect -1276 30408 -1242 30440
rect -1276 30406 -1242 30408
rect -1276 30340 -1242 30368
rect -1276 30334 -1242 30340
rect -1276 30272 -1242 30296
rect -1276 30262 -1242 30272
rect -1276 30204 -1242 30224
rect -1276 30190 -1242 30204
rect -1276 30136 -1242 30152
rect -1276 30118 -1242 30136
rect -1276 30068 -1242 30080
rect -1276 30046 -1242 30068
rect -1276 30000 -1242 30008
rect -1276 29974 -1242 30000
rect -1118 30918 -1084 30944
rect -1118 30910 -1084 30918
rect -1118 30850 -1084 30872
rect -1118 30838 -1084 30850
rect -1118 30782 -1084 30800
rect -1118 30766 -1084 30782
rect -1118 30714 -1084 30728
rect -1118 30694 -1084 30714
rect -1118 30646 -1084 30656
rect -1118 30622 -1084 30646
rect -1118 30578 -1084 30584
rect -1118 30550 -1084 30578
rect -1118 30510 -1084 30512
rect -1118 30478 -1084 30510
rect -1118 30408 -1084 30440
rect -1118 30406 -1084 30408
rect -1118 30340 -1084 30368
rect -1118 30334 -1084 30340
rect -1118 30272 -1084 30296
rect -1118 30262 -1084 30272
rect -1118 30204 -1084 30224
rect -1118 30190 -1084 30204
rect -1118 30136 -1084 30152
rect -1118 30118 -1084 30136
rect -1118 30068 -1084 30080
rect -1118 30046 -1084 30068
rect -1118 30000 -1084 30008
rect -1118 29974 -1084 30000
rect -960 30918 -926 30944
rect -960 30910 -926 30918
rect -960 30850 -926 30872
rect -960 30838 -926 30850
rect -960 30782 -926 30800
rect -960 30766 -926 30782
rect -960 30714 -926 30728
rect -960 30694 -926 30714
rect -960 30646 -926 30656
rect -960 30622 -926 30646
rect -960 30578 -926 30584
rect -960 30550 -926 30578
rect -960 30510 -926 30512
rect -960 30478 -926 30510
rect -960 30408 -926 30440
rect -960 30406 -926 30408
rect -960 30340 -926 30368
rect -960 30334 -926 30340
rect -960 30272 -926 30296
rect -960 30262 -926 30272
rect -960 30204 -926 30224
rect -960 30190 -926 30204
rect -960 30136 -926 30152
rect -960 30118 -926 30136
rect -960 30068 -926 30080
rect -960 30046 -926 30068
rect -960 30000 -926 30008
rect -960 29974 -926 30000
rect -802 30918 -768 30944
rect -802 30910 -768 30918
rect -802 30850 -768 30872
rect -802 30838 -768 30850
rect -802 30782 -768 30800
rect -802 30766 -768 30782
rect -802 30714 -768 30728
rect -802 30694 -768 30714
rect -802 30646 -768 30656
rect -802 30622 -768 30646
rect -802 30578 -768 30584
rect -802 30550 -768 30578
rect -802 30510 -768 30512
rect -802 30478 -768 30510
rect -802 30408 -768 30440
rect -802 30406 -768 30408
rect -802 30340 -768 30368
rect -802 30334 -768 30340
rect -802 30272 -768 30296
rect -802 30262 -768 30272
rect -802 30204 -768 30224
rect -802 30190 -768 30204
rect -802 30136 -768 30152
rect -802 30118 -768 30136
rect -802 30068 -768 30080
rect -802 30046 -768 30068
rect -802 30000 -768 30008
rect -802 29974 -768 30000
rect -644 30918 -610 30944
rect -644 30910 -610 30918
rect -644 30850 -610 30872
rect -644 30838 -610 30850
rect -644 30782 -610 30800
rect -644 30766 -610 30782
rect -644 30714 -610 30728
rect -644 30694 -610 30714
rect -644 30646 -610 30656
rect -644 30622 -610 30646
rect -644 30578 -610 30584
rect -644 30550 -610 30578
rect -644 30510 -610 30512
rect -644 30478 -610 30510
rect -644 30408 -610 30440
rect -644 30406 -610 30408
rect -644 30340 -610 30368
rect -644 30334 -610 30340
rect -644 30272 -610 30296
rect -644 30262 -610 30272
rect -644 30204 -610 30224
rect -644 30190 -610 30204
rect -644 30136 -610 30152
rect -644 30118 -610 30136
rect -644 30068 -610 30080
rect -644 30046 -610 30068
rect -644 30000 -610 30008
rect -644 29974 -610 30000
rect -486 30918 -452 30944
rect -486 30910 -452 30918
rect -486 30850 -452 30872
rect -486 30838 -452 30850
rect -486 30782 -452 30800
rect -486 30766 -452 30782
rect -486 30714 -452 30728
rect -486 30694 -452 30714
rect -486 30646 -452 30656
rect -486 30622 -452 30646
rect -486 30578 -452 30584
rect -486 30550 -452 30578
rect -486 30510 -452 30512
rect -486 30478 -452 30510
rect -486 30408 -452 30440
rect -486 30406 -452 30408
rect -486 30340 -452 30368
rect -486 30334 -452 30340
rect -486 30272 -452 30296
rect -486 30262 -452 30272
rect -486 30204 -452 30224
rect -486 30190 -452 30204
rect -486 30136 -452 30152
rect -486 30118 -452 30136
rect -486 30068 -452 30080
rect -486 30046 -452 30068
rect -486 30000 -452 30008
rect -486 29974 -452 30000
rect -328 30918 -294 30944
rect -328 30910 -294 30918
rect -328 30850 -294 30872
rect -328 30838 -294 30850
rect -328 30782 -294 30800
rect -328 30766 -294 30782
rect -328 30714 -294 30728
rect -328 30694 -294 30714
rect -328 30646 -294 30656
rect -328 30622 -294 30646
rect -328 30578 -294 30584
rect -328 30550 -294 30578
rect -328 30510 -294 30512
rect -328 30478 -294 30510
rect -328 30408 -294 30440
rect -328 30406 -294 30408
rect -328 30340 -294 30368
rect -328 30334 -294 30340
rect -328 30272 -294 30296
rect -328 30262 -294 30272
rect -328 30204 -294 30224
rect -328 30190 -294 30204
rect -328 30136 -294 30152
rect -328 30118 -294 30136
rect -328 30068 -294 30080
rect -328 30046 -294 30068
rect -328 30000 -294 30008
rect -328 29974 -294 30000
rect -170 30918 -136 30944
rect -170 30910 -136 30918
rect -170 30850 -136 30872
rect -170 30838 -136 30850
rect -170 30782 -136 30800
rect -170 30766 -136 30782
rect -170 30714 -136 30728
rect -170 30694 -136 30714
rect -170 30646 -136 30656
rect -170 30622 -136 30646
rect -170 30578 -136 30584
rect -170 30550 -136 30578
rect -170 30510 -136 30512
rect -170 30478 -136 30510
rect -170 30408 -136 30440
rect -170 30406 -136 30408
rect -170 30340 -136 30368
rect -170 30334 -136 30340
rect -170 30272 -136 30296
rect -170 30262 -136 30272
rect -170 30204 -136 30224
rect -170 30190 -136 30204
rect -170 30136 -136 30152
rect -170 30118 -136 30136
rect -170 30068 -136 30080
rect -170 30046 -136 30068
rect -170 30000 -136 30008
rect -170 29974 -136 30000
rect -12 30918 22 30944
rect -12 30910 22 30918
rect -12 30850 22 30872
rect -12 30838 22 30850
rect -12 30782 22 30800
rect -12 30766 22 30782
rect -12 30714 22 30728
rect -12 30694 22 30714
rect -12 30646 22 30656
rect -12 30622 22 30646
rect -12 30578 22 30584
rect -12 30550 22 30578
rect -12 30510 22 30512
rect -12 30478 22 30510
rect -12 30408 22 30440
rect -12 30406 22 30408
rect -12 30340 22 30368
rect -12 30334 22 30340
rect -12 30272 22 30296
rect -12 30262 22 30272
rect -12 30204 22 30224
rect -12 30190 22 30204
rect -12 30136 22 30152
rect -12 30118 22 30136
rect -12 30068 22 30080
rect -12 30046 22 30068
rect -12 30000 22 30008
rect -12 29974 22 30000
rect 146 30918 180 30944
rect 146 30910 180 30918
rect 146 30850 180 30872
rect 146 30838 180 30850
rect 146 30782 180 30800
rect 146 30766 180 30782
rect 146 30714 180 30728
rect 146 30694 180 30714
rect 146 30646 180 30656
rect 146 30622 180 30646
rect 146 30578 180 30584
rect 146 30550 180 30578
rect 146 30510 180 30512
rect 146 30478 180 30510
rect 146 30408 180 30440
rect 146 30406 180 30408
rect 146 30340 180 30368
rect 146 30334 180 30340
rect 146 30272 180 30296
rect 146 30262 180 30272
rect 146 30204 180 30224
rect 146 30190 180 30204
rect 146 30136 180 30152
rect 146 30118 180 30136
rect 146 30068 180 30080
rect 146 30046 180 30068
rect 146 30000 180 30008
rect 146 29974 180 30000
rect 304 30918 338 30944
rect 304 30910 338 30918
rect 304 30850 338 30872
rect 304 30838 338 30850
rect 304 30782 338 30800
rect 304 30766 338 30782
rect 304 30714 338 30728
rect 304 30694 338 30714
rect 304 30646 338 30656
rect 304 30622 338 30646
rect 304 30578 338 30584
rect 304 30550 338 30578
rect 304 30510 338 30512
rect 304 30478 338 30510
rect 304 30408 338 30440
rect 304 30406 338 30408
rect 304 30340 338 30368
rect 304 30334 338 30340
rect 304 30272 338 30296
rect 304 30262 338 30272
rect 304 30204 338 30224
rect 304 30190 338 30204
rect 304 30136 338 30152
rect 304 30118 338 30136
rect 304 30068 338 30080
rect 304 30046 338 30068
rect 304 30000 338 30008
rect 304 29974 338 30000
rect 462 30918 496 30944
rect 462 30910 496 30918
rect 462 30850 496 30872
rect 462 30838 496 30850
rect 462 30782 496 30800
rect 462 30766 496 30782
rect 462 30714 496 30728
rect 462 30694 496 30714
rect 462 30646 496 30656
rect 462 30622 496 30646
rect 462 30578 496 30584
rect 462 30550 496 30578
rect 462 30510 496 30512
rect 462 30478 496 30510
rect 462 30408 496 30440
rect 462 30406 496 30408
rect 462 30340 496 30368
rect 462 30334 496 30340
rect 462 30272 496 30296
rect 462 30262 496 30272
rect 462 30204 496 30224
rect 462 30190 496 30204
rect 462 30136 496 30152
rect 462 30118 496 30136
rect 462 30068 496 30080
rect 462 30046 496 30068
rect 462 30000 496 30008
rect 462 29974 496 30000
rect 620 30918 654 30944
rect 620 30910 654 30918
rect 620 30850 654 30872
rect 620 30838 654 30850
rect 620 30782 654 30800
rect 620 30766 654 30782
rect 620 30714 654 30728
rect 620 30694 654 30714
rect 620 30646 654 30656
rect 620 30622 654 30646
rect 620 30578 654 30584
rect 620 30550 654 30578
rect 620 30510 654 30512
rect 620 30478 654 30510
rect 620 30408 654 30440
rect 620 30406 654 30408
rect 620 30340 654 30368
rect 620 30334 654 30340
rect 620 30272 654 30296
rect 620 30262 654 30272
rect 620 30204 654 30224
rect 620 30190 654 30204
rect 620 30136 654 30152
rect 620 30118 654 30136
rect 620 30068 654 30080
rect 620 30046 654 30068
rect 620 30000 654 30008
rect 620 29974 654 30000
rect 778 30918 812 30944
rect 778 30910 812 30918
rect 778 30850 812 30872
rect 778 30838 812 30850
rect 778 30782 812 30800
rect 778 30766 812 30782
rect 778 30714 812 30728
rect 778 30694 812 30714
rect 778 30646 812 30656
rect 778 30622 812 30646
rect 778 30578 812 30584
rect 778 30550 812 30578
rect 778 30510 812 30512
rect 778 30478 812 30510
rect 778 30408 812 30440
rect 778 30406 812 30408
rect 778 30340 812 30368
rect 778 30334 812 30340
rect 778 30272 812 30296
rect 778 30262 812 30272
rect 778 30204 812 30224
rect 778 30190 812 30204
rect 778 30136 812 30152
rect 778 30118 812 30136
rect 778 30068 812 30080
rect 778 30046 812 30068
rect 778 30000 812 30008
rect 778 29974 812 30000
rect 936 30918 970 30944
rect 936 30910 970 30918
rect 936 30850 970 30872
rect 936 30838 970 30850
rect 936 30782 970 30800
rect 936 30766 970 30782
rect 936 30714 970 30728
rect 936 30694 970 30714
rect 936 30646 970 30656
rect 936 30622 970 30646
rect 936 30578 970 30584
rect 936 30550 970 30578
rect 936 30510 970 30512
rect 936 30478 970 30510
rect 936 30408 970 30440
rect 936 30406 970 30408
rect 936 30340 970 30368
rect 936 30334 970 30340
rect 936 30272 970 30296
rect 936 30262 970 30272
rect 936 30204 970 30224
rect 936 30190 970 30204
rect 936 30136 970 30152
rect 936 30118 970 30136
rect 936 30068 970 30080
rect 936 30046 970 30068
rect 936 30000 970 30008
rect 936 29974 970 30000
rect 1094 30918 1128 30944
rect 1094 30910 1128 30918
rect 1094 30850 1128 30872
rect 1094 30838 1128 30850
rect 1094 30782 1128 30800
rect 1094 30766 1128 30782
rect 1094 30714 1128 30728
rect 1094 30694 1128 30714
rect 1094 30646 1128 30656
rect 1094 30622 1128 30646
rect 1094 30578 1128 30584
rect 1094 30550 1128 30578
rect 1094 30510 1128 30512
rect 1094 30478 1128 30510
rect 1094 30408 1128 30440
rect 1094 30406 1128 30408
rect 1094 30340 1128 30368
rect 1094 30334 1128 30340
rect 1094 30272 1128 30296
rect 1094 30262 1128 30272
rect 1094 30204 1128 30224
rect 1094 30190 1128 30204
rect 1094 30136 1128 30152
rect 1094 30118 1128 30136
rect 1094 30068 1128 30080
rect 1094 30046 1128 30068
rect 1094 30000 1128 30008
rect 1094 29974 1128 30000
rect 1252 30918 1286 30944
rect 1252 30910 1286 30918
rect 1252 30850 1286 30872
rect 1252 30838 1286 30850
rect 1252 30782 1286 30800
rect 1252 30766 1286 30782
rect 1252 30714 1286 30728
rect 1252 30694 1286 30714
rect 1252 30646 1286 30656
rect 1252 30622 1286 30646
rect 1252 30578 1286 30584
rect 1252 30550 1286 30578
rect 1252 30510 1286 30512
rect 1252 30478 1286 30510
rect 1252 30408 1286 30440
rect 1252 30406 1286 30408
rect 1252 30340 1286 30368
rect 1252 30334 1286 30340
rect 1252 30272 1286 30296
rect 1252 30262 1286 30272
rect 1252 30204 1286 30224
rect 1252 30190 1286 30204
rect 1252 30136 1286 30152
rect 1252 30118 1286 30136
rect 1252 30068 1286 30080
rect 1252 30046 1286 30068
rect 1252 30000 1286 30008
rect 1252 29974 1286 30000
rect 1410 30918 1444 30944
rect 1410 30910 1444 30918
rect 1410 30850 1444 30872
rect 1410 30838 1444 30850
rect 1410 30782 1444 30800
rect 1410 30766 1444 30782
rect 1410 30714 1444 30728
rect 1410 30694 1444 30714
rect 1410 30646 1444 30656
rect 1410 30622 1444 30646
rect 1410 30578 1444 30584
rect 1410 30550 1444 30578
rect 1410 30510 1444 30512
rect 1410 30478 1444 30510
rect 1410 30408 1444 30440
rect 1410 30406 1444 30408
rect 1410 30340 1444 30368
rect 1410 30334 1444 30340
rect 1410 30272 1444 30296
rect 1410 30262 1444 30272
rect 1410 30204 1444 30224
rect 1410 30190 1444 30204
rect 1410 30136 1444 30152
rect 1410 30118 1444 30136
rect 1410 30068 1444 30080
rect 1410 30046 1444 30068
rect 1410 30000 1444 30008
rect 1410 29974 1444 30000
rect 1568 30918 1602 30944
rect 1568 30910 1602 30918
rect 1568 30850 1602 30872
rect 1568 30838 1602 30850
rect 1568 30782 1602 30800
rect 1568 30766 1602 30782
rect 1568 30714 1602 30728
rect 1568 30694 1602 30714
rect 1568 30646 1602 30656
rect 1568 30622 1602 30646
rect 1568 30578 1602 30584
rect 1568 30550 1602 30578
rect 1568 30510 1602 30512
rect 1568 30478 1602 30510
rect 1568 30408 1602 30440
rect 1568 30406 1602 30408
rect 1568 30340 1602 30368
rect 1568 30334 1602 30340
rect 1568 30272 1602 30296
rect 1568 30262 1602 30272
rect 1568 30204 1602 30224
rect 1568 30190 1602 30204
rect 1568 30136 1602 30152
rect 1568 30118 1602 30136
rect 1568 30068 1602 30080
rect 1568 30046 1602 30068
rect 1568 30000 1602 30008
rect 1568 29974 1602 30000
rect 1726 30918 1760 30944
rect 1726 30910 1760 30918
rect 1726 30850 1760 30872
rect 1726 30838 1760 30850
rect 1726 30782 1760 30800
rect 1726 30766 1760 30782
rect 1726 30714 1760 30728
rect 1726 30694 1760 30714
rect 1726 30646 1760 30656
rect 1726 30622 1760 30646
rect 1726 30578 1760 30584
rect 1726 30550 1760 30578
rect 1726 30510 1760 30512
rect 1726 30478 1760 30510
rect 1726 30408 1760 30440
rect 1726 30406 1760 30408
rect 1726 30340 1760 30368
rect 1726 30334 1760 30340
rect 1726 30272 1760 30296
rect 1726 30262 1760 30272
rect 1726 30204 1760 30224
rect 1726 30190 1760 30204
rect 1726 30136 1760 30152
rect 1726 30118 1760 30136
rect 1726 30068 1760 30080
rect 1726 30046 1760 30068
rect 1726 30000 1760 30008
rect 1726 29974 1760 30000
rect 1884 30918 1918 30944
rect 1884 30910 1918 30918
rect 1884 30850 1918 30872
rect 1884 30838 1918 30850
rect 1884 30782 1918 30800
rect 1884 30766 1918 30782
rect 1884 30714 1918 30728
rect 1884 30694 1918 30714
rect 1884 30646 1918 30656
rect 1884 30622 1918 30646
rect 1884 30578 1918 30584
rect 1884 30550 1918 30578
rect 1884 30510 1918 30512
rect 1884 30478 1918 30510
rect 1884 30408 1918 30440
rect 1884 30406 1918 30408
rect 1884 30340 1918 30368
rect 1884 30334 1918 30340
rect 1884 30272 1918 30296
rect 1884 30262 1918 30272
rect 1884 30204 1918 30224
rect 1884 30190 1918 30204
rect 1884 30136 1918 30152
rect 1884 30118 1918 30136
rect 1884 30068 1918 30080
rect 1884 30046 1918 30068
rect 1884 30000 1918 30008
rect 1884 29974 1918 30000
rect 2042 30918 2076 30944
rect 2042 30910 2076 30918
rect 2042 30850 2076 30872
rect 2042 30838 2076 30850
rect 2042 30782 2076 30800
rect 2042 30766 2076 30782
rect 2042 30714 2076 30728
rect 2042 30694 2076 30714
rect 2042 30646 2076 30656
rect 2042 30622 2076 30646
rect 2042 30578 2076 30584
rect 2042 30550 2076 30578
rect 2042 30510 2076 30512
rect 2042 30478 2076 30510
rect 2042 30408 2076 30440
rect 2042 30406 2076 30408
rect 2042 30340 2076 30368
rect 2042 30334 2076 30340
rect 2042 30272 2076 30296
rect 2042 30262 2076 30272
rect 2042 30204 2076 30224
rect 2042 30190 2076 30204
rect 2042 30136 2076 30152
rect 2042 30118 2076 30136
rect 2042 30068 2076 30080
rect 2042 30046 2076 30068
rect 2042 30000 2076 30008
rect 2042 29974 2076 30000
rect 2200 30918 2234 30944
rect 2200 30910 2234 30918
rect 2200 30850 2234 30872
rect 2200 30838 2234 30850
rect 2200 30782 2234 30800
rect 2200 30766 2234 30782
rect 2200 30714 2234 30728
rect 2200 30694 2234 30714
rect 2200 30646 2234 30656
rect 2200 30622 2234 30646
rect 2200 30578 2234 30584
rect 2200 30550 2234 30578
rect 2200 30510 2234 30512
rect 2200 30478 2234 30510
rect 2200 30408 2234 30440
rect 2200 30406 2234 30408
rect 2200 30340 2234 30368
rect 2200 30334 2234 30340
rect 2200 30272 2234 30296
rect 2200 30262 2234 30272
rect 2200 30204 2234 30224
rect 2200 30190 2234 30204
rect 2200 30136 2234 30152
rect 2200 30118 2234 30136
rect 2200 30068 2234 30080
rect 2200 30046 2234 30068
rect 2200 30000 2234 30008
rect 2200 29974 2234 30000
rect 2358 30918 2392 30944
rect 2358 30910 2392 30918
rect 2358 30850 2392 30872
rect 2358 30838 2392 30850
rect 2358 30782 2392 30800
rect 2358 30766 2392 30782
rect 2358 30714 2392 30728
rect 2358 30694 2392 30714
rect 2358 30646 2392 30656
rect 2358 30622 2392 30646
rect 2358 30578 2392 30584
rect 2358 30550 2392 30578
rect 2358 30510 2392 30512
rect 2358 30478 2392 30510
rect 2358 30408 2392 30440
rect 2358 30406 2392 30408
rect 2358 30340 2392 30368
rect 2358 30334 2392 30340
rect 2358 30272 2392 30296
rect 2358 30262 2392 30272
rect 2358 30204 2392 30224
rect 2358 30190 2392 30204
rect 2358 30136 2392 30152
rect 2358 30118 2392 30136
rect 2358 30068 2392 30080
rect 2358 30046 2392 30068
rect 2358 30000 2392 30008
rect 2358 29974 2392 30000
rect 2516 30918 2550 30944
rect 2516 30910 2550 30918
rect 2516 30850 2550 30872
rect 2516 30838 2550 30850
rect 2516 30782 2550 30800
rect 2516 30766 2550 30782
rect 2516 30714 2550 30728
rect 2516 30694 2550 30714
rect 2516 30646 2550 30656
rect 2516 30622 2550 30646
rect 2516 30578 2550 30584
rect 2516 30550 2550 30578
rect 2516 30510 2550 30512
rect 2516 30478 2550 30510
rect 2516 30408 2550 30440
rect 2516 30406 2550 30408
rect 2516 30340 2550 30368
rect 2516 30334 2550 30340
rect 2516 30272 2550 30296
rect 2516 30262 2550 30272
rect 2516 30204 2550 30224
rect 2516 30190 2550 30204
rect 2516 30136 2550 30152
rect 2516 30118 2550 30136
rect 2516 30068 2550 30080
rect 2516 30046 2550 30068
rect 2516 30000 2550 30008
rect 2516 29974 2550 30000
rect 2674 30918 2708 30944
rect 2674 30910 2708 30918
rect 2674 30850 2708 30872
rect 2674 30838 2708 30850
rect 2674 30782 2708 30800
rect 2674 30766 2708 30782
rect 2674 30714 2708 30728
rect 2674 30694 2708 30714
rect 2674 30646 2708 30656
rect 2674 30622 2708 30646
rect 2674 30578 2708 30584
rect 2674 30550 2708 30578
rect 2674 30510 2708 30512
rect 2674 30478 2708 30510
rect 2674 30408 2708 30440
rect 2674 30406 2708 30408
rect 2674 30340 2708 30368
rect 2674 30334 2708 30340
rect 2674 30272 2708 30296
rect 2674 30262 2708 30272
rect 2674 30204 2708 30224
rect 2674 30190 2708 30204
rect 2674 30136 2708 30152
rect 2674 30118 2708 30136
rect 2674 30068 2708 30080
rect 2674 30046 2708 30068
rect 2674 30000 2708 30008
rect 2674 29974 2708 30000
rect 2832 30918 2866 30944
rect 2832 30910 2866 30918
rect 2832 30850 2866 30872
rect 2832 30838 2866 30850
rect 2832 30782 2866 30800
rect 2832 30766 2866 30782
rect 2832 30714 2866 30728
rect 2832 30694 2866 30714
rect 2832 30646 2866 30656
rect 2832 30622 2866 30646
rect 2832 30578 2866 30584
rect 2832 30550 2866 30578
rect 2832 30510 2866 30512
rect 2832 30478 2866 30510
rect 2832 30408 2866 30440
rect 2832 30406 2866 30408
rect 2832 30340 2866 30368
rect 2832 30334 2866 30340
rect 2832 30272 2866 30296
rect 2832 30262 2866 30272
rect 2832 30204 2866 30224
rect 2832 30190 2866 30204
rect 2832 30136 2866 30152
rect 2832 30118 2866 30136
rect 2832 30068 2866 30080
rect 2832 30046 2866 30068
rect 2832 30000 2866 30008
rect 2832 29974 2866 30000
rect 2990 30918 3024 30944
rect 2990 30910 3024 30918
rect 2990 30850 3024 30872
rect 2990 30838 3024 30850
rect 2990 30782 3024 30800
rect 2990 30766 3024 30782
rect 2990 30714 3024 30728
rect 2990 30694 3024 30714
rect 2990 30646 3024 30656
rect 2990 30622 3024 30646
rect 2990 30578 3024 30584
rect 2990 30550 3024 30578
rect 2990 30510 3024 30512
rect 2990 30478 3024 30510
rect 2990 30408 3024 30440
rect 2990 30406 3024 30408
rect 2990 30340 3024 30368
rect 2990 30334 3024 30340
rect 2990 30272 3024 30296
rect 2990 30262 3024 30272
rect 2990 30204 3024 30224
rect 2990 30190 3024 30204
rect 2990 30136 3024 30152
rect 2990 30118 3024 30136
rect 2990 30068 3024 30080
rect 2990 30046 3024 30068
rect 2990 30000 3024 30008
rect 2990 29974 3024 30000
rect 3148 30918 3182 30944
rect 3148 30910 3182 30918
rect 3148 30850 3182 30872
rect 3148 30838 3182 30850
rect 3148 30782 3182 30800
rect 3148 30766 3182 30782
rect 3148 30714 3182 30728
rect 3148 30694 3182 30714
rect 3148 30646 3182 30656
rect 3148 30622 3182 30646
rect 3148 30578 3182 30584
rect 3148 30550 3182 30578
rect 3148 30510 3182 30512
rect 3148 30478 3182 30510
rect 3148 30408 3182 30440
rect 3148 30406 3182 30408
rect 3148 30340 3182 30368
rect 3148 30334 3182 30340
rect 3148 30272 3182 30296
rect 3148 30262 3182 30272
rect 3148 30204 3182 30224
rect 3148 30190 3182 30204
rect 3148 30136 3182 30152
rect 3148 30118 3182 30136
rect 3148 30068 3182 30080
rect 3148 30046 3182 30068
rect 3148 30000 3182 30008
rect 3148 29974 3182 30000
rect 4293 30782 4687 31896
rect 6724 30782 7118 31896
rect -3093 29878 -3059 29912
rect -2935 29878 -2901 29912
rect -2777 29878 -2743 29912
rect -2619 29878 -2585 29912
rect -2461 29878 -2427 29912
rect -2303 29878 -2269 29912
rect -2145 29878 -2111 29912
rect -1987 29878 -1953 29912
rect -1829 29878 -1795 29912
rect -1671 29878 -1637 29912
rect -1513 29878 -1479 29912
rect -1355 29878 -1321 29912
rect -1197 29878 -1163 29912
rect -1039 29878 -1005 29912
rect -881 29878 -847 29912
rect -723 29878 -689 29912
rect -565 29878 -531 29912
rect -407 29878 -373 29912
rect -249 29878 -215 29912
rect -91 29878 -57 29912
rect 67 29878 101 29912
rect 225 29878 259 29912
rect 383 29878 417 29912
rect 541 29878 575 29912
rect 699 29878 733 29912
rect 857 29878 891 29912
rect 1015 29878 1049 29912
rect 1173 29878 1207 29912
rect 1331 29878 1365 29912
rect 1489 29878 1523 29912
rect 1647 29878 1681 29912
rect 1805 29878 1839 29912
rect 1963 29878 1997 29912
rect 2121 29878 2155 29912
rect 2279 29878 2313 29912
rect 2437 29878 2471 29912
rect 2595 29878 2629 29912
rect 2753 29878 2787 29912
rect 2911 29878 2945 29912
rect 3069 29878 3103 29912
rect -1596 29776 -1576 29810
rect -1576 29776 -1562 29810
rect -1524 29776 -1508 29810
rect -1508 29776 -1490 29810
rect -1452 29776 -1440 29810
rect -1440 29776 -1418 29810
rect -1380 29776 -1372 29810
rect -1372 29776 -1346 29810
rect -1308 29776 -1304 29810
rect -1304 29776 -1274 29810
rect -1236 29776 -1202 29810
rect -1164 29776 -1134 29810
rect -1134 29776 -1130 29810
rect -1092 29776 -1066 29810
rect -1066 29776 -1058 29810
rect -1020 29776 -998 29810
rect -998 29776 -986 29810
rect -948 29776 -930 29810
rect -930 29776 -914 29810
rect -876 29776 -862 29810
rect -862 29776 -842 29810
rect -804 29776 -794 29810
rect -794 29776 -770 29810
rect -732 29776 -726 29810
rect -726 29776 -698 29810
rect -660 29776 -658 29810
rect -658 29776 -626 29810
rect -588 29776 -556 29810
rect -556 29776 -554 29810
rect -516 29776 -488 29810
rect -488 29776 -482 29810
rect -444 29776 -420 29810
rect -420 29776 -410 29810
rect -372 29776 -352 29810
rect -352 29776 -338 29810
rect -300 29776 -284 29810
rect -284 29776 -266 29810
rect -228 29776 -216 29810
rect -216 29776 -194 29810
rect -156 29776 -148 29810
rect -148 29776 -122 29810
rect -84 29776 -80 29810
rect -80 29776 -50 29810
rect -12 29776 22 29810
rect 60 29776 90 29810
rect 90 29776 94 29810
rect 132 29776 158 29810
rect 158 29776 166 29810
rect 204 29776 226 29810
rect 226 29776 238 29810
rect 276 29776 294 29810
rect 294 29776 310 29810
rect 348 29776 362 29810
rect 362 29776 382 29810
rect 420 29776 430 29810
rect 430 29776 454 29810
rect 492 29776 498 29810
rect 498 29776 526 29810
rect 564 29776 566 29810
rect 566 29776 598 29810
rect 636 29776 668 29810
rect 668 29776 670 29810
rect 708 29776 736 29810
rect 736 29776 742 29810
rect 780 29776 804 29810
rect 804 29776 814 29810
rect 852 29776 872 29810
rect 872 29776 886 29810
rect 924 29776 940 29810
rect 940 29776 958 29810
rect 996 29776 1008 29810
rect 1008 29776 1030 29810
rect 1068 29776 1076 29810
rect 1076 29776 1102 29810
rect 1140 29776 1144 29810
rect 1144 29776 1174 29810
rect 1212 29776 1246 29810
rect 1284 29776 1314 29810
rect 1314 29776 1318 29810
rect 1356 29776 1382 29810
rect 1382 29776 1390 29810
rect 1428 29776 1450 29810
rect 1450 29776 1462 29810
rect 1500 29776 1518 29810
rect 1518 29776 1534 29810
rect 1572 29776 1586 29810
rect 1586 29776 1606 29810
rect -6350 29166 -6190 29190
rect -6000 29166 -5840 29190
rect -5630 29166 -5470 29190
rect -841 29438 -829 29472
rect -829 29438 -807 29472
rect -769 29438 -761 29472
rect -761 29438 -735 29472
rect -697 29438 -693 29472
rect -693 29438 -663 29472
rect -625 29438 -591 29472
rect -553 29438 -523 29472
rect -523 29438 -519 29472
rect -481 29438 -455 29472
rect -455 29438 -447 29472
rect -409 29438 -387 29472
rect -387 29438 -375 29472
rect -337 29438 -319 29472
rect -319 29438 -303 29472
rect -265 29438 -251 29472
rect -251 29438 -231 29472
rect -193 29438 -183 29472
rect -183 29438 -159 29472
rect -121 29438 -115 29472
rect -115 29438 -87 29472
rect -49 29438 -47 29472
rect -47 29438 -15 29472
rect 23 29438 55 29472
rect 55 29438 57 29472
rect 95 29438 123 29472
rect 123 29438 129 29472
rect 167 29438 191 29472
rect 191 29438 201 29472
rect 239 29438 259 29472
rect 259 29438 273 29472
rect 311 29438 327 29472
rect 327 29438 345 29472
rect 383 29438 395 29472
rect 395 29438 417 29472
rect 455 29438 463 29472
rect 463 29438 489 29472
rect 527 29438 531 29472
rect 531 29438 561 29472
rect 599 29438 633 29472
rect 671 29438 701 29472
rect 701 29438 705 29472
rect 743 29438 769 29472
rect 769 29438 777 29472
rect 815 29438 837 29472
rect 837 29438 849 29472
rect -1593 29336 -1559 29370
rect -1435 29336 -1401 29370
rect -1277 29336 -1243 29370
rect -1119 29336 -1085 29370
rect -961 29336 -927 29370
rect -803 29336 -769 29370
rect -645 29336 -611 29370
rect -487 29336 -453 29370
rect -329 29336 -295 29370
rect -171 29336 -137 29370
rect -13 29336 21 29370
rect 145 29336 179 29370
rect 303 29336 337 29370
rect 461 29336 495 29370
rect 619 29336 653 29370
rect 777 29336 811 29370
rect 935 29336 969 29370
rect 1093 29336 1127 29370
rect 1251 29336 1285 29370
rect 1409 29336 1443 29370
rect 1567 29336 1601 29370
rect -6350 29140 -6190 29166
rect -6000 29140 -5840 29166
rect -5630 29140 -5470 29166
rect -1672 29248 -1638 29274
rect -1672 29240 -1638 29248
rect -1672 29180 -1638 29202
rect -1672 29168 -1638 29180
rect -1672 29112 -1638 29130
rect -1672 29096 -1638 29112
rect -1672 29044 -1638 29058
rect -1672 29024 -1638 29044
rect -1672 28976 -1638 28986
rect -1672 28952 -1638 28976
rect -1672 28908 -1638 28914
rect -1672 28880 -1638 28908
rect -1672 28840 -1638 28842
rect -1672 28808 -1638 28840
rect -1672 28738 -1638 28770
rect -1672 28736 -1638 28738
rect -1672 28670 -1638 28698
rect -1672 28664 -1638 28670
rect -1672 28602 -1638 28626
rect -1672 28592 -1638 28602
rect -1672 28534 -1638 28554
rect -1672 28520 -1638 28534
rect -1672 28466 -1638 28482
rect -1672 28448 -1638 28466
rect -1672 28398 -1638 28410
rect -1672 28376 -1638 28398
rect -1672 28330 -1638 28338
rect -1672 28304 -1638 28330
rect -1514 29248 -1480 29274
rect -1514 29240 -1480 29248
rect -1514 29180 -1480 29202
rect -1514 29168 -1480 29180
rect -1514 29112 -1480 29130
rect -1514 29096 -1480 29112
rect -1514 29044 -1480 29058
rect -1514 29024 -1480 29044
rect -1514 28976 -1480 28986
rect -1514 28952 -1480 28976
rect -1514 28908 -1480 28914
rect -1514 28880 -1480 28908
rect -1514 28840 -1480 28842
rect -1514 28808 -1480 28840
rect -1514 28738 -1480 28770
rect -1514 28736 -1480 28738
rect -1514 28670 -1480 28698
rect -1514 28664 -1480 28670
rect -1514 28602 -1480 28626
rect -1514 28592 -1480 28602
rect -1514 28534 -1480 28554
rect -1514 28520 -1480 28534
rect -1514 28466 -1480 28482
rect -1514 28448 -1480 28466
rect -1514 28398 -1480 28410
rect -1514 28376 -1480 28398
rect -1514 28330 -1480 28338
rect -1514 28304 -1480 28330
rect -1356 29248 -1322 29274
rect -1356 29240 -1322 29248
rect -1356 29180 -1322 29202
rect -1356 29168 -1322 29180
rect -1356 29112 -1322 29130
rect -1356 29096 -1322 29112
rect -1356 29044 -1322 29058
rect -1356 29024 -1322 29044
rect -1356 28976 -1322 28986
rect -1356 28952 -1322 28976
rect -1356 28908 -1322 28914
rect -1356 28880 -1322 28908
rect -1356 28840 -1322 28842
rect -1356 28808 -1322 28840
rect -1356 28738 -1322 28770
rect -1356 28736 -1322 28738
rect -1356 28670 -1322 28698
rect -1356 28664 -1322 28670
rect -1356 28602 -1322 28626
rect -1356 28592 -1322 28602
rect -1356 28534 -1322 28554
rect -1356 28520 -1322 28534
rect -1356 28466 -1322 28482
rect -1356 28448 -1322 28466
rect -1356 28398 -1322 28410
rect -1356 28376 -1322 28398
rect -1356 28330 -1322 28338
rect -1356 28304 -1322 28330
rect -1198 29248 -1164 29274
rect -1198 29240 -1164 29248
rect -1198 29180 -1164 29202
rect -1198 29168 -1164 29180
rect -1198 29112 -1164 29130
rect -1198 29096 -1164 29112
rect -1198 29044 -1164 29058
rect -1198 29024 -1164 29044
rect -1198 28976 -1164 28986
rect -1198 28952 -1164 28976
rect -1198 28908 -1164 28914
rect -1198 28880 -1164 28908
rect -1198 28840 -1164 28842
rect -1198 28808 -1164 28840
rect -1198 28738 -1164 28770
rect -1198 28736 -1164 28738
rect -1198 28670 -1164 28698
rect -1198 28664 -1164 28670
rect -1198 28602 -1164 28626
rect -1198 28592 -1164 28602
rect -1198 28534 -1164 28554
rect -1198 28520 -1164 28534
rect -1198 28466 -1164 28482
rect -1198 28448 -1164 28466
rect -1198 28398 -1164 28410
rect -1198 28376 -1164 28398
rect -1198 28330 -1164 28338
rect -1198 28304 -1164 28330
rect -1040 29248 -1006 29274
rect -1040 29240 -1006 29248
rect -1040 29180 -1006 29202
rect -1040 29168 -1006 29180
rect -1040 29112 -1006 29130
rect -1040 29096 -1006 29112
rect -1040 29044 -1006 29058
rect -1040 29024 -1006 29044
rect -1040 28976 -1006 28986
rect -1040 28952 -1006 28976
rect -1040 28908 -1006 28914
rect -1040 28880 -1006 28908
rect -1040 28840 -1006 28842
rect -1040 28808 -1006 28840
rect -1040 28738 -1006 28770
rect -1040 28736 -1006 28738
rect -1040 28670 -1006 28698
rect -1040 28664 -1006 28670
rect -1040 28602 -1006 28626
rect -1040 28592 -1006 28602
rect -1040 28534 -1006 28554
rect -1040 28520 -1006 28534
rect -1040 28466 -1006 28482
rect -1040 28448 -1006 28466
rect -1040 28398 -1006 28410
rect -1040 28376 -1006 28398
rect -1040 28330 -1006 28338
rect -1040 28304 -1006 28330
rect -882 29248 -848 29274
rect -882 29240 -848 29248
rect -882 29180 -848 29202
rect -882 29168 -848 29180
rect -882 29112 -848 29130
rect -882 29096 -848 29112
rect -882 29044 -848 29058
rect -882 29024 -848 29044
rect -882 28976 -848 28986
rect -882 28952 -848 28976
rect -882 28908 -848 28914
rect -882 28880 -848 28908
rect -882 28840 -848 28842
rect -882 28808 -848 28840
rect -882 28738 -848 28770
rect -882 28736 -848 28738
rect -882 28670 -848 28698
rect -882 28664 -848 28670
rect -882 28602 -848 28626
rect -882 28592 -848 28602
rect -882 28534 -848 28554
rect -882 28520 -848 28534
rect -882 28466 -848 28482
rect -882 28448 -848 28466
rect -882 28398 -848 28410
rect -882 28376 -848 28398
rect -882 28330 -848 28338
rect -882 28304 -848 28330
rect -724 29248 -690 29274
rect -724 29240 -690 29248
rect -724 29180 -690 29202
rect -724 29168 -690 29180
rect -724 29112 -690 29130
rect -724 29096 -690 29112
rect -724 29044 -690 29058
rect -724 29024 -690 29044
rect -724 28976 -690 28986
rect -724 28952 -690 28976
rect -724 28908 -690 28914
rect -724 28880 -690 28908
rect -724 28840 -690 28842
rect -724 28808 -690 28840
rect -724 28738 -690 28770
rect -724 28736 -690 28738
rect -724 28670 -690 28698
rect -724 28664 -690 28670
rect -724 28602 -690 28626
rect -724 28592 -690 28602
rect -724 28534 -690 28554
rect -724 28520 -690 28534
rect -724 28466 -690 28482
rect -724 28448 -690 28466
rect -724 28398 -690 28410
rect -724 28376 -690 28398
rect -724 28330 -690 28338
rect -724 28304 -690 28330
rect -566 29248 -532 29274
rect -566 29240 -532 29248
rect -566 29180 -532 29202
rect -566 29168 -532 29180
rect -566 29112 -532 29130
rect -566 29096 -532 29112
rect -566 29044 -532 29058
rect -566 29024 -532 29044
rect -566 28976 -532 28986
rect -566 28952 -532 28976
rect -566 28908 -532 28914
rect -566 28880 -532 28908
rect -566 28840 -532 28842
rect -566 28808 -532 28840
rect -566 28738 -532 28770
rect -566 28736 -532 28738
rect -566 28670 -532 28698
rect -566 28664 -532 28670
rect -566 28602 -532 28626
rect -566 28592 -532 28602
rect -566 28534 -532 28554
rect -566 28520 -532 28534
rect -566 28466 -532 28482
rect -566 28448 -532 28466
rect -566 28398 -532 28410
rect -566 28376 -532 28398
rect -566 28330 -532 28338
rect -566 28304 -532 28330
rect -408 29248 -374 29274
rect -408 29240 -374 29248
rect -408 29180 -374 29202
rect -408 29168 -374 29180
rect -408 29112 -374 29130
rect -408 29096 -374 29112
rect -408 29044 -374 29058
rect -408 29024 -374 29044
rect -408 28976 -374 28986
rect -408 28952 -374 28976
rect -408 28908 -374 28914
rect -408 28880 -374 28908
rect -408 28840 -374 28842
rect -408 28808 -374 28840
rect -408 28738 -374 28770
rect -408 28736 -374 28738
rect -408 28670 -374 28698
rect -408 28664 -374 28670
rect -408 28602 -374 28626
rect -408 28592 -374 28602
rect -408 28534 -374 28554
rect -408 28520 -374 28534
rect -408 28466 -374 28482
rect -408 28448 -374 28466
rect -408 28398 -374 28410
rect -408 28376 -374 28398
rect -408 28330 -374 28338
rect -408 28304 -374 28330
rect -250 29248 -216 29274
rect -250 29240 -216 29248
rect -250 29180 -216 29202
rect -250 29168 -216 29180
rect -250 29112 -216 29130
rect -250 29096 -216 29112
rect -250 29044 -216 29058
rect -250 29024 -216 29044
rect -250 28976 -216 28986
rect -250 28952 -216 28976
rect -250 28908 -216 28914
rect -250 28880 -216 28908
rect -250 28840 -216 28842
rect -250 28808 -216 28840
rect -250 28738 -216 28770
rect -250 28736 -216 28738
rect -250 28670 -216 28698
rect -250 28664 -216 28670
rect -250 28602 -216 28626
rect -250 28592 -216 28602
rect -250 28534 -216 28554
rect -250 28520 -216 28534
rect -250 28466 -216 28482
rect -250 28448 -216 28466
rect -250 28398 -216 28410
rect -250 28376 -216 28398
rect -250 28330 -216 28338
rect -250 28304 -216 28330
rect -92 29248 -58 29274
rect -92 29240 -58 29248
rect -92 29180 -58 29202
rect -92 29168 -58 29180
rect -92 29112 -58 29130
rect -92 29096 -58 29112
rect -92 29044 -58 29058
rect -92 29024 -58 29044
rect -92 28976 -58 28986
rect -92 28952 -58 28976
rect -92 28908 -58 28914
rect -92 28880 -58 28908
rect -92 28840 -58 28842
rect -92 28808 -58 28840
rect -92 28738 -58 28770
rect -92 28736 -58 28738
rect -92 28670 -58 28698
rect -92 28664 -58 28670
rect -92 28602 -58 28626
rect -92 28592 -58 28602
rect -92 28534 -58 28554
rect -92 28520 -58 28534
rect -92 28466 -58 28482
rect -92 28448 -58 28466
rect -92 28398 -58 28410
rect -92 28376 -58 28398
rect -92 28330 -58 28338
rect -92 28304 -58 28330
rect 66 29248 100 29274
rect 66 29240 100 29248
rect 66 29180 100 29202
rect 66 29168 100 29180
rect 66 29112 100 29130
rect 66 29096 100 29112
rect 66 29044 100 29058
rect 66 29024 100 29044
rect 66 28976 100 28986
rect 66 28952 100 28976
rect 66 28908 100 28914
rect 66 28880 100 28908
rect 66 28840 100 28842
rect 66 28808 100 28840
rect 66 28738 100 28770
rect 66 28736 100 28738
rect 66 28670 100 28698
rect 66 28664 100 28670
rect 66 28602 100 28626
rect 66 28592 100 28602
rect 66 28534 100 28554
rect 66 28520 100 28534
rect 66 28466 100 28482
rect 66 28448 100 28466
rect 66 28398 100 28410
rect 66 28376 100 28398
rect 66 28330 100 28338
rect 66 28304 100 28330
rect 224 29248 258 29274
rect 224 29240 258 29248
rect 224 29180 258 29202
rect 224 29168 258 29180
rect 224 29112 258 29130
rect 224 29096 258 29112
rect 224 29044 258 29058
rect 224 29024 258 29044
rect 224 28976 258 28986
rect 224 28952 258 28976
rect 224 28908 258 28914
rect 224 28880 258 28908
rect 224 28840 258 28842
rect 224 28808 258 28840
rect 224 28738 258 28770
rect 224 28736 258 28738
rect 224 28670 258 28698
rect 224 28664 258 28670
rect 224 28602 258 28626
rect 224 28592 258 28602
rect 224 28534 258 28554
rect 224 28520 258 28534
rect 224 28466 258 28482
rect 224 28448 258 28466
rect 224 28398 258 28410
rect 224 28376 258 28398
rect 224 28330 258 28338
rect 224 28304 258 28330
rect 382 29248 416 29274
rect 382 29240 416 29248
rect 382 29180 416 29202
rect 382 29168 416 29180
rect 382 29112 416 29130
rect 382 29096 416 29112
rect 382 29044 416 29058
rect 382 29024 416 29044
rect 382 28976 416 28986
rect 382 28952 416 28976
rect 382 28908 416 28914
rect 382 28880 416 28908
rect 382 28840 416 28842
rect 382 28808 416 28840
rect 382 28738 416 28770
rect 382 28736 416 28738
rect 382 28670 416 28698
rect 382 28664 416 28670
rect 382 28602 416 28626
rect 382 28592 416 28602
rect 382 28534 416 28554
rect 382 28520 416 28534
rect 382 28466 416 28482
rect 382 28448 416 28466
rect 382 28398 416 28410
rect 382 28376 416 28398
rect 382 28330 416 28338
rect 382 28304 416 28330
rect 540 29248 574 29274
rect 540 29240 574 29248
rect 540 29180 574 29202
rect 540 29168 574 29180
rect 540 29112 574 29130
rect 540 29096 574 29112
rect 540 29044 574 29058
rect 540 29024 574 29044
rect 540 28976 574 28986
rect 540 28952 574 28976
rect 540 28908 574 28914
rect 540 28880 574 28908
rect 540 28840 574 28842
rect 540 28808 574 28840
rect 540 28738 574 28770
rect 540 28736 574 28738
rect 540 28670 574 28698
rect 540 28664 574 28670
rect 540 28602 574 28626
rect 540 28592 574 28602
rect 540 28534 574 28554
rect 540 28520 574 28534
rect 540 28466 574 28482
rect 540 28448 574 28466
rect 540 28398 574 28410
rect 540 28376 574 28398
rect 540 28330 574 28338
rect 540 28304 574 28330
rect 698 29248 732 29274
rect 698 29240 732 29248
rect 698 29180 732 29202
rect 698 29168 732 29180
rect 698 29112 732 29130
rect 698 29096 732 29112
rect 698 29044 732 29058
rect 698 29024 732 29044
rect 698 28976 732 28986
rect 698 28952 732 28976
rect 698 28908 732 28914
rect 698 28880 732 28908
rect 698 28840 732 28842
rect 698 28808 732 28840
rect 698 28738 732 28770
rect 698 28736 732 28738
rect 698 28670 732 28698
rect 698 28664 732 28670
rect 698 28602 732 28626
rect 698 28592 732 28602
rect 698 28534 732 28554
rect 698 28520 732 28534
rect 698 28466 732 28482
rect 698 28448 732 28466
rect 698 28398 732 28410
rect 698 28376 732 28398
rect 698 28330 732 28338
rect 698 28304 732 28330
rect 856 29248 890 29274
rect 856 29240 890 29248
rect 856 29180 890 29202
rect 856 29168 890 29180
rect 856 29112 890 29130
rect 856 29096 890 29112
rect 856 29044 890 29058
rect 856 29024 890 29044
rect 856 28976 890 28986
rect 856 28952 890 28976
rect 856 28908 890 28914
rect 856 28880 890 28908
rect 856 28840 890 28842
rect 856 28808 890 28840
rect 856 28738 890 28770
rect 856 28736 890 28738
rect 856 28670 890 28698
rect 856 28664 890 28670
rect 856 28602 890 28626
rect 856 28592 890 28602
rect 856 28534 890 28554
rect 856 28520 890 28534
rect 856 28466 890 28482
rect 856 28448 890 28466
rect 856 28398 890 28410
rect 856 28376 890 28398
rect 856 28330 890 28338
rect 856 28304 890 28330
rect 1014 29248 1048 29274
rect 1014 29240 1048 29248
rect 1014 29180 1048 29202
rect 1014 29168 1048 29180
rect 1014 29112 1048 29130
rect 1014 29096 1048 29112
rect 1014 29044 1048 29058
rect 1014 29024 1048 29044
rect 1014 28976 1048 28986
rect 1014 28952 1048 28976
rect 1014 28908 1048 28914
rect 1014 28880 1048 28908
rect 1014 28840 1048 28842
rect 1014 28808 1048 28840
rect 1014 28738 1048 28770
rect 1014 28736 1048 28738
rect 1014 28670 1048 28698
rect 1014 28664 1048 28670
rect 1014 28602 1048 28626
rect 1014 28592 1048 28602
rect 1014 28534 1048 28554
rect 1014 28520 1048 28534
rect 1014 28466 1048 28482
rect 1014 28448 1048 28466
rect 1014 28398 1048 28410
rect 1014 28376 1048 28398
rect 1014 28330 1048 28338
rect 1014 28304 1048 28330
rect 1172 29248 1206 29274
rect 1172 29240 1206 29248
rect 1172 29180 1206 29202
rect 1172 29168 1206 29180
rect 1172 29112 1206 29130
rect 1172 29096 1206 29112
rect 1172 29044 1206 29058
rect 1172 29024 1206 29044
rect 1172 28976 1206 28986
rect 1172 28952 1206 28976
rect 1172 28908 1206 28914
rect 1172 28880 1206 28908
rect 1172 28840 1206 28842
rect 1172 28808 1206 28840
rect 1172 28738 1206 28770
rect 1172 28736 1206 28738
rect 1172 28670 1206 28698
rect 1172 28664 1206 28670
rect 1172 28602 1206 28626
rect 1172 28592 1206 28602
rect 1172 28534 1206 28554
rect 1172 28520 1206 28534
rect 1172 28466 1206 28482
rect 1172 28448 1206 28466
rect 1172 28398 1206 28410
rect 1172 28376 1206 28398
rect 1172 28330 1206 28338
rect 1172 28304 1206 28330
rect 1330 29248 1364 29274
rect 1330 29240 1364 29248
rect 1330 29180 1364 29202
rect 1330 29168 1364 29180
rect 1330 29112 1364 29130
rect 1330 29096 1364 29112
rect 1330 29044 1364 29058
rect 1330 29024 1364 29044
rect 1330 28976 1364 28986
rect 1330 28952 1364 28976
rect 1330 28908 1364 28914
rect 1330 28880 1364 28908
rect 1330 28840 1364 28842
rect 1330 28808 1364 28840
rect 1330 28738 1364 28770
rect 1330 28736 1364 28738
rect 1330 28670 1364 28698
rect 1330 28664 1364 28670
rect 1330 28602 1364 28626
rect 1330 28592 1364 28602
rect 1330 28534 1364 28554
rect 1330 28520 1364 28534
rect 1330 28466 1364 28482
rect 1330 28448 1364 28466
rect 1330 28398 1364 28410
rect 1330 28376 1364 28398
rect 1330 28330 1364 28338
rect 1330 28304 1364 28330
rect 1488 29248 1522 29274
rect 1488 29240 1522 29248
rect 1488 29180 1522 29202
rect 1488 29168 1522 29180
rect 1488 29112 1522 29130
rect 1488 29096 1522 29112
rect 1488 29044 1522 29058
rect 1488 29024 1522 29044
rect 1488 28976 1522 28986
rect 1488 28952 1522 28976
rect 1488 28908 1522 28914
rect 1488 28880 1522 28908
rect 1488 28840 1522 28842
rect 1488 28808 1522 28840
rect 1488 28738 1522 28770
rect 1488 28736 1522 28738
rect 1488 28670 1522 28698
rect 1488 28664 1522 28670
rect 1488 28602 1522 28626
rect 1488 28592 1522 28602
rect 1488 28534 1522 28554
rect 1488 28520 1522 28534
rect 1488 28466 1522 28482
rect 1488 28448 1522 28466
rect 1488 28398 1522 28410
rect 1488 28376 1522 28398
rect 1488 28330 1522 28338
rect 1488 28304 1522 28330
rect 1646 29248 1680 29274
rect 1646 29240 1680 29248
rect 1646 29180 1680 29202
rect 1646 29168 1680 29180
rect 1646 29112 1680 29130
rect 1646 29096 1680 29112
rect 1646 29044 1680 29058
rect 1646 29024 1680 29044
rect 1646 28976 1680 28986
rect 1646 28952 1680 28976
rect 1646 28908 1680 28914
rect 1646 28880 1680 28908
rect 1646 28840 1680 28842
rect 1646 28808 1680 28840
rect 1646 28738 1680 28770
rect 1646 28736 1680 28738
rect 1646 28670 1680 28698
rect 1646 28664 1680 28670
rect 1646 28602 1680 28626
rect 1646 28592 1680 28602
rect 1646 28534 1680 28554
rect 1646 28520 1680 28534
rect 1646 28466 1680 28482
rect 1646 28448 1680 28466
rect 1646 28398 1680 28410
rect 1646 28376 1680 28398
rect 1646 28330 1680 28338
rect 1646 28304 1680 28330
rect 4293 29302 4687 30416
rect 6724 29302 7118 30416
rect 5438 29156 5451 29180
rect 5451 29156 5485 29180
rect 5485 29156 5519 29180
rect 5519 29156 5553 29180
rect 5553 29156 5587 29180
rect 5587 29156 5621 29180
rect 5621 29156 5638 29180
rect 6098 29156 6131 29180
rect 6131 29156 6165 29180
rect 6165 29156 6199 29180
rect 6199 29156 6233 29180
rect 6233 29156 6267 29180
rect 6267 29156 6298 29180
rect 5438 29120 5638 29156
rect 6098 29120 6298 29156
rect -1593 28208 -1559 28242
rect -1435 28208 -1401 28242
rect -1277 28208 -1243 28242
rect -1119 28208 -1085 28242
rect -961 28208 -927 28242
rect -803 28208 -769 28242
rect -645 28208 -611 28242
rect -487 28208 -453 28242
rect -329 28208 -295 28242
rect -171 28208 -137 28242
rect -13 28208 21 28242
rect 145 28208 179 28242
rect 303 28208 337 28242
rect 461 28208 495 28242
rect 619 28208 653 28242
rect 777 28208 811 28242
rect 935 28208 969 28242
rect 1093 28208 1127 28242
rect 1251 28208 1285 28242
rect 1409 28208 1443 28242
rect 1567 28208 1601 28242
rect -996 28106 -965 28109
rect -965 28106 -931 28109
rect -931 28106 -897 28109
rect -897 28106 -863 28109
rect -863 28106 -829 28109
rect -829 28106 -795 28109
rect -795 28106 -761 28109
rect -761 28106 -727 28109
rect -727 28106 -693 28109
rect -693 28106 -659 28109
rect -659 28106 -625 28109
rect -625 28106 -591 28109
rect -591 28106 -557 28109
rect -557 28106 -523 28109
rect -523 28106 -489 28109
rect -489 28106 -458 28109
rect 474 28106 497 28109
rect 497 28106 531 28109
rect 531 28106 565 28109
rect 565 28106 599 28109
rect 599 28106 633 28109
rect 633 28106 667 28109
rect 667 28106 701 28109
rect 701 28106 735 28109
rect 735 28106 769 28109
rect 769 28106 803 28109
rect 803 28106 837 28109
rect 837 28106 871 28109
rect 871 28106 905 28109
rect 905 28106 939 28109
rect 939 28106 973 28109
rect 973 28106 1007 28109
rect 1007 28106 1012 28109
rect -996 27932 -458 28106
rect 474 27932 1012 28106
rect -996 27931 -965 27932
rect -965 27931 -931 27932
rect -931 27931 -897 27932
rect -897 27931 -863 27932
rect -863 27931 -829 27932
rect -829 27931 -795 27932
rect -795 27931 -761 27932
rect -761 27931 -727 27932
rect -727 27931 -693 27932
rect -693 27931 -659 27932
rect -659 27931 -625 27932
rect -625 27931 -591 27932
rect -591 27931 -557 27932
rect -557 27931 -523 27932
rect -523 27931 -489 27932
rect -489 27931 -458 27932
rect 474 27931 497 27932
rect 497 27931 531 27932
rect 531 27931 565 27932
rect 565 27931 599 27932
rect 599 27931 633 27932
rect 633 27931 667 27932
rect 667 27931 701 27932
rect 701 27931 735 27932
rect 735 27931 769 27932
rect 769 27931 803 27932
rect 803 27931 837 27932
rect 837 27931 871 27932
rect 871 27931 905 27932
rect 905 27931 939 27932
rect 939 27931 973 27932
rect 973 27931 1007 27932
rect 1007 27931 1012 27932
rect -1593 27796 -1559 27830
rect -1435 27796 -1401 27830
rect -1277 27796 -1243 27830
rect -1119 27796 -1085 27830
rect -961 27796 -927 27830
rect -803 27796 -769 27830
rect -645 27796 -611 27830
rect -487 27796 -453 27830
rect -329 27796 -295 27830
rect -171 27796 -137 27830
rect -13 27796 21 27830
rect 145 27796 179 27830
rect 303 27796 337 27830
rect 461 27796 495 27830
rect 619 27796 653 27830
rect 777 27796 811 27830
rect 935 27796 969 27830
rect 1093 27796 1127 27830
rect 1251 27796 1285 27830
rect 1409 27796 1443 27830
rect 1567 27796 1601 27830
rect -1672 27708 -1638 27734
rect -1672 27700 -1638 27708
rect -1672 27640 -1638 27662
rect -1672 27628 -1638 27640
rect -1672 27572 -1638 27590
rect -1672 27556 -1638 27572
rect -1672 27504 -1638 27518
rect -1672 27484 -1638 27504
rect -1672 27436 -1638 27446
rect -1672 27412 -1638 27436
rect -1672 27368 -1638 27374
rect -1672 27340 -1638 27368
rect -1672 27300 -1638 27302
rect -1672 27268 -1638 27300
rect -1672 27198 -1638 27230
rect -1672 27196 -1638 27198
rect -1672 27130 -1638 27158
rect -1672 27124 -1638 27130
rect -1672 27062 -1638 27086
rect -1672 27052 -1638 27062
rect -1672 26994 -1638 27014
rect -1672 26980 -1638 26994
rect -1672 26926 -1638 26942
rect -1672 26908 -1638 26926
rect -1672 26858 -1638 26870
rect -1672 26836 -1638 26858
rect -1672 26790 -1638 26798
rect -1672 26764 -1638 26790
rect -1514 27708 -1480 27734
rect -1514 27700 -1480 27708
rect -1514 27640 -1480 27662
rect -1514 27628 -1480 27640
rect -1514 27572 -1480 27590
rect -1514 27556 -1480 27572
rect -1514 27504 -1480 27518
rect -1514 27484 -1480 27504
rect -1514 27436 -1480 27446
rect -1514 27412 -1480 27436
rect -1514 27368 -1480 27374
rect -1514 27340 -1480 27368
rect -1514 27300 -1480 27302
rect -1514 27268 -1480 27300
rect -1514 27198 -1480 27230
rect -1514 27196 -1480 27198
rect -1514 27130 -1480 27158
rect -1514 27124 -1480 27130
rect -1514 27062 -1480 27086
rect -1514 27052 -1480 27062
rect -1514 26994 -1480 27014
rect -1514 26980 -1480 26994
rect -1514 26926 -1480 26942
rect -1514 26908 -1480 26926
rect -1514 26858 -1480 26870
rect -1514 26836 -1480 26858
rect -1514 26790 -1480 26798
rect -1514 26764 -1480 26790
rect -1356 27708 -1322 27734
rect -1356 27700 -1322 27708
rect -1356 27640 -1322 27662
rect -1356 27628 -1322 27640
rect -1356 27572 -1322 27590
rect -1356 27556 -1322 27572
rect -1356 27504 -1322 27518
rect -1356 27484 -1322 27504
rect -1356 27436 -1322 27446
rect -1356 27412 -1322 27436
rect -1356 27368 -1322 27374
rect -1356 27340 -1322 27368
rect -1356 27300 -1322 27302
rect -1356 27268 -1322 27300
rect -1356 27198 -1322 27230
rect -1356 27196 -1322 27198
rect -1356 27130 -1322 27158
rect -1356 27124 -1322 27130
rect -1356 27062 -1322 27086
rect -1356 27052 -1322 27062
rect -1356 26994 -1322 27014
rect -1356 26980 -1322 26994
rect -1356 26926 -1322 26942
rect -1356 26908 -1322 26926
rect -1356 26858 -1322 26870
rect -1356 26836 -1322 26858
rect -1356 26790 -1322 26798
rect -1356 26764 -1322 26790
rect -1198 27708 -1164 27734
rect -1198 27700 -1164 27708
rect -1198 27640 -1164 27662
rect -1198 27628 -1164 27640
rect -1198 27572 -1164 27590
rect -1198 27556 -1164 27572
rect -1198 27504 -1164 27518
rect -1198 27484 -1164 27504
rect -1198 27436 -1164 27446
rect -1198 27412 -1164 27436
rect -1198 27368 -1164 27374
rect -1198 27340 -1164 27368
rect -1198 27300 -1164 27302
rect -1198 27268 -1164 27300
rect -1198 27198 -1164 27230
rect -1198 27196 -1164 27198
rect -1198 27130 -1164 27158
rect -1198 27124 -1164 27130
rect -1198 27062 -1164 27086
rect -1198 27052 -1164 27062
rect -1198 26994 -1164 27014
rect -1198 26980 -1164 26994
rect -1198 26926 -1164 26942
rect -1198 26908 -1164 26926
rect -1198 26858 -1164 26870
rect -1198 26836 -1164 26858
rect -1198 26790 -1164 26798
rect -1198 26764 -1164 26790
rect -1040 27708 -1006 27734
rect -1040 27700 -1006 27708
rect -1040 27640 -1006 27662
rect -1040 27628 -1006 27640
rect -1040 27572 -1006 27590
rect -1040 27556 -1006 27572
rect -1040 27504 -1006 27518
rect -1040 27484 -1006 27504
rect -1040 27436 -1006 27446
rect -1040 27412 -1006 27436
rect -1040 27368 -1006 27374
rect -1040 27340 -1006 27368
rect -1040 27300 -1006 27302
rect -1040 27268 -1006 27300
rect -1040 27198 -1006 27230
rect -1040 27196 -1006 27198
rect -1040 27130 -1006 27158
rect -1040 27124 -1006 27130
rect -1040 27062 -1006 27086
rect -1040 27052 -1006 27062
rect -1040 26994 -1006 27014
rect -1040 26980 -1006 26994
rect -1040 26926 -1006 26942
rect -1040 26908 -1006 26926
rect -1040 26858 -1006 26870
rect -1040 26836 -1006 26858
rect -1040 26790 -1006 26798
rect -1040 26764 -1006 26790
rect -882 27708 -848 27734
rect -882 27700 -848 27708
rect -882 27640 -848 27662
rect -882 27628 -848 27640
rect -882 27572 -848 27590
rect -882 27556 -848 27572
rect -882 27504 -848 27518
rect -882 27484 -848 27504
rect -882 27436 -848 27446
rect -882 27412 -848 27436
rect -882 27368 -848 27374
rect -882 27340 -848 27368
rect -882 27300 -848 27302
rect -882 27268 -848 27300
rect -882 27198 -848 27230
rect -882 27196 -848 27198
rect -882 27130 -848 27158
rect -882 27124 -848 27130
rect -882 27062 -848 27086
rect -882 27052 -848 27062
rect -882 26994 -848 27014
rect -882 26980 -848 26994
rect -882 26926 -848 26942
rect -882 26908 -848 26926
rect -882 26858 -848 26870
rect -882 26836 -848 26858
rect -882 26790 -848 26798
rect -882 26764 -848 26790
rect -724 27708 -690 27734
rect -724 27700 -690 27708
rect -724 27640 -690 27662
rect -724 27628 -690 27640
rect -724 27572 -690 27590
rect -724 27556 -690 27572
rect -724 27504 -690 27518
rect -724 27484 -690 27504
rect -724 27436 -690 27446
rect -724 27412 -690 27436
rect -724 27368 -690 27374
rect -724 27340 -690 27368
rect -724 27300 -690 27302
rect -724 27268 -690 27300
rect -724 27198 -690 27230
rect -724 27196 -690 27198
rect -724 27130 -690 27158
rect -724 27124 -690 27130
rect -724 27062 -690 27086
rect -724 27052 -690 27062
rect -724 26994 -690 27014
rect -724 26980 -690 26994
rect -724 26926 -690 26942
rect -724 26908 -690 26926
rect -724 26858 -690 26870
rect -724 26836 -690 26858
rect -724 26790 -690 26798
rect -724 26764 -690 26790
rect -566 27708 -532 27734
rect -566 27700 -532 27708
rect -566 27640 -532 27662
rect -566 27628 -532 27640
rect -566 27572 -532 27590
rect -566 27556 -532 27572
rect -566 27504 -532 27518
rect -566 27484 -532 27504
rect -566 27436 -532 27446
rect -566 27412 -532 27436
rect -566 27368 -532 27374
rect -566 27340 -532 27368
rect -566 27300 -532 27302
rect -566 27268 -532 27300
rect -566 27198 -532 27230
rect -566 27196 -532 27198
rect -566 27130 -532 27158
rect -566 27124 -532 27130
rect -566 27062 -532 27086
rect -566 27052 -532 27062
rect -566 26994 -532 27014
rect -566 26980 -532 26994
rect -566 26926 -532 26942
rect -566 26908 -532 26926
rect -566 26858 -532 26870
rect -566 26836 -532 26858
rect -566 26790 -532 26798
rect -566 26764 -532 26790
rect -408 27708 -374 27734
rect -408 27700 -374 27708
rect -408 27640 -374 27662
rect -408 27628 -374 27640
rect -408 27572 -374 27590
rect -408 27556 -374 27572
rect -408 27504 -374 27518
rect -408 27484 -374 27504
rect -408 27436 -374 27446
rect -408 27412 -374 27436
rect -408 27368 -374 27374
rect -408 27340 -374 27368
rect -408 27300 -374 27302
rect -408 27268 -374 27300
rect -408 27198 -374 27230
rect -408 27196 -374 27198
rect -408 27130 -374 27158
rect -408 27124 -374 27130
rect -408 27062 -374 27086
rect -408 27052 -374 27062
rect -408 26994 -374 27014
rect -408 26980 -374 26994
rect -408 26926 -374 26942
rect -408 26908 -374 26926
rect -408 26858 -374 26870
rect -408 26836 -374 26858
rect -408 26790 -374 26798
rect -408 26764 -374 26790
rect -250 27708 -216 27734
rect -250 27700 -216 27708
rect -250 27640 -216 27662
rect -250 27628 -216 27640
rect -250 27572 -216 27590
rect -250 27556 -216 27572
rect -250 27504 -216 27518
rect -250 27484 -216 27504
rect -250 27436 -216 27446
rect -250 27412 -216 27436
rect -250 27368 -216 27374
rect -250 27340 -216 27368
rect -250 27300 -216 27302
rect -250 27268 -216 27300
rect -250 27198 -216 27230
rect -250 27196 -216 27198
rect -250 27130 -216 27158
rect -250 27124 -216 27130
rect -250 27062 -216 27086
rect -250 27052 -216 27062
rect -250 26994 -216 27014
rect -250 26980 -216 26994
rect -250 26926 -216 26942
rect -250 26908 -216 26926
rect -250 26858 -216 26870
rect -250 26836 -216 26858
rect -250 26790 -216 26798
rect -250 26764 -216 26790
rect -92 27708 -58 27734
rect -92 27700 -58 27708
rect -92 27640 -58 27662
rect -92 27628 -58 27640
rect -92 27572 -58 27590
rect -92 27556 -58 27572
rect -92 27504 -58 27518
rect -92 27484 -58 27504
rect -92 27436 -58 27446
rect -92 27412 -58 27436
rect -92 27368 -58 27374
rect -92 27340 -58 27368
rect -92 27300 -58 27302
rect -92 27268 -58 27300
rect -92 27198 -58 27230
rect -92 27196 -58 27198
rect -92 27130 -58 27158
rect -92 27124 -58 27130
rect -92 27062 -58 27086
rect -92 27052 -58 27062
rect -92 26994 -58 27014
rect -92 26980 -58 26994
rect -92 26926 -58 26942
rect -92 26908 -58 26926
rect -92 26858 -58 26870
rect -92 26836 -58 26858
rect -92 26790 -58 26798
rect -92 26764 -58 26790
rect 66 27708 100 27734
rect 66 27700 100 27708
rect 66 27640 100 27662
rect 66 27628 100 27640
rect 66 27572 100 27590
rect 66 27556 100 27572
rect 66 27504 100 27518
rect 66 27484 100 27504
rect 66 27436 100 27446
rect 66 27412 100 27436
rect 66 27368 100 27374
rect 66 27340 100 27368
rect 66 27300 100 27302
rect 66 27268 100 27300
rect 66 27198 100 27230
rect 66 27196 100 27198
rect 66 27130 100 27158
rect 66 27124 100 27130
rect 66 27062 100 27086
rect 66 27052 100 27062
rect 66 26994 100 27014
rect 66 26980 100 26994
rect 66 26926 100 26942
rect 66 26908 100 26926
rect 66 26858 100 26870
rect 66 26836 100 26858
rect 66 26790 100 26798
rect 66 26764 100 26790
rect 224 27708 258 27734
rect 224 27700 258 27708
rect 224 27640 258 27662
rect 224 27628 258 27640
rect 224 27572 258 27590
rect 224 27556 258 27572
rect 224 27504 258 27518
rect 224 27484 258 27504
rect 224 27436 258 27446
rect 224 27412 258 27436
rect 224 27368 258 27374
rect 224 27340 258 27368
rect 224 27300 258 27302
rect 224 27268 258 27300
rect 224 27198 258 27230
rect 224 27196 258 27198
rect 224 27130 258 27158
rect 224 27124 258 27130
rect 224 27062 258 27086
rect 224 27052 258 27062
rect 224 26994 258 27014
rect 224 26980 258 26994
rect 224 26926 258 26942
rect 224 26908 258 26926
rect 224 26858 258 26870
rect 224 26836 258 26858
rect 224 26790 258 26798
rect 224 26764 258 26790
rect 382 27708 416 27734
rect 382 27700 416 27708
rect 382 27640 416 27662
rect 382 27628 416 27640
rect 382 27572 416 27590
rect 382 27556 416 27572
rect 382 27504 416 27518
rect 382 27484 416 27504
rect 382 27436 416 27446
rect 382 27412 416 27436
rect 382 27368 416 27374
rect 382 27340 416 27368
rect 382 27300 416 27302
rect 382 27268 416 27300
rect 382 27198 416 27230
rect 382 27196 416 27198
rect 382 27130 416 27158
rect 382 27124 416 27130
rect 382 27062 416 27086
rect 382 27052 416 27062
rect 382 26994 416 27014
rect 382 26980 416 26994
rect 382 26926 416 26942
rect 382 26908 416 26926
rect 382 26858 416 26870
rect 382 26836 416 26858
rect 382 26790 416 26798
rect 382 26764 416 26790
rect 540 27708 574 27734
rect 540 27700 574 27708
rect 540 27640 574 27662
rect 540 27628 574 27640
rect 540 27572 574 27590
rect 540 27556 574 27572
rect 540 27504 574 27518
rect 540 27484 574 27504
rect 540 27436 574 27446
rect 540 27412 574 27436
rect 540 27368 574 27374
rect 540 27340 574 27368
rect 540 27300 574 27302
rect 540 27268 574 27300
rect 540 27198 574 27230
rect 540 27196 574 27198
rect 540 27130 574 27158
rect 540 27124 574 27130
rect 540 27062 574 27086
rect 540 27052 574 27062
rect 540 26994 574 27014
rect 540 26980 574 26994
rect 540 26926 574 26942
rect 540 26908 574 26926
rect 540 26858 574 26870
rect 540 26836 574 26858
rect 540 26790 574 26798
rect 540 26764 574 26790
rect 698 27708 732 27734
rect 698 27700 732 27708
rect 698 27640 732 27662
rect 698 27628 732 27640
rect 698 27572 732 27590
rect 698 27556 732 27572
rect 698 27504 732 27518
rect 698 27484 732 27504
rect 698 27436 732 27446
rect 698 27412 732 27436
rect 698 27368 732 27374
rect 698 27340 732 27368
rect 698 27300 732 27302
rect 698 27268 732 27300
rect 698 27198 732 27230
rect 698 27196 732 27198
rect 698 27130 732 27158
rect 698 27124 732 27130
rect 698 27062 732 27086
rect 698 27052 732 27062
rect 698 26994 732 27014
rect 698 26980 732 26994
rect 698 26926 732 26942
rect 698 26908 732 26926
rect 698 26858 732 26870
rect 698 26836 732 26858
rect 698 26790 732 26798
rect 698 26764 732 26790
rect 856 27708 890 27734
rect 856 27700 890 27708
rect 856 27640 890 27662
rect 856 27628 890 27640
rect 856 27572 890 27590
rect 856 27556 890 27572
rect 856 27504 890 27518
rect 856 27484 890 27504
rect 856 27436 890 27446
rect 856 27412 890 27436
rect 856 27368 890 27374
rect 856 27340 890 27368
rect 856 27300 890 27302
rect 856 27268 890 27300
rect 856 27198 890 27230
rect 856 27196 890 27198
rect 856 27130 890 27158
rect 856 27124 890 27130
rect 856 27062 890 27086
rect 856 27052 890 27062
rect 856 26994 890 27014
rect 856 26980 890 26994
rect 856 26926 890 26942
rect 856 26908 890 26926
rect 856 26858 890 26870
rect 856 26836 890 26858
rect 856 26790 890 26798
rect 856 26764 890 26790
rect 1014 27708 1048 27734
rect 1014 27700 1048 27708
rect 1014 27640 1048 27662
rect 1014 27628 1048 27640
rect 1014 27572 1048 27590
rect 1014 27556 1048 27572
rect 1014 27504 1048 27518
rect 1014 27484 1048 27504
rect 1014 27436 1048 27446
rect 1014 27412 1048 27436
rect 1014 27368 1048 27374
rect 1014 27340 1048 27368
rect 1014 27300 1048 27302
rect 1014 27268 1048 27300
rect 1014 27198 1048 27230
rect 1014 27196 1048 27198
rect 1014 27130 1048 27158
rect 1014 27124 1048 27130
rect 1014 27062 1048 27086
rect 1014 27052 1048 27062
rect 1014 26994 1048 27014
rect 1014 26980 1048 26994
rect 1014 26926 1048 26942
rect 1014 26908 1048 26926
rect 1014 26858 1048 26870
rect 1014 26836 1048 26858
rect 1014 26790 1048 26798
rect 1014 26764 1048 26790
rect 1172 27708 1206 27734
rect 1172 27700 1206 27708
rect 1172 27640 1206 27662
rect 1172 27628 1206 27640
rect 1172 27572 1206 27590
rect 1172 27556 1206 27572
rect 1172 27504 1206 27518
rect 1172 27484 1206 27504
rect 1172 27436 1206 27446
rect 1172 27412 1206 27436
rect 1172 27368 1206 27374
rect 1172 27340 1206 27368
rect 1172 27300 1206 27302
rect 1172 27268 1206 27300
rect 1172 27198 1206 27230
rect 1172 27196 1206 27198
rect 1172 27130 1206 27158
rect 1172 27124 1206 27130
rect 1172 27062 1206 27086
rect 1172 27052 1206 27062
rect 1172 26994 1206 27014
rect 1172 26980 1206 26994
rect 1172 26926 1206 26942
rect 1172 26908 1206 26926
rect 1172 26858 1206 26870
rect 1172 26836 1206 26858
rect 1172 26790 1206 26798
rect 1172 26764 1206 26790
rect 1330 27708 1364 27734
rect 1330 27700 1364 27708
rect 1330 27640 1364 27662
rect 1330 27628 1364 27640
rect 1330 27572 1364 27590
rect 1330 27556 1364 27572
rect 1330 27504 1364 27518
rect 1330 27484 1364 27504
rect 1330 27436 1364 27446
rect 1330 27412 1364 27436
rect 1330 27368 1364 27374
rect 1330 27340 1364 27368
rect 1330 27300 1364 27302
rect 1330 27268 1364 27300
rect 1330 27198 1364 27230
rect 1330 27196 1364 27198
rect 1330 27130 1364 27158
rect 1330 27124 1364 27130
rect 1330 27062 1364 27086
rect 1330 27052 1364 27062
rect 1330 26994 1364 27014
rect 1330 26980 1364 26994
rect 1330 26926 1364 26942
rect 1330 26908 1364 26926
rect 1330 26858 1364 26870
rect 1330 26836 1364 26858
rect 1330 26790 1364 26798
rect 1330 26764 1364 26790
rect 1488 27708 1522 27734
rect 1488 27700 1522 27708
rect 1488 27640 1522 27662
rect 1488 27628 1522 27640
rect 1488 27572 1522 27590
rect 1488 27556 1522 27572
rect 1488 27504 1522 27518
rect 1488 27484 1522 27504
rect 1488 27436 1522 27446
rect 1488 27412 1522 27436
rect 1488 27368 1522 27374
rect 1488 27340 1522 27368
rect 1488 27300 1522 27302
rect 1488 27268 1522 27300
rect 1488 27198 1522 27230
rect 1488 27196 1522 27198
rect 1488 27130 1522 27158
rect 1488 27124 1522 27130
rect 1488 27062 1522 27086
rect 1488 27052 1522 27062
rect 1488 26994 1522 27014
rect 1488 26980 1522 26994
rect 1488 26926 1522 26942
rect 1488 26908 1522 26926
rect 1488 26858 1522 26870
rect 1488 26836 1522 26858
rect 1488 26790 1522 26798
rect 1488 26764 1522 26790
rect 1646 27708 1680 27734
rect 1646 27700 1680 27708
rect 1646 27640 1680 27662
rect 1646 27628 1680 27640
rect 1646 27572 1680 27590
rect 1646 27556 1680 27572
rect 1646 27504 1680 27518
rect 1646 27484 1680 27504
rect 1646 27436 1680 27446
rect 1646 27412 1680 27436
rect 1646 27368 1680 27374
rect 1646 27340 1680 27368
rect 1646 27300 1680 27302
rect 1646 27268 1680 27300
rect 1646 27198 1680 27230
rect 1646 27196 1680 27198
rect 1646 27130 1680 27158
rect 1646 27124 1680 27130
rect 1646 27062 1680 27086
rect 1646 27052 1680 27062
rect 1646 26994 1680 27014
rect 1646 26980 1680 26994
rect 1646 26926 1680 26942
rect 1646 26908 1680 26926
rect 1646 26858 1680 26870
rect 1646 26836 1680 26858
rect 1646 26790 1680 26798
rect 1646 26764 1680 26790
rect -1593 26668 -1559 26702
rect -1435 26668 -1401 26702
rect -1277 26668 -1243 26702
rect -1119 26668 -1085 26702
rect -961 26668 -927 26702
rect -803 26668 -769 26702
rect -645 26668 -611 26702
rect -487 26668 -453 26702
rect -329 26668 -295 26702
rect -171 26668 -137 26702
rect -13 26668 21 26702
rect 145 26668 179 26702
rect 303 26668 337 26702
rect 461 26668 495 26702
rect 619 26668 653 26702
rect 777 26668 811 26702
rect 935 26668 969 26702
rect 1093 26668 1127 26702
rect 1251 26668 1285 26702
rect 1409 26668 1443 26702
rect 1567 26668 1601 26702
rect -306 26321 -290 26355
rect -290 26321 -272 26355
rect -234 26321 -222 26355
rect -222 26321 -200 26355
rect -162 26321 -154 26355
rect -154 26321 -128 26355
rect -90 26321 -86 26355
rect -86 26321 -56 26355
rect -18 26321 16 26355
rect 54 26321 84 26355
rect 84 26321 88 26355
rect 126 26321 152 26355
rect 152 26321 160 26355
rect 198 26321 220 26355
rect 220 26321 232 26355
rect 270 26321 288 26355
rect 288 26321 304 26355
rect -492 26219 -458 26253
rect -334 26219 -300 26253
rect -176 26219 -142 26253
rect -18 26219 16 26253
rect 140 26219 174 26253
rect 298 26219 332 26253
rect 456 26219 490 26253
rect -571 26140 -537 26166
rect -571 26132 -537 26140
rect -571 26072 -537 26094
rect -571 26060 -537 26072
rect -571 26004 -537 26022
rect -571 25988 -537 26004
rect -571 25936 -537 25950
rect -571 25916 -537 25936
rect -571 25868 -537 25878
rect -571 25844 -537 25868
rect -571 25800 -537 25806
rect -571 25772 -537 25800
rect -571 25732 -537 25734
rect -571 25700 -537 25732
rect -571 25630 -537 25662
rect -571 25628 -537 25630
rect -571 25562 -537 25590
rect -571 25556 -537 25562
rect -571 25494 -537 25518
rect -571 25484 -537 25494
rect -571 25426 -537 25446
rect -571 25412 -537 25426
rect -571 25358 -537 25374
rect -571 25340 -537 25358
rect -571 25290 -537 25302
rect -571 25268 -537 25290
rect -571 25222 -537 25230
rect -571 25196 -537 25222
rect -413 26140 -379 26166
rect -413 26132 -379 26140
rect -413 26072 -379 26094
rect -413 26060 -379 26072
rect -413 26004 -379 26022
rect -413 25988 -379 26004
rect -413 25936 -379 25950
rect -413 25916 -379 25936
rect -413 25868 -379 25878
rect -413 25844 -379 25868
rect -413 25800 -379 25806
rect -413 25772 -379 25800
rect -413 25732 -379 25734
rect -413 25700 -379 25732
rect -413 25630 -379 25662
rect -413 25628 -379 25630
rect -413 25562 -379 25590
rect -413 25556 -379 25562
rect -413 25494 -379 25518
rect -413 25484 -379 25494
rect -413 25426 -379 25446
rect -413 25412 -379 25426
rect -413 25358 -379 25374
rect -413 25340 -379 25358
rect -413 25290 -379 25302
rect -413 25268 -379 25290
rect -413 25222 -379 25230
rect -413 25196 -379 25222
rect -255 26140 -221 26166
rect -255 26132 -221 26140
rect -255 26072 -221 26094
rect -255 26060 -221 26072
rect -255 26004 -221 26022
rect -255 25988 -221 26004
rect -255 25936 -221 25950
rect -255 25916 -221 25936
rect -255 25868 -221 25878
rect -255 25844 -221 25868
rect -255 25800 -221 25806
rect -255 25772 -221 25800
rect -255 25732 -221 25734
rect -255 25700 -221 25732
rect -255 25630 -221 25662
rect -255 25628 -221 25630
rect -255 25562 -221 25590
rect -255 25556 -221 25562
rect -255 25494 -221 25518
rect -255 25484 -221 25494
rect -255 25426 -221 25446
rect -255 25412 -221 25426
rect -255 25358 -221 25374
rect -255 25340 -221 25358
rect -255 25290 -221 25302
rect -255 25268 -221 25290
rect -255 25222 -221 25230
rect -255 25196 -221 25222
rect -97 26140 -63 26166
rect -97 26132 -63 26140
rect -97 26072 -63 26094
rect -97 26060 -63 26072
rect -97 26004 -63 26022
rect -97 25988 -63 26004
rect -97 25936 -63 25950
rect -97 25916 -63 25936
rect -97 25868 -63 25878
rect -97 25844 -63 25868
rect -97 25800 -63 25806
rect -97 25772 -63 25800
rect -97 25732 -63 25734
rect -97 25700 -63 25732
rect -97 25630 -63 25662
rect -97 25628 -63 25630
rect -97 25562 -63 25590
rect -97 25556 -63 25562
rect -97 25494 -63 25518
rect -97 25484 -63 25494
rect -97 25426 -63 25446
rect -97 25412 -63 25426
rect -97 25358 -63 25374
rect -97 25340 -63 25358
rect -97 25290 -63 25302
rect -97 25268 -63 25290
rect -97 25222 -63 25230
rect -97 25196 -63 25222
rect 61 26140 95 26166
rect 61 26132 95 26140
rect 61 26072 95 26094
rect 61 26060 95 26072
rect 61 26004 95 26022
rect 61 25988 95 26004
rect 61 25936 95 25950
rect 61 25916 95 25936
rect 61 25868 95 25878
rect 61 25844 95 25868
rect 61 25800 95 25806
rect 61 25772 95 25800
rect 61 25732 95 25734
rect 61 25700 95 25732
rect 61 25630 95 25662
rect 61 25628 95 25630
rect 61 25562 95 25590
rect 61 25556 95 25562
rect 61 25494 95 25518
rect 61 25484 95 25494
rect 61 25426 95 25446
rect 61 25412 95 25426
rect 61 25358 95 25374
rect 61 25340 95 25358
rect 61 25290 95 25302
rect 61 25268 95 25290
rect 61 25222 95 25230
rect 61 25196 95 25222
rect 219 26140 253 26166
rect 219 26132 253 26140
rect 219 26072 253 26094
rect 219 26060 253 26072
rect 219 26004 253 26022
rect 219 25988 253 26004
rect 219 25936 253 25950
rect 219 25916 253 25936
rect 219 25868 253 25878
rect 219 25844 253 25868
rect 219 25800 253 25806
rect 219 25772 253 25800
rect 219 25732 253 25734
rect 219 25700 253 25732
rect 219 25630 253 25662
rect 219 25628 253 25630
rect 219 25562 253 25590
rect 219 25556 253 25562
rect 219 25494 253 25518
rect 219 25484 253 25494
rect 219 25426 253 25446
rect 219 25412 253 25426
rect 219 25358 253 25374
rect 219 25340 253 25358
rect 219 25290 253 25302
rect 219 25268 253 25290
rect 219 25222 253 25230
rect 219 25196 253 25222
rect 377 26140 411 26166
rect 377 26132 411 26140
rect 377 26072 411 26094
rect 377 26060 411 26072
rect 377 26004 411 26022
rect 377 25988 411 26004
rect 377 25936 411 25950
rect 377 25916 411 25936
rect 377 25868 411 25878
rect 377 25844 411 25868
rect 377 25800 411 25806
rect 377 25772 411 25800
rect 377 25732 411 25734
rect 377 25700 411 25732
rect 377 25630 411 25662
rect 377 25628 411 25630
rect 377 25562 411 25590
rect 377 25556 411 25562
rect 377 25494 411 25518
rect 377 25484 411 25494
rect 377 25426 411 25446
rect 377 25412 411 25426
rect 377 25358 411 25374
rect 377 25340 411 25358
rect 377 25290 411 25302
rect 377 25268 411 25290
rect 377 25222 411 25230
rect 377 25196 411 25222
rect 535 26140 569 26166
rect 535 26132 569 26140
rect 535 26072 569 26094
rect 535 26060 569 26072
rect 535 26004 569 26022
rect 535 25988 569 26004
rect 535 25936 569 25950
rect 535 25916 569 25936
rect 535 25868 569 25878
rect 535 25844 569 25868
rect 535 25800 569 25806
rect 535 25772 569 25800
rect 535 25732 569 25734
rect 535 25700 569 25732
rect 535 25630 569 25662
rect 535 25628 569 25630
rect 535 25562 569 25590
rect 535 25556 569 25562
rect 535 25494 569 25518
rect 535 25484 569 25494
rect 535 25426 569 25446
rect 535 25412 569 25426
rect 535 25358 569 25374
rect 535 25340 569 25358
rect 535 25290 569 25302
rect 535 25268 569 25290
rect 535 25222 569 25230
rect 535 25196 569 25222
rect -492 25109 -458 25143
rect -334 25109 -300 25143
rect -176 25109 -142 25143
rect -18 25109 16 25143
rect 140 25109 174 25143
rect 298 25109 332 25143
rect 456 25109 490 25143
rect -306 25007 -290 25041
rect -290 25007 -272 25041
rect -234 25007 -222 25041
rect -222 25007 -200 25041
rect -162 25007 -154 25041
rect -154 25007 -128 25041
rect -90 25007 -86 25041
rect -86 25007 -56 25041
rect -18 25007 16 25041
rect 54 25007 84 25041
rect 84 25007 88 25041
rect 126 25007 152 25041
rect 152 25007 160 25041
rect 198 25007 220 25041
rect 220 25007 232 25041
rect 270 25007 288 25041
rect 288 25007 304 25041
rect -306 24801 -290 24835
rect -290 24801 -272 24835
rect -234 24801 -222 24835
rect -222 24801 -200 24835
rect -162 24801 -154 24835
rect -154 24801 -128 24835
rect -90 24801 -86 24835
rect -86 24801 -56 24835
rect -18 24801 16 24835
rect 54 24801 84 24835
rect 84 24801 88 24835
rect 126 24801 152 24835
rect 152 24801 160 24835
rect 198 24801 220 24835
rect 220 24801 232 24835
rect 270 24801 288 24835
rect 288 24801 304 24835
rect -492 24699 -458 24733
rect -334 24699 -300 24733
rect -176 24699 -142 24733
rect -18 24699 16 24733
rect 140 24699 174 24733
rect 298 24699 332 24733
rect 456 24699 490 24733
rect -571 24620 -537 24646
rect -571 24612 -537 24620
rect -571 24552 -537 24574
rect -571 24540 -537 24552
rect -571 24484 -537 24502
rect -571 24468 -537 24484
rect -571 24416 -537 24430
rect -571 24396 -537 24416
rect -571 24348 -537 24358
rect -571 24324 -537 24348
rect -571 24280 -537 24286
rect -571 24252 -537 24280
rect -571 24212 -537 24214
rect -571 24180 -537 24212
rect -571 24110 -537 24142
rect -571 24108 -537 24110
rect -571 24042 -537 24070
rect -571 24036 -537 24042
rect -571 23974 -537 23998
rect -571 23964 -537 23974
rect -571 23906 -537 23926
rect -571 23892 -537 23906
rect -571 23838 -537 23854
rect -571 23820 -537 23838
rect -571 23770 -537 23782
rect -571 23748 -537 23770
rect -571 23702 -537 23710
rect -571 23676 -537 23702
rect -413 24620 -379 24646
rect -413 24612 -379 24620
rect -413 24552 -379 24574
rect -413 24540 -379 24552
rect -413 24484 -379 24502
rect -413 24468 -379 24484
rect -413 24416 -379 24430
rect -413 24396 -379 24416
rect -413 24348 -379 24358
rect -413 24324 -379 24348
rect -413 24280 -379 24286
rect -413 24252 -379 24280
rect -413 24212 -379 24214
rect -413 24180 -379 24212
rect -413 24110 -379 24142
rect -413 24108 -379 24110
rect -413 24042 -379 24070
rect -413 24036 -379 24042
rect -413 23974 -379 23998
rect -413 23964 -379 23974
rect -413 23906 -379 23926
rect -413 23892 -379 23906
rect -413 23838 -379 23854
rect -413 23820 -379 23838
rect -413 23770 -379 23782
rect -413 23748 -379 23770
rect -413 23702 -379 23710
rect -413 23676 -379 23702
rect -255 24620 -221 24646
rect -255 24612 -221 24620
rect -255 24552 -221 24574
rect -255 24540 -221 24552
rect -255 24484 -221 24502
rect -255 24468 -221 24484
rect -255 24416 -221 24430
rect -255 24396 -221 24416
rect -255 24348 -221 24358
rect -255 24324 -221 24348
rect -255 24280 -221 24286
rect -255 24252 -221 24280
rect -255 24212 -221 24214
rect -255 24180 -221 24212
rect -255 24110 -221 24142
rect -255 24108 -221 24110
rect -255 24042 -221 24070
rect -255 24036 -221 24042
rect -255 23974 -221 23998
rect -255 23964 -221 23974
rect -255 23906 -221 23926
rect -255 23892 -221 23906
rect -255 23838 -221 23854
rect -255 23820 -221 23838
rect -255 23770 -221 23782
rect -255 23748 -221 23770
rect -255 23702 -221 23710
rect -255 23676 -221 23702
rect -97 24620 -63 24646
rect -97 24612 -63 24620
rect -97 24552 -63 24574
rect -97 24540 -63 24552
rect -97 24484 -63 24502
rect -97 24468 -63 24484
rect -97 24416 -63 24430
rect -97 24396 -63 24416
rect -97 24348 -63 24358
rect -97 24324 -63 24348
rect -97 24280 -63 24286
rect -97 24252 -63 24280
rect -97 24212 -63 24214
rect -97 24180 -63 24212
rect -97 24110 -63 24142
rect -97 24108 -63 24110
rect -97 24042 -63 24070
rect -97 24036 -63 24042
rect -97 23974 -63 23998
rect -97 23964 -63 23974
rect -97 23906 -63 23926
rect -97 23892 -63 23906
rect -97 23838 -63 23854
rect -97 23820 -63 23838
rect -97 23770 -63 23782
rect -97 23748 -63 23770
rect -97 23702 -63 23710
rect -97 23676 -63 23702
rect 61 24620 95 24646
rect 61 24612 95 24620
rect 61 24552 95 24574
rect 61 24540 95 24552
rect 61 24484 95 24502
rect 61 24468 95 24484
rect 61 24416 95 24430
rect 61 24396 95 24416
rect 61 24348 95 24358
rect 61 24324 95 24348
rect 61 24280 95 24286
rect 61 24252 95 24280
rect 61 24212 95 24214
rect 61 24180 95 24212
rect 61 24110 95 24142
rect 61 24108 95 24110
rect 61 24042 95 24070
rect 61 24036 95 24042
rect 61 23974 95 23998
rect 61 23964 95 23974
rect 61 23906 95 23926
rect 61 23892 95 23906
rect 61 23838 95 23854
rect 61 23820 95 23838
rect 61 23770 95 23782
rect 61 23748 95 23770
rect 61 23702 95 23710
rect 61 23676 95 23702
rect 219 24620 253 24646
rect 219 24612 253 24620
rect 219 24552 253 24574
rect 219 24540 253 24552
rect 219 24484 253 24502
rect 219 24468 253 24484
rect 219 24416 253 24430
rect 219 24396 253 24416
rect 219 24348 253 24358
rect 219 24324 253 24348
rect 219 24280 253 24286
rect 219 24252 253 24280
rect 219 24212 253 24214
rect 219 24180 253 24212
rect 219 24110 253 24142
rect 219 24108 253 24110
rect 219 24042 253 24070
rect 219 24036 253 24042
rect 219 23974 253 23998
rect 219 23964 253 23974
rect 219 23906 253 23926
rect 219 23892 253 23906
rect 219 23838 253 23854
rect 219 23820 253 23838
rect 219 23770 253 23782
rect 219 23748 253 23770
rect 219 23702 253 23710
rect 219 23676 253 23702
rect 377 24620 411 24646
rect 377 24612 411 24620
rect 377 24552 411 24574
rect 377 24540 411 24552
rect 377 24484 411 24502
rect 377 24468 411 24484
rect 377 24416 411 24430
rect 377 24396 411 24416
rect 377 24348 411 24358
rect 377 24324 411 24348
rect 377 24280 411 24286
rect 377 24252 411 24280
rect 377 24212 411 24214
rect 377 24180 411 24212
rect 377 24110 411 24142
rect 377 24108 411 24110
rect 377 24042 411 24070
rect 377 24036 411 24042
rect 377 23974 411 23998
rect 377 23964 411 23974
rect 377 23906 411 23926
rect 377 23892 411 23906
rect 377 23838 411 23854
rect 377 23820 411 23838
rect 377 23770 411 23782
rect 377 23748 411 23770
rect 377 23702 411 23710
rect 377 23676 411 23702
rect 535 24620 569 24646
rect 535 24612 569 24620
rect 535 24552 569 24574
rect 535 24540 569 24552
rect 535 24484 569 24502
rect 535 24468 569 24484
rect 535 24416 569 24430
rect 535 24396 569 24416
rect 535 24348 569 24358
rect 535 24324 569 24348
rect 535 24280 569 24286
rect 535 24252 569 24280
rect 535 24212 569 24214
rect 535 24180 569 24212
rect 535 24110 569 24142
rect 535 24108 569 24110
rect 535 24042 569 24070
rect 535 24036 569 24042
rect 535 23974 569 23998
rect 535 23964 569 23974
rect 535 23906 569 23926
rect 535 23892 569 23906
rect 535 23838 569 23854
rect 535 23820 569 23838
rect 535 23770 569 23782
rect 535 23748 569 23770
rect 535 23702 569 23710
rect 535 23676 569 23702
rect -492 23589 -458 23623
rect -334 23589 -300 23623
rect -176 23589 -142 23623
rect -18 23589 16 23623
rect 140 23589 174 23623
rect 298 23589 332 23623
rect 456 23589 490 23623
rect -306 23487 -290 23521
rect -290 23487 -272 23521
rect -234 23487 -222 23521
rect -222 23487 -200 23521
rect -162 23487 -154 23521
rect -154 23487 -128 23521
rect -90 23487 -86 23521
rect -86 23487 -56 23521
rect -18 23487 16 23521
rect 54 23487 84 23521
rect 84 23487 88 23521
rect 126 23487 152 23521
rect 152 23487 160 23521
rect 198 23487 220 23521
rect 220 23487 232 23521
rect 270 23487 288 23521
rect 288 23487 304 23521
rect -806 23280 -796 23314
rect -796 23280 -772 23314
rect -734 23280 -728 23314
rect -728 23280 -700 23314
rect -662 23280 -660 23314
rect -660 23280 -628 23314
rect -590 23280 -558 23314
rect -558 23280 -556 23314
rect -518 23280 -490 23314
rect -490 23280 -484 23314
rect -446 23280 -422 23314
rect -422 23280 -412 23314
rect -374 23280 -354 23314
rect -354 23280 -340 23314
rect -302 23280 -286 23314
rect -286 23280 -268 23314
rect -230 23280 -218 23314
rect -218 23280 -196 23314
rect -158 23280 -150 23314
rect -150 23280 -124 23314
rect -86 23280 -82 23314
rect -82 23280 -52 23314
rect -14 23280 20 23314
rect 58 23280 88 23314
rect 88 23280 92 23314
rect 130 23280 156 23314
rect 156 23280 164 23314
rect 202 23280 224 23314
rect 224 23280 236 23314
rect 274 23280 292 23314
rect 292 23280 308 23314
rect 346 23280 360 23314
rect 360 23280 380 23314
rect 418 23280 428 23314
rect 428 23280 452 23314
rect 490 23280 496 23314
rect 496 23280 524 23314
rect 562 23280 564 23314
rect 564 23280 596 23314
rect 634 23280 666 23314
rect 666 23280 668 23314
rect 706 23280 734 23314
rect 734 23280 740 23314
rect 778 23280 802 23314
rect 802 23280 812 23314
rect -1469 23178 -1467 23212
rect -1467 23178 -1435 23212
rect -1397 23178 -1365 23212
rect -1365 23178 -1363 23212
rect -1211 23178 -1209 23212
rect -1209 23178 -1177 23212
rect -1139 23178 -1107 23212
rect -1107 23178 -1105 23212
rect -953 23178 -951 23212
rect -951 23178 -919 23212
rect -881 23178 -849 23212
rect -849 23178 -847 23212
rect -695 23178 -693 23212
rect -693 23178 -661 23212
rect -623 23178 -591 23212
rect -591 23178 -589 23212
rect -437 23178 -435 23212
rect -435 23178 -403 23212
rect -365 23178 -333 23212
rect -333 23178 -331 23212
rect -179 23178 -177 23212
rect -177 23178 -145 23212
rect -107 23178 -75 23212
rect -75 23178 -73 23212
rect 79 23178 81 23212
rect 81 23178 113 23212
rect 151 23178 183 23212
rect 183 23178 185 23212
rect 337 23178 339 23212
rect 339 23178 371 23212
rect 409 23178 441 23212
rect 441 23178 443 23212
rect 595 23178 597 23212
rect 597 23178 629 23212
rect 667 23178 699 23212
rect 699 23178 701 23212
rect 853 23178 855 23212
rect 855 23178 887 23212
rect 925 23178 957 23212
rect 957 23178 959 23212
rect 1111 23178 1113 23212
rect 1113 23178 1145 23212
rect 1183 23178 1215 23212
rect 1215 23178 1217 23212
rect 1369 23178 1371 23212
rect 1371 23178 1403 23212
rect 1441 23178 1473 23212
rect 1473 23178 1475 23212
rect -1562 23099 -1528 23125
rect -1562 23091 -1528 23099
rect -1562 23031 -1528 23053
rect -1562 23019 -1528 23031
rect -1562 22963 -1528 22981
rect -1562 22947 -1528 22963
rect -1562 22895 -1528 22909
rect -1562 22875 -1528 22895
rect -1562 22827 -1528 22837
rect -1562 22803 -1528 22827
rect -1562 22759 -1528 22765
rect -1562 22731 -1528 22759
rect -1562 22691 -1528 22693
rect -1562 22659 -1528 22691
rect -1562 22589 -1528 22621
rect -1562 22587 -1528 22589
rect -1562 22521 -1528 22549
rect -1562 22515 -1528 22521
rect -1562 22453 -1528 22477
rect -1562 22443 -1528 22453
rect -1562 22385 -1528 22405
rect -1562 22371 -1528 22385
rect -1562 22317 -1528 22333
rect -1562 22299 -1528 22317
rect -1562 22249 -1528 22261
rect -1562 22227 -1528 22249
rect -1562 22181 -1528 22189
rect -1562 22155 -1528 22181
rect -1304 23099 -1270 23125
rect -1304 23091 -1270 23099
rect -1304 23031 -1270 23053
rect -1304 23019 -1270 23031
rect -1304 22963 -1270 22981
rect -1304 22947 -1270 22963
rect -1304 22895 -1270 22909
rect -1304 22875 -1270 22895
rect -1304 22827 -1270 22837
rect -1304 22803 -1270 22827
rect -1304 22759 -1270 22765
rect -1304 22731 -1270 22759
rect -1304 22691 -1270 22693
rect -1304 22659 -1270 22691
rect -1304 22589 -1270 22621
rect -1304 22587 -1270 22589
rect -1304 22521 -1270 22549
rect -1304 22515 -1270 22521
rect -1304 22453 -1270 22477
rect -1304 22443 -1270 22453
rect -1304 22385 -1270 22405
rect -1304 22371 -1270 22385
rect -1304 22317 -1270 22333
rect -1304 22299 -1270 22317
rect -1304 22249 -1270 22261
rect -1304 22227 -1270 22249
rect -1304 22181 -1270 22189
rect -1304 22155 -1270 22181
rect -1046 23099 -1012 23125
rect -1046 23091 -1012 23099
rect -1046 23031 -1012 23053
rect -1046 23019 -1012 23031
rect -1046 22963 -1012 22981
rect -1046 22947 -1012 22963
rect -1046 22895 -1012 22909
rect -1046 22875 -1012 22895
rect -1046 22827 -1012 22837
rect -1046 22803 -1012 22827
rect -1046 22759 -1012 22765
rect -1046 22731 -1012 22759
rect -1046 22691 -1012 22693
rect -1046 22659 -1012 22691
rect -1046 22589 -1012 22621
rect -1046 22587 -1012 22589
rect -1046 22521 -1012 22549
rect -1046 22515 -1012 22521
rect -1046 22453 -1012 22477
rect -1046 22443 -1012 22453
rect -1046 22385 -1012 22405
rect -1046 22371 -1012 22385
rect -1046 22317 -1012 22333
rect -1046 22299 -1012 22317
rect -1046 22249 -1012 22261
rect -1046 22227 -1012 22249
rect -1046 22181 -1012 22189
rect -1046 22155 -1012 22181
rect -788 23099 -754 23125
rect -788 23091 -754 23099
rect -788 23031 -754 23053
rect -788 23019 -754 23031
rect -788 22963 -754 22981
rect -788 22947 -754 22963
rect -788 22895 -754 22909
rect -788 22875 -754 22895
rect -788 22827 -754 22837
rect -788 22803 -754 22827
rect -788 22759 -754 22765
rect -788 22731 -754 22759
rect -788 22691 -754 22693
rect -788 22659 -754 22691
rect -788 22589 -754 22621
rect -788 22587 -754 22589
rect -788 22521 -754 22549
rect -788 22515 -754 22521
rect -788 22453 -754 22477
rect -788 22443 -754 22453
rect -788 22385 -754 22405
rect -788 22371 -754 22385
rect -788 22317 -754 22333
rect -788 22299 -754 22317
rect -788 22249 -754 22261
rect -788 22227 -754 22249
rect -788 22181 -754 22189
rect -788 22155 -754 22181
rect -530 23099 -496 23125
rect -530 23091 -496 23099
rect -530 23031 -496 23053
rect -530 23019 -496 23031
rect -530 22963 -496 22981
rect -530 22947 -496 22963
rect -530 22895 -496 22909
rect -530 22875 -496 22895
rect -530 22827 -496 22837
rect -530 22803 -496 22827
rect -530 22759 -496 22765
rect -530 22731 -496 22759
rect -530 22691 -496 22693
rect -530 22659 -496 22691
rect -530 22589 -496 22621
rect -530 22587 -496 22589
rect -530 22521 -496 22549
rect -530 22515 -496 22521
rect -530 22453 -496 22477
rect -530 22443 -496 22453
rect -530 22385 -496 22405
rect -530 22371 -496 22385
rect -530 22317 -496 22333
rect -530 22299 -496 22317
rect -530 22249 -496 22261
rect -530 22227 -496 22249
rect -530 22181 -496 22189
rect -530 22155 -496 22181
rect -272 23099 -238 23125
rect -272 23091 -238 23099
rect -272 23031 -238 23053
rect -272 23019 -238 23031
rect -272 22963 -238 22981
rect -272 22947 -238 22963
rect -272 22895 -238 22909
rect -272 22875 -238 22895
rect -272 22827 -238 22837
rect -272 22803 -238 22827
rect -272 22759 -238 22765
rect -272 22731 -238 22759
rect -272 22691 -238 22693
rect -272 22659 -238 22691
rect -272 22589 -238 22621
rect -272 22587 -238 22589
rect -272 22521 -238 22549
rect -272 22515 -238 22521
rect -272 22453 -238 22477
rect -272 22443 -238 22453
rect -272 22385 -238 22405
rect -272 22371 -238 22385
rect -272 22317 -238 22333
rect -272 22299 -238 22317
rect -272 22249 -238 22261
rect -272 22227 -238 22249
rect -272 22181 -238 22189
rect -272 22155 -238 22181
rect -14 23099 20 23125
rect -14 23091 20 23099
rect -14 23031 20 23053
rect -14 23019 20 23031
rect -14 22963 20 22981
rect -14 22947 20 22963
rect -14 22895 20 22909
rect -14 22875 20 22895
rect -14 22827 20 22837
rect -14 22803 20 22827
rect -14 22759 20 22765
rect -14 22731 20 22759
rect -14 22691 20 22693
rect -14 22659 20 22691
rect -14 22589 20 22621
rect -14 22587 20 22589
rect -14 22521 20 22549
rect -14 22515 20 22521
rect -14 22453 20 22477
rect -14 22443 20 22453
rect -14 22385 20 22405
rect -14 22371 20 22385
rect -14 22317 20 22333
rect -14 22299 20 22317
rect -14 22249 20 22261
rect -14 22227 20 22249
rect -14 22181 20 22189
rect -14 22155 20 22181
rect 244 23099 278 23125
rect 244 23091 278 23099
rect 244 23031 278 23053
rect 244 23019 278 23031
rect 244 22963 278 22981
rect 244 22947 278 22963
rect 244 22895 278 22909
rect 244 22875 278 22895
rect 244 22827 278 22837
rect 244 22803 278 22827
rect 244 22759 278 22765
rect 244 22731 278 22759
rect 244 22691 278 22693
rect 244 22659 278 22691
rect 244 22589 278 22621
rect 244 22587 278 22589
rect 244 22521 278 22549
rect 244 22515 278 22521
rect 244 22453 278 22477
rect 244 22443 278 22453
rect 244 22385 278 22405
rect 244 22371 278 22385
rect 244 22317 278 22333
rect 244 22299 278 22317
rect 244 22249 278 22261
rect 244 22227 278 22249
rect 244 22181 278 22189
rect 244 22155 278 22181
rect 502 23099 536 23125
rect 502 23091 536 23099
rect 502 23031 536 23053
rect 502 23019 536 23031
rect 502 22963 536 22981
rect 502 22947 536 22963
rect 502 22895 536 22909
rect 502 22875 536 22895
rect 502 22827 536 22837
rect 502 22803 536 22827
rect 502 22759 536 22765
rect 502 22731 536 22759
rect 502 22691 536 22693
rect 502 22659 536 22691
rect 502 22589 536 22621
rect 502 22587 536 22589
rect 502 22521 536 22549
rect 502 22515 536 22521
rect 502 22453 536 22477
rect 502 22443 536 22453
rect 502 22385 536 22405
rect 502 22371 536 22385
rect 502 22317 536 22333
rect 502 22299 536 22317
rect 502 22249 536 22261
rect 502 22227 536 22249
rect 502 22181 536 22189
rect 502 22155 536 22181
rect 760 23099 794 23125
rect 760 23091 794 23099
rect 760 23031 794 23053
rect 760 23019 794 23031
rect 760 22963 794 22981
rect 760 22947 794 22963
rect 760 22895 794 22909
rect 760 22875 794 22895
rect 760 22827 794 22837
rect 760 22803 794 22827
rect 760 22759 794 22765
rect 760 22731 794 22759
rect 760 22691 794 22693
rect 760 22659 794 22691
rect 760 22589 794 22621
rect 760 22587 794 22589
rect 760 22521 794 22549
rect 760 22515 794 22521
rect 760 22453 794 22477
rect 760 22443 794 22453
rect 760 22385 794 22405
rect 760 22371 794 22385
rect 760 22317 794 22333
rect 760 22299 794 22317
rect 760 22249 794 22261
rect 760 22227 794 22249
rect 760 22181 794 22189
rect 760 22155 794 22181
rect 1018 23099 1052 23125
rect 1018 23091 1052 23099
rect 1018 23031 1052 23053
rect 1018 23019 1052 23031
rect 1018 22963 1052 22981
rect 1018 22947 1052 22963
rect 1018 22895 1052 22909
rect 1018 22875 1052 22895
rect 1018 22827 1052 22837
rect 1018 22803 1052 22827
rect 1018 22759 1052 22765
rect 1018 22731 1052 22759
rect 1018 22691 1052 22693
rect 1018 22659 1052 22691
rect 1018 22589 1052 22621
rect 1018 22587 1052 22589
rect 1018 22521 1052 22549
rect 1018 22515 1052 22521
rect 1018 22453 1052 22477
rect 1018 22443 1052 22453
rect 1018 22385 1052 22405
rect 1018 22371 1052 22385
rect 1018 22317 1052 22333
rect 1018 22299 1052 22317
rect 1018 22249 1052 22261
rect 1018 22227 1052 22249
rect 1018 22181 1052 22189
rect 1018 22155 1052 22181
rect 1276 23099 1310 23125
rect 1276 23091 1310 23099
rect 1276 23031 1310 23053
rect 1276 23019 1310 23031
rect 1276 22963 1310 22981
rect 1276 22947 1310 22963
rect 1276 22895 1310 22909
rect 1276 22875 1310 22895
rect 1276 22827 1310 22837
rect 1276 22803 1310 22827
rect 1276 22759 1310 22765
rect 1276 22731 1310 22759
rect 1276 22691 1310 22693
rect 1276 22659 1310 22691
rect 1276 22589 1310 22621
rect 1276 22587 1310 22589
rect 1276 22521 1310 22549
rect 1276 22515 1310 22521
rect 1276 22453 1310 22477
rect 1276 22443 1310 22453
rect 1276 22385 1310 22405
rect 1276 22371 1310 22385
rect 1276 22317 1310 22333
rect 1276 22299 1310 22317
rect 1276 22249 1310 22261
rect 1276 22227 1310 22249
rect 1276 22181 1310 22189
rect 1276 22155 1310 22181
rect 1534 23099 1568 23125
rect 1534 23091 1568 23099
rect 1534 23031 1568 23053
rect 1534 23019 1568 23031
rect 1534 22963 1568 22981
rect 1534 22947 1568 22963
rect 1534 22895 1568 22909
rect 1534 22875 1568 22895
rect 1534 22827 1568 22837
rect 1534 22803 1568 22827
rect 1534 22759 1568 22765
rect 1534 22731 1568 22759
rect 1534 22691 1568 22693
rect 1534 22659 1568 22691
rect 1534 22589 1568 22621
rect 1534 22587 1568 22589
rect 1534 22521 1568 22549
rect 1534 22515 1568 22521
rect 1534 22453 1568 22477
rect 1534 22443 1568 22453
rect 1534 22385 1568 22405
rect 1534 22371 1568 22385
rect 1534 22317 1568 22333
rect 1534 22299 1568 22317
rect 1534 22249 1568 22261
rect 1534 22227 1568 22249
rect 1534 22181 1568 22189
rect 1534 22155 1568 22181
rect -1469 22068 -1467 22102
rect -1467 22068 -1435 22102
rect -1397 22068 -1365 22102
rect -1365 22068 -1363 22102
rect -1211 22068 -1209 22102
rect -1209 22068 -1177 22102
rect -1139 22068 -1107 22102
rect -1107 22068 -1105 22102
rect -953 22068 -951 22102
rect -951 22068 -919 22102
rect -881 22068 -849 22102
rect -849 22068 -847 22102
rect -695 22068 -693 22102
rect -693 22068 -661 22102
rect -623 22068 -591 22102
rect -591 22068 -589 22102
rect -437 22068 -435 22102
rect -435 22068 -403 22102
rect -365 22068 -333 22102
rect -333 22068 -331 22102
rect -179 22068 -177 22102
rect -177 22068 -145 22102
rect -107 22068 -75 22102
rect -75 22068 -73 22102
rect 79 22068 81 22102
rect 81 22068 113 22102
rect 151 22068 183 22102
rect 183 22068 185 22102
rect 337 22068 339 22102
rect 339 22068 371 22102
rect 409 22068 441 22102
rect 441 22068 443 22102
rect 595 22068 597 22102
rect 597 22068 629 22102
rect 667 22068 699 22102
rect 699 22068 701 22102
rect 853 22068 855 22102
rect 855 22068 887 22102
rect 925 22068 957 22102
rect 957 22068 959 22102
rect 1111 22068 1113 22102
rect 1113 22068 1145 22102
rect 1183 22068 1215 22102
rect 1215 22068 1217 22102
rect 1369 22068 1371 22102
rect 1371 22068 1403 22102
rect 1441 22068 1473 22102
rect 1473 22068 1475 22102
rect -806 21966 -796 22000
rect -796 21966 -772 22000
rect -734 21966 -728 22000
rect -728 21966 -700 22000
rect -662 21966 -660 22000
rect -660 21966 -628 22000
rect -590 21966 -558 22000
rect -558 21966 -556 22000
rect -518 21966 -490 22000
rect -490 21966 -484 22000
rect -446 21966 -422 22000
rect -422 21966 -412 22000
rect -374 21966 -354 22000
rect -354 21966 -340 22000
rect -302 21966 -286 22000
rect -286 21966 -268 22000
rect -230 21966 -218 22000
rect -218 21966 -196 22000
rect -158 21966 -150 22000
rect -150 21966 -124 22000
rect -86 21966 -82 22000
rect -82 21966 -52 22000
rect -14 21966 20 22000
rect 58 21966 88 22000
rect 88 21966 92 22000
rect 130 21966 156 22000
rect 156 21966 164 22000
rect 202 21966 224 22000
rect 224 21966 236 22000
rect 274 21966 292 22000
rect 292 21966 308 22000
rect 346 21966 360 22000
rect 360 21966 380 22000
rect 418 21966 428 22000
rect 428 21966 452 22000
rect 490 21966 496 22000
rect 496 21966 524 22000
rect 562 21966 564 22000
rect 564 21966 596 22000
rect 634 21966 666 22000
rect 666 21966 668 22000
rect 706 21966 734 22000
rect 734 21966 740 22000
rect 778 21966 802 22000
rect 802 21966 812 22000
rect -916 21760 -900 21794
rect -900 21760 -882 21794
rect -844 21760 -832 21794
rect -832 21760 -810 21794
rect -772 21760 -764 21794
rect -764 21760 -738 21794
rect -700 21760 -696 21794
rect -696 21760 -666 21794
rect -628 21760 -594 21794
rect -556 21760 -526 21794
rect -526 21760 -522 21794
rect -484 21760 -458 21794
rect -458 21760 -450 21794
rect -412 21760 -390 21794
rect -390 21760 -378 21794
rect -340 21760 -322 21794
rect -322 21760 -306 21794
rect -268 21760 -254 21794
rect -254 21760 -234 21794
rect -196 21760 -186 21794
rect -186 21760 -162 21794
rect -124 21760 -118 21794
rect -118 21760 -90 21794
rect -52 21760 -50 21794
rect -50 21760 -18 21794
rect 20 21760 52 21794
rect 52 21760 54 21794
rect 92 21760 120 21794
rect 120 21760 126 21794
rect 164 21760 188 21794
rect 188 21760 198 21794
rect 236 21760 256 21794
rect 256 21760 270 21794
rect 308 21760 324 21794
rect 324 21760 342 21794
rect 380 21760 392 21794
rect 392 21760 414 21794
rect 452 21760 460 21794
rect 460 21760 486 21794
rect 524 21760 528 21794
rect 528 21760 558 21794
rect 596 21760 630 21794
rect 668 21760 698 21794
rect 698 21760 702 21794
rect 740 21760 766 21794
rect 766 21760 774 21794
rect 812 21760 834 21794
rect 834 21760 846 21794
rect 884 21760 902 21794
rect 902 21760 918 21794
rect -1729 21658 -1727 21692
rect -1727 21658 -1695 21692
rect -1657 21658 -1625 21692
rect -1625 21658 -1623 21692
rect -1471 21658 -1469 21692
rect -1469 21658 -1437 21692
rect -1399 21658 -1367 21692
rect -1367 21658 -1365 21692
rect -1213 21658 -1211 21692
rect -1211 21658 -1179 21692
rect -1141 21658 -1109 21692
rect -1109 21658 -1107 21692
rect -955 21658 -953 21692
rect -953 21658 -921 21692
rect -883 21658 -851 21692
rect -851 21658 -849 21692
rect -697 21658 -695 21692
rect -695 21658 -663 21692
rect -625 21658 -593 21692
rect -593 21658 -591 21692
rect -439 21658 -437 21692
rect -437 21658 -405 21692
rect -367 21658 -335 21692
rect -335 21658 -333 21692
rect -181 21658 -179 21692
rect -179 21658 -147 21692
rect -109 21658 -77 21692
rect -77 21658 -75 21692
rect 77 21658 79 21692
rect 79 21658 111 21692
rect 149 21658 181 21692
rect 181 21658 183 21692
rect 335 21658 337 21692
rect 337 21658 369 21692
rect 407 21658 439 21692
rect 439 21658 441 21692
rect 593 21658 595 21692
rect 595 21658 627 21692
rect 665 21658 697 21692
rect 697 21658 699 21692
rect 851 21658 853 21692
rect 853 21658 885 21692
rect 923 21658 955 21692
rect 955 21658 957 21692
rect 1109 21658 1111 21692
rect 1111 21658 1143 21692
rect 1181 21658 1213 21692
rect 1213 21658 1215 21692
rect 1367 21658 1369 21692
rect 1369 21658 1401 21692
rect 1439 21658 1471 21692
rect 1471 21658 1473 21692
rect 1625 21658 1627 21692
rect 1627 21658 1659 21692
rect 1697 21658 1729 21692
rect 1729 21658 1731 21692
rect -1822 21579 -1788 21605
rect -1822 21571 -1788 21579
rect -1822 21511 -1788 21533
rect -1822 21499 -1788 21511
rect -1822 21443 -1788 21461
rect -1822 21427 -1788 21443
rect -1822 21375 -1788 21389
rect -1822 21355 -1788 21375
rect -1822 21307 -1788 21317
rect -1822 21283 -1788 21307
rect -1822 21239 -1788 21245
rect -1822 21211 -1788 21239
rect -1822 21171 -1788 21173
rect -1822 21139 -1788 21171
rect -1822 21069 -1788 21101
rect -1822 21067 -1788 21069
rect -1822 21001 -1788 21029
rect -1822 20995 -1788 21001
rect -1822 20933 -1788 20957
rect -1822 20923 -1788 20933
rect -1822 20865 -1788 20885
rect -1822 20851 -1788 20865
rect -1822 20797 -1788 20813
rect -1822 20779 -1788 20797
rect -1822 20729 -1788 20741
rect -1822 20707 -1788 20729
rect -1822 20661 -1788 20669
rect -1822 20635 -1788 20661
rect -1564 21579 -1530 21605
rect -1564 21571 -1530 21579
rect -1564 21511 -1530 21533
rect -1564 21499 -1530 21511
rect -1564 21443 -1530 21461
rect -1564 21427 -1530 21443
rect -1564 21375 -1530 21389
rect -1564 21355 -1530 21375
rect -1564 21307 -1530 21317
rect -1564 21283 -1530 21307
rect -1564 21239 -1530 21245
rect -1564 21211 -1530 21239
rect -1564 21171 -1530 21173
rect -1564 21139 -1530 21171
rect -1564 21069 -1530 21101
rect -1564 21067 -1530 21069
rect -1564 21001 -1530 21029
rect -1564 20995 -1530 21001
rect -1564 20933 -1530 20957
rect -1564 20923 -1530 20933
rect -1564 20865 -1530 20885
rect -1564 20851 -1530 20865
rect -1564 20797 -1530 20813
rect -1564 20779 -1530 20797
rect -1564 20729 -1530 20741
rect -1564 20707 -1530 20729
rect -1564 20661 -1530 20669
rect -1564 20635 -1530 20661
rect -1306 21579 -1272 21605
rect -1306 21571 -1272 21579
rect -1306 21511 -1272 21533
rect -1306 21499 -1272 21511
rect -1306 21443 -1272 21461
rect -1306 21427 -1272 21443
rect -1306 21375 -1272 21389
rect -1306 21355 -1272 21375
rect -1306 21307 -1272 21317
rect -1306 21283 -1272 21307
rect -1306 21239 -1272 21245
rect -1306 21211 -1272 21239
rect -1306 21171 -1272 21173
rect -1306 21139 -1272 21171
rect -1306 21069 -1272 21101
rect -1306 21067 -1272 21069
rect -1306 21001 -1272 21029
rect -1306 20995 -1272 21001
rect -1306 20933 -1272 20957
rect -1306 20923 -1272 20933
rect -1306 20865 -1272 20885
rect -1306 20851 -1272 20865
rect -1306 20797 -1272 20813
rect -1306 20779 -1272 20797
rect -1306 20729 -1272 20741
rect -1306 20707 -1272 20729
rect -1306 20661 -1272 20669
rect -1306 20635 -1272 20661
rect -1048 21579 -1014 21605
rect -1048 21571 -1014 21579
rect -1048 21511 -1014 21533
rect -1048 21499 -1014 21511
rect -1048 21443 -1014 21461
rect -1048 21427 -1014 21443
rect -1048 21375 -1014 21389
rect -1048 21355 -1014 21375
rect -1048 21307 -1014 21317
rect -1048 21283 -1014 21307
rect -1048 21239 -1014 21245
rect -1048 21211 -1014 21239
rect -1048 21171 -1014 21173
rect -1048 21139 -1014 21171
rect -1048 21069 -1014 21101
rect -1048 21067 -1014 21069
rect -1048 21001 -1014 21029
rect -1048 20995 -1014 21001
rect -1048 20933 -1014 20957
rect -1048 20923 -1014 20933
rect -1048 20865 -1014 20885
rect -1048 20851 -1014 20865
rect -1048 20797 -1014 20813
rect -1048 20779 -1014 20797
rect -1048 20729 -1014 20741
rect -1048 20707 -1014 20729
rect -1048 20661 -1014 20669
rect -1048 20635 -1014 20661
rect -790 21579 -756 21605
rect -790 21571 -756 21579
rect -790 21511 -756 21533
rect -790 21499 -756 21511
rect -790 21443 -756 21461
rect -790 21427 -756 21443
rect -790 21375 -756 21389
rect -790 21355 -756 21375
rect -790 21307 -756 21317
rect -790 21283 -756 21307
rect -790 21239 -756 21245
rect -790 21211 -756 21239
rect -790 21171 -756 21173
rect -790 21139 -756 21171
rect -790 21069 -756 21101
rect -790 21067 -756 21069
rect -790 21001 -756 21029
rect -790 20995 -756 21001
rect -790 20933 -756 20957
rect -790 20923 -756 20933
rect -790 20865 -756 20885
rect -790 20851 -756 20865
rect -790 20797 -756 20813
rect -790 20779 -756 20797
rect -790 20729 -756 20741
rect -790 20707 -756 20729
rect -790 20661 -756 20669
rect -790 20635 -756 20661
rect -532 21579 -498 21605
rect -532 21571 -498 21579
rect -532 21511 -498 21533
rect -532 21499 -498 21511
rect -532 21443 -498 21461
rect -532 21427 -498 21443
rect -532 21375 -498 21389
rect -532 21355 -498 21375
rect -532 21307 -498 21317
rect -532 21283 -498 21307
rect -532 21239 -498 21245
rect -532 21211 -498 21239
rect -532 21171 -498 21173
rect -532 21139 -498 21171
rect -532 21069 -498 21101
rect -532 21067 -498 21069
rect -532 21001 -498 21029
rect -532 20995 -498 21001
rect -532 20933 -498 20957
rect -532 20923 -498 20933
rect -532 20865 -498 20885
rect -532 20851 -498 20865
rect -532 20797 -498 20813
rect -532 20779 -498 20797
rect -532 20729 -498 20741
rect -532 20707 -498 20729
rect -532 20661 -498 20669
rect -532 20635 -498 20661
rect -274 21579 -240 21605
rect -274 21571 -240 21579
rect -274 21511 -240 21533
rect -274 21499 -240 21511
rect -274 21443 -240 21461
rect -274 21427 -240 21443
rect -274 21375 -240 21389
rect -274 21355 -240 21375
rect -274 21307 -240 21317
rect -274 21283 -240 21307
rect -274 21239 -240 21245
rect -274 21211 -240 21239
rect -274 21171 -240 21173
rect -274 21139 -240 21171
rect -274 21069 -240 21101
rect -274 21067 -240 21069
rect -274 21001 -240 21029
rect -274 20995 -240 21001
rect -274 20933 -240 20957
rect -274 20923 -240 20933
rect -274 20865 -240 20885
rect -274 20851 -240 20865
rect -274 20797 -240 20813
rect -274 20779 -240 20797
rect -274 20729 -240 20741
rect -274 20707 -240 20729
rect -274 20661 -240 20669
rect -274 20635 -240 20661
rect -16 21579 18 21605
rect -16 21571 18 21579
rect -16 21511 18 21533
rect -16 21499 18 21511
rect -16 21443 18 21461
rect -16 21427 18 21443
rect -16 21375 18 21389
rect -16 21355 18 21375
rect -16 21307 18 21317
rect -16 21283 18 21307
rect -16 21239 18 21245
rect -16 21211 18 21239
rect -16 21171 18 21173
rect -16 21139 18 21171
rect -16 21069 18 21101
rect -16 21067 18 21069
rect -16 21001 18 21029
rect -16 20995 18 21001
rect -16 20933 18 20957
rect -16 20923 18 20933
rect -16 20865 18 20885
rect -16 20851 18 20865
rect -16 20797 18 20813
rect -16 20779 18 20797
rect -16 20729 18 20741
rect -16 20707 18 20729
rect -16 20661 18 20669
rect -16 20635 18 20661
rect 242 21579 276 21605
rect 242 21571 276 21579
rect 242 21511 276 21533
rect 242 21499 276 21511
rect 242 21443 276 21461
rect 242 21427 276 21443
rect 242 21375 276 21389
rect 242 21355 276 21375
rect 242 21307 276 21317
rect 242 21283 276 21307
rect 242 21239 276 21245
rect 242 21211 276 21239
rect 242 21171 276 21173
rect 242 21139 276 21171
rect 242 21069 276 21101
rect 242 21067 276 21069
rect 242 21001 276 21029
rect 242 20995 276 21001
rect 242 20933 276 20957
rect 242 20923 276 20933
rect 242 20865 276 20885
rect 242 20851 276 20865
rect 242 20797 276 20813
rect 242 20779 276 20797
rect 242 20729 276 20741
rect 242 20707 276 20729
rect 242 20661 276 20669
rect 242 20635 276 20661
rect 500 21579 534 21605
rect 500 21571 534 21579
rect 500 21511 534 21533
rect 500 21499 534 21511
rect 500 21443 534 21461
rect 500 21427 534 21443
rect 500 21375 534 21389
rect 500 21355 534 21375
rect 500 21307 534 21317
rect 500 21283 534 21307
rect 500 21239 534 21245
rect 500 21211 534 21239
rect 500 21171 534 21173
rect 500 21139 534 21171
rect 500 21069 534 21101
rect 500 21067 534 21069
rect 500 21001 534 21029
rect 500 20995 534 21001
rect 500 20933 534 20957
rect 500 20923 534 20933
rect 500 20865 534 20885
rect 500 20851 534 20865
rect 500 20797 534 20813
rect 500 20779 534 20797
rect 500 20729 534 20741
rect 500 20707 534 20729
rect 500 20661 534 20669
rect 500 20635 534 20661
rect 758 21579 792 21605
rect 758 21571 792 21579
rect 758 21511 792 21533
rect 758 21499 792 21511
rect 758 21443 792 21461
rect 758 21427 792 21443
rect 758 21375 792 21389
rect 758 21355 792 21375
rect 758 21307 792 21317
rect 758 21283 792 21307
rect 758 21239 792 21245
rect 758 21211 792 21239
rect 758 21171 792 21173
rect 758 21139 792 21171
rect 758 21069 792 21101
rect 758 21067 792 21069
rect 758 21001 792 21029
rect 758 20995 792 21001
rect 758 20933 792 20957
rect 758 20923 792 20933
rect 758 20865 792 20885
rect 758 20851 792 20865
rect 758 20797 792 20813
rect 758 20779 792 20797
rect 758 20729 792 20741
rect 758 20707 792 20729
rect 758 20661 792 20669
rect 758 20635 792 20661
rect 1016 21579 1050 21605
rect 1016 21571 1050 21579
rect 1016 21511 1050 21533
rect 1016 21499 1050 21511
rect 1016 21443 1050 21461
rect 1016 21427 1050 21443
rect 1016 21375 1050 21389
rect 1016 21355 1050 21375
rect 1016 21307 1050 21317
rect 1016 21283 1050 21307
rect 1016 21239 1050 21245
rect 1016 21211 1050 21239
rect 1016 21171 1050 21173
rect 1016 21139 1050 21171
rect 1016 21069 1050 21101
rect 1016 21067 1050 21069
rect 1016 21001 1050 21029
rect 1016 20995 1050 21001
rect 1016 20933 1050 20957
rect 1016 20923 1050 20933
rect 1016 20865 1050 20885
rect 1016 20851 1050 20865
rect 1016 20797 1050 20813
rect 1016 20779 1050 20797
rect 1016 20729 1050 20741
rect 1016 20707 1050 20729
rect 1016 20661 1050 20669
rect 1016 20635 1050 20661
rect 1274 21579 1308 21605
rect 1274 21571 1308 21579
rect 1274 21511 1308 21533
rect 1274 21499 1308 21511
rect 1274 21443 1308 21461
rect 1274 21427 1308 21443
rect 1274 21375 1308 21389
rect 1274 21355 1308 21375
rect 1274 21307 1308 21317
rect 1274 21283 1308 21307
rect 1274 21239 1308 21245
rect 1274 21211 1308 21239
rect 1274 21171 1308 21173
rect 1274 21139 1308 21171
rect 1274 21069 1308 21101
rect 1274 21067 1308 21069
rect 1274 21001 1308 21029
rect 1274 20995 1308 21001
rect 1274 20933 1308 20957
rect 1274 20923 1308 20933
rect 1274 20865 1308 20885
rect 1274 20851 1308 20865
rect 1274 20797 1308 20813
rect 1274 20779 1308 20797
rect 1274 20729 1308 20741
rect 1274 20707 1308 20729
rect 1274 20661 1308 20669
rect 1274 20635 1308 20661
rect 1532 21579 1566 21605
rect 1532 21571 1566 21579
rect 1532 21511 1566 21533
rect 1532 21499 1566 21511
rect 1532 21443 1566 21461
rect 1532 21427 1566 21443
rect 1532 21375 1566 21389
rect 1532 21355 1566 21375
rect 1532 21307 1566 21317
rect 1532 21283 1566 21307
rect 1532 21239 1566 21245
rect 1532 21211 1566 21239
rect 1532 21171 1566 21173
rect 1532 21139 1566 21171
rect 1532 21069 1566 21101
rect 1532 21067 1566 21069
rect 1532 21001 1566 21029
rect 1532 20995 1566 21001
rect 1532 20933 1566 20957
rect 1532 20923 1566 20933
rect 1532 20865 1566 20885
rect 1532 20851 1566 20865
rect 1532 20797 1566 20813
rect 1532 20779 1566 20797
rect 1532 20729 1566 20741
rect 1532 20707 1566 20729
rect 1532 20661 1566 20669
rect 1532 20635 1566 20661
rect 1790 21579 1824 21605
rect 1790 21571 1824 21579
rect 1790 21511 1824 21533
rect 1790 21499 1824 21511
rect 1790 21443 1824 21461
rect 1790 21427 1824 21443
rect 1790 21375 1824 21389
rect 1790 21355 1824 21375
rect 1790 21307 1824 21317
rect 1790 21283 1824 21307
rect 1790 21239 1824 21245
rect 1790 21211 1824 21239
rect 1790 21171 1824 21173
rect 1790 21139 1824 21171
rect 1790 21069 1824 21101
rect 1790 21067 1824 21069
rect 1790 21001 1824 21029
rect 1790 20995 1824 21001
rect 1790 20933 1824 20957
rect 1790 20923 1824 20933
rect 1790 20865 1824 20885
rect 1790 20851 1824 20865
rect 1790 20797 1824 20813
rect 1790 20779 1824 20797
rect 1790 20729 1824 20741
rect 1790 20707 1824 20729
rect 1790 20661 1824 20669
rect 1790 20635 1824 20661
rect -1729 20548 -1727 20582
rect -1727 20548 -1695 20582
rect -1657 20548 -1625 20582
rect -1625 20548 -1623 20582
rect -1471 20548 -1469 20582
rect -1469 20548 -1437 20582
rect -1399 20548 -1367 20582
rect -1367 20548 -1365 20582
rect -1213 20548 -1211 20582
rect -1211 20548 -1179 20582
rect -1141 20548 -1109 20582
rect -1109 20548 -1107 20582
rect -955 20548 -953 20582
rect -953 20548 -921 20582
rect -883 20548 -851 20582
rect -851 20548 -849 20582
rect -697 20548 -695 20582
rect -695 20548 -663 20582
rect -625 20548 -593 20582
rect -593 20548 -591 20582
rect -439 20548 -437 20582
rect -437 20548 -405 20582
rect -367 20548 -335 20582
rect -335 20548 -333 20582
rect -181 20548 -179 20582
rect -179 20548 -147 20582
rect -109 20548 -77 20582
rect -77 20548 -75 20582
rect 77 20548 79 20582
rect 79 20548 111 20582
rect 149 20548 181 20582
rect 181 20548 183 20582
rect 335 20548 337 20582
rect 337 20548 369 20582
rect 407 20548 439 20582
rect 439 20548 441 20582
rect 593 20548 595 20582
rect 595 20548 627 20582
rect 665 20548 697 20582
rect 697 20548 699 20582
rect 851 20548 853 20582
rect 853 20548 885 20582
rect 923 20548 955 20582
rect 955 20548 957 20582
rect 1109 20548 1111 20582
rect 1111 20548 1143 20582
rect 1181 20548 1213 20582
rect 1213 20548 1215 20582
rect 1367 20548 1369 20582
rect 1369 20548 1401 20582
rect 1439 20548 1471 20582
rect 1471 20548 1473 20582
rect 1625 20548 1627 20582
rect 1627 20548 1659 20582
rect 1697 20548 1729 20582
rect 1729 20548 1731 20582
rect -916 20446 -900 20480
rect -900 20446 -882 20480
rect -844 20446 -832 20480
rect -832 20446 -810 20480
rect -772 20446 -764 20480
rect -764 20446 -738 20480
rect -700 20446 -696 20480
rect -696 20446 -666 20480
rect -628 20446 -594 20480
rect -556 20446 -526 20480
rect -526 20446 -522 20480
rect -484 20446 -458 20480
rect -458 20446 -450 20480
rect -412 20446 -390 20480
rect -390 20446 -378 20480
rect -340 20446 -322 20480
rect -322 20446 -306 20480
rect -268 20446 -254 20480
rect -254 20446 -234 20480
rect -196 20446 -186 20480
rect -186 20446 -162 20480
rect -124 20446 -118 20480
rect -118 20446 -90 20480
rect -52 20446 -50 20480
rect -50 20446 -18 20480
rect 20 20446 52 20480
rect 52 20446 54 20480
rect 92 20446 120 20480
rect 120 20446 126 20480
rect 164 20446 188 20480
rect 188 20446 198 20480
rect 236 20446 256 20480
rect 256 20446 270 20480
rect 308 20446 324 20480
rect 324 20446 342 20480
rect 380 20446 392 20480
rect 392 20446 414 20480
rect 452 20446 460 20480
rect 460 20446 486 20480
rect 524 20446 528 20480
rect 528 20446 558 20480
rect 596 20446 630 20480
rect 668 20446 698 20480
rect 698 20446 702 20480
rect 740 20446 766 20480
rect 766 20446 774 20480
rect 812 20446 834 20480
rect 834 20446 846 20480
rect 884 20446 902 20480
rect 902 20446 918 20480
rect -3220 19546 -3060 19640
rect -2160 19546 -2000 19640
rect -700 19546 -540 19640
rect 520 19546 680 19640
rect 2000 19546 2160 19640
rect 3000 19546 3160 19640
rect -3220 19512 -3060 19546
rect -2160 19512 -2000 19546
rect -700 19512 -540 19546
rect 520 19512 680 19546
rect 2000 19512 2160 19546
rect 3000 19512 3160 19546
rect -3220 19480 -3060 19512
rect -2160 19480 -2000 19512
rect -700 19480 -540 19512
rect 520 19480 680 19512
rect 2000 19480 2160 19512
rect 3000 19480 3160 19512
rect -3579 19398 -2603 19432
rect -2343 19398 -1367 19432
rect -1107 19398 -131 19432
rect 129 19398 1105 19432
rect 1365 19398 2341 19432
rect 2601 19398 3577 19432
rect -3672 19202 -3638 19370
rect -2544 19202 -2510 19370
rect -2436 19202 -2402 19370
rect -1308 19202 -1274 19370
rect -1200 19202 -1166 19370
rect -72 19202 -38 19370
rect 36 19202 70 19370
rect 1164 19202 1198 19370
rect 1272 19202 1306 19370
rect 2400 19202 2434 19370
rect 2508 19202 2542 19370
rect 3636 19202 3670 19370
rect -3579 19140 -2603 19174
rect -2343 19140 -1367 19174
rect -1107 19140 -131 19174
rect 129 19140 1105 19174
rect 1365 19140 2341 19174
rect 2601 19140 3577 19174
rect -3220 19026 -3060 19060
rect -2160 19026 -2000 19060
rect -700 19026 -540 19060
rect 520 19026 680 19060
rect 2000 19026 2160 19060
rect 3000 19026 3160 19060
rect -3220 18956 -3060 19026
rect -2160 18956 -2000 19026
rect -700 18956 -540 19026
rect 520 18956 680 19026
rect 2000 18956 2160 19026
rect 3000 18956 3160 19026
rect -3220 18922 -3060 18956
rect -2160 18922 -2000 18956
rect -700 18922 -540 18956
rect 520 18922 680 18956
rect 2000 18922 2160 18956
rect 3000 18922 3160 18956
rect -3220 18900 -3060 18922
rect -2160 18900 -2000 18922
rect -700 18900 -540 18922
rect 520 18900 680 18922
rect 2000 18900 2160 18922
rect 3000 18900 3160 18922
rect -3579 18808 -2603 18842
rect -2343 18808 -1367 18842
rect -1107 18808 -131 18842
rect 129 18808 1105 18842
rect 1365 18808 2341 18842
rect 2601 18808 3577 18842
rect -3672 18612 -3638 18780
rect -2544 18612 -2510 18780
rect -2436 18612 -2402 18780
rect -1308 18612 -1274 18780
rect -1200 18612 -1166 18780
rect -72 18612 -38 18780
rect 36 18612 70 18780
rect 1164 18612 1198 18780
rect 1272 18612 1306 18780
rect 2400 18612 2434 18780
rect 2508 18612 2542 18780
rect 3636 18612 3670 18780
rect -3579 18550 -2603 18584
rect -2343 18550 -1367 18584
rect -1107 18550 -131 18584
rect 129 18550 1105 18584
rect 1365 18550 2341 18584
rect 2601 18550 3577 18584
rect -818 18018 -592 18052
rect -350 18018 -124 18052
rect 118 18018 344 18052
rect 586 18018 812 18052
rect -902 17822 -868 17990
rect -542 17822 -508 17990
rect -434 17822 -400 17990
rect -74 17822 -40 17990
rect 34 17822 68 17990
rect 394 17822 428 17990
rect 502 17822 536 17990
rect 862 17822 896 17990
rect -818 17760 -592 17794
rect -350 17760 -124 17794
rect 118 17760 344 17794
rect 586 17760 812 17794
rect -840 17646 -620 17680
rect -320 17646 -100 17680
rect 100 17646 320 17680
rect 650 17646 870 17680
rect -840 17541 -620 17646
rect -320 17541 -100 17646
rect 100 17541 320 17646
rect 650 17541 870 17646
rect -840 17530 -688 17541
rect -688 17530 -620 17541
rect -320 17530 -100 17541
rect 100 17530 320 17541
rect 650 17530 686 17541
rect 686 17530 870 17541
rect -598 17393 -122 17427
rect 120 17393 596 17427
rect -682 17297 -648 17365
rect -72 17297 -38 17365
rect 36 17297 70 17365
rect 646 17297 680 17365
rect -598 17235 -122 17269
rect 120 17235 596 17269
rect -3200 17016 -3020 17120
rect -2060 17016 -1880 17120
rect -1080 17016 -900 17130
rect -310 17121 -130 17130
rect 130 17121 310 17130
rect -310 17016 -130 17121
rect 130 17016 310 17121
rect 850 17016 1030 17120
rect 1920 17016 2100 17130
rect 2920 17016 3100 17130
rect -3200 16990 -3020 17016
rect -2060 16990 -1880 17016
rect -1080 17000 -900 17016
rect -310 17000 -130 17016
rect 130 17000 310 17016
rect 850 16990 1030 17016
rect 1920 17000 2100 17016
rect 2920 17000 3100 17016
rect -3533 16868 -2557 16902
rect -2315 16868 -1339 16902
rect -1097 16868 -121 16902
rect 121 16868 1097 16902
rect 1339 16868 2315 16902
rect 2557 16868 3533 16902
rect -3617 16672 -3583 16840
rect -2507 16672 -2473 16840
rect -2399 16672 -2365 16840
rect -1289 16672 -1255 16840
rect -1181 16672 -1147 16840
rect -71 16672 -37 16840
rect 37 16672 71 16840
rect 1147 16672 1181 16840
rect 1255 16672 1289 16840
rect 2365 16672 2399 16840
rect 2473 16672 2507 16840
rect 3583 16672 3617 16840
rect -3533 16610 -2557 16644
rect -2315 16610 -1339 16644
rect -1097 16610 -121 16644
rect 121 16610 1097 16644
rect 1339 16610 2315 16644
rect 2557 16610 3533 16644
rect -2827 15749 -1713 16146
rect -1307 15749 -193 16146
rect 203 15755 1317 16152
rect 1713 15755 2827 16152
rect -3240 15100 -3120 15220
rect 3130 15100 3250 15220
rect -3240 12100 -3120 12220
rect 3130 12100 3250 12220
rect -3240 9100 -3120 9220
rect 3130 9100 3250 9220
rect -3240 6100 -3120 6220
rect 3130 6100 3250 6220
rect -3240 3100 -3120 3220
rect 3130 3100 3250 3220
rect -2827 1518 -1713 1915
rect -1307 1518 -193 1915
rect 203 1524 1317 1921
rect 1713 1524 2827 1921
<< metal1 >>
rect -7130 31926 -6700 31950
rect -7130 30812 -7116 31926
rect -6719 30812 -6700 31926
rect -7130 30660 -6700 30812
rect -7922 30620 -6700 30660
rect -7922 30560 -7912 30620
rect -7852 30560 -7792 30620
rect -7732 30560 -6700 30620
rect -7922 30520 -6700 30560
rect -7130 30426 -6700 30520
rect -7130 29312 -7116 30426
rect -6719 29312 -6700 30426
rect -7130 29300 -6700 29312
rect -4710 31926 -4270 31950
rect -4710 30812 -4685 31926
rect -4288 30812 -4270 31926
rect 4148 31896 4698 31930
rect -672 31387 708 31450
rect -672 31148 -629 31387
rect -1635 31143 -629 31148
rect -385 31143 421 31387
rect 665 31148 708 31387
rect 665 31143 1645 31148
rect -1635 31142 1645 31143
rect -1635 31108 -1596 31142
rect -1562 31108 -1524 31142
rect -1490 31108 -1452 31142
rect -1418 31108 -1380 31142
rect -1346 31108 -1308 31142
rect -1274 31108 -1236 31142
rect -1202 31108 -1164 31142
rect -1130 31108 -1092 31142
rect -1058 31108 -1020 31142
rect -986 31108 -948 31142
rect -914 31108 -876 31142
rect -842 31108 -804 31142
rect -770 31108 -732 31142
rect -698 31108 -660 31142
rect -626 31108 -588 31142
rect -554 31108 -516 31142
rect -482 31108 -444 31142
rect -410 31108 -372 31142
rect -338 31108 -300 31142
rect -266 31108 -228 31142
rect -194 31108 -156 31142
rect -122 31108 -84 31142
rect -50 31108 -12 31142
rect 22 31108 60 31142
rect 94 31108 132 31142
rect 166 31108 204 31142
rect 238 31108 276 31142
rect 310 31108 348 31142
rect 382 31108 420 31142
rect 454 31108 492 31142
rect 526 31108 564 31142
rect 598 31108 636 31142
rect 670 31108 708 31142
rect 742 31108 780 31142
rect 814 31108 852 31142
rect 886 31108 924 31142
rect 958 31108 996 31142
rect 1030 31108 1068 31142
rect 1102 31108 1140 31142
rect 1174 31108 1212 31142
rect 1246 31108 1284 31142
rect 1318 31108 1356 31142
rect 1390 31108 1428 31142
rect 1462 31108 1500 31142
rect 1534 31108 1572 31142
rect 1606 31108 1645 31142
rect -1635 31102 1645 31108
rect -4710 30620 -4270 30812
rect -3322 31040 3338 31050
rect -3322 31006 -3093 31040
rect -3059 31006 -2935 31040
rect -2901 31006 -2777 31040
rect -2743 31006 -2619 31040
rect -2585 31006 -2461 31040
rect -2427 31006 -2303 31040
rect -2269 31006 -2145 31040
rect -2111 31006 -1987 31040
rect -1953 31006 -1829 31040
rect -1795 31006 -1671 31040
rect -1637 31006 -1513 31040
rect -1479 31006 -1355 31040
rect -1321 31006 -1197 31040
rect -1163 31006 -1039 31040
rect -1005 31006 -881 31040
rect -847 31006 -723 31040
rect -689 31006 -565 31040
rect -531 31006 -407 31040
rect -373 31006 -249 31040
rect -215 31006 -91 31040
rect -57 31006 67 31040
rect 101 31006 225 31040
rect 259 31006 383 31040
rect 417 31006 541 31040
rect 575 31006 699 31040
rect 733 31006 857 31040
rect 891 31006 1015 31040
rect 1049 31006 1173 31040
rect 1207 31006 1331 31040
rect 1365 31006 1489 31040
rect 1523 31006 1647 31040
rect 1681 31006 1805 31040
rect 1839 31006 1963 31040
rect 1997 31006 2121 31040
rect 2155 31006 2279 31040
rect 2313 31006 2437 31040
rect 2471 31006 2595 31040
rect 2629 31006 2753 31040
rect 2787 31006 2911 31040
rect 2945 31006 3069 31040
rect 3103 31006 3338 31040
rect -3322 31000 3338 31006
rect -3322 30620 -3242 31000
rect -3178 30944 -3132 30959
rect -3178 30920 -3172 30944
rect -3202 30911 -3172 30920
rect -3138 30920 -3132 30944
rect -3020 30944 -2974 30959
rect -3138 30911 -3112 30920
rect -3202 30859 -3183 30911
rect -3131 30859 -3112 30911
rect -3202 30850 -3172 30859
rect -3178 30838 -3172 30850
rect -3138 30850 -3112 30859
rect -3020 30910 -3014 30944
rect -2980 30910 -2974 30944
rect -2862 30944 -2816 30959
rect -2862 30920 -2856 30944
rect -3020 30872 -2974 30910
rect -3138 30838 -3132 30850
rect -3178 30800 -3132 30838
rect -3178 30766 -3172 30800
rect -3138 30766 -3132 30800
rect -3178 30728 -3132 30766
rect -3178 30694 -3172 30728
rect -3138 30694 -3132 30728
rect -3178 30680 -3132 30694
rect -3020 30838 -3014 30872
rect -2980 30838 -2974 30872
rect -2882 30911 -2856 30920
rect -2822 30920 -2816 30944
rect -2704 30944 -2658 30959
rect -2822 30911 -2792 30920
rect -2882 30859 -2863 30911
rect -2811 30859 -2792 30911
rect -2882 30850 -2856 30859
rect -3020 30800 -2974 30838
rect -3020 30766 -3014 30800
rect -2980 30766 -2974 30800
rect -3020 30728 -2974 30766
rect -3020 30694 -3014 30728
rect -2980 30694 -2974 30728
rect -4710 30426 -3242 30620
rect -3202 30671 -3112 30680
rect -3202 30619 -3183 30671
rect -3131 30619 -3112 30671
rect -3202 30610 -3112 30619
rect -3020 30656 -2974 30694
rect -2862 30838 -2856 30850
rect -2822 30850 -2792 30859
rect -2704 30910 -2698 30944
rect -2664 30910 -2658 30944
rect -2546 30944 -2500 30959
rect -2546 30920 -2540 30944
rect -2704 30872 -2658 30910
rect -2822 30838 -2816 30850
rect -2862 30800 -2816 30838
rect -2862 30766 -2856 30800
rect -2822 30766 -2816 30800
rect -2862 30728 -2816 30766
rect -2862 30694 -2856 30728
rect -2822 30694 -2816 30728
rect -2862 30680 -2816 30694
rect -2704 30838 -2698 30872
rect -2664 30838 -2658 30872
rect -2572 30911 -2540 30920
rect -2506 30920 -2500 30944
rect -2388 30944 -2342 30959
rect -2506 30911 -2482 30920
rect -2572 30859 -2553 30911
rect -2501 30859 -2482 30911
rect -2572 30850 -2540 30859
rect -2704 30800 -2658 30838
rect -2704 30766 -2698 30800
rect -2664 30766 -2658 30800
rect -2704 30728 -2658 30766
rect -2704 30694 -2698 30728
rect -2664 30694 -2658 30728
rect -3020 30622 -3014 30656
rect -2980 30622 -2974 30656
rect -4710 29312 -4685 30426
rect -4288 30330 -3242 30426
rect -4288 29312 -4270 30330
rect -3322 29920 -3242 30330
rect -3178 30584 -3132 30610
rect -3178 30550 -3172 30584
rect -3138 30550 -3132 30584
rect -3178 30512 -3132 30550
rect -3178 30478 -3172 30512
rect -3138 30478 -3132 30512
rect -3178 30440 -3132 30478
rect -3178 30406 -3172 30440
rect -3138 30406 -3132 30440
rect -3178 30368 -3132 30406
rect -3178 30334 -3172 30368
rect -3138 30334 -3132 30368
rect -3178 30296 -3132 30334
rect -3020 30584 -2974 30622
rect -2882 30671 -2792 30680
rect -2882 30619 -2863 30671
rect -2811 30619 -2792 30671
rect -2882 30610 -2792 30619
rect -2704 30656 -2658 30694
rect -2546 30838 -2540 30850
rect -2506 30850 -2482 30859
rect -2388 30910 -2382 30944
rect -2348 30910 -2342 30944
rect -2230 30944 -2184 30959
rect -2230 30920 -2224 30944
rect -2388 30872 -2342 30910
rect -2506 30838 -2500 30850
rect -2546 30800 -2500 30838
rect -2546 30766 -2540 30800
rect -2506 30766 -2500 30800
rect -2546 30728 -2500 30766
rect -2546 30694 -2540 30728
rect -2506 30694 -2500 30728
rect -2546 30680 -2500 30694
rect -2388 30838 -2382 30872
rect -2348 30838 -2342 30872
rect -2252 30911 -2224 30920
rect -2190 30920 -2184 30944
rect -2072 30944 -2026 30959
rect -2190 30911 -2162 30920
rect -2252 30859 -2233 30911
rect -2181 30859 -2162 30911
rect -2252 30850 -2224 30859
rect -2388 30800 -2342 30838
rect -2388 30766 -2382 30800
rect -2348 30766 -2342 30800
rect -2388 30728 -2342 30766
rect -2388 30694 -2382 30728
rect -2348 30694 -2342 30728
rect -2704 30622 -2698 30656
rect -2664 30622 -2658 30656
rect -3020 30550 -3014 30584
rect -2980 30550 -2974 30584
rect -3020 30512 -2974 30550
rect -3020 30478 -3014 30512
rect -2980 30478 -2974 30512
rect -3020 30440 -2974 30478
rect -3020 30406 -3014 30440
rect -2980 30406 -2974 30440
rect -3020 30368 -2974 30406
rect -3020 30334 -3014 30368
rect -2980 30334 -2974 30368
rect -3020 30310 -2974 30334
rect -2862 30584 -2816 30610
rect -2862 30550 -2856 30584
rect -2822 30550 -2816 30584
rect -2862 30512 -2816 30550
rect -2862 30478 -2856 30512
rect -2822 30478 -2816 30512
rect -2862 30440 -2816 30478
rect -2862 30406 -2856 30440
rect -2822 30406 -2816 30440
rect -2862 30368 -2816 30406
rect -2862 30334 -2856 30368
rect -2822 30334 -2816 30368
rect -3178 30262 -3172 30296
rect -3138 30262 -3132 30296
rect -3178 30224 -3132 30262
rect -3042 30301 -2952 30310
rect -3042 30249 -3023 30301
rect -2971 30249 -2952 30301
rect -3042 30240 -2952 30249
rect -2862 30296 -2816 30334
rect -2704 30584 -2658 30622
rect -2572 30671 -2482 30680
rect -2572 30619 -2553 30671
rect -2501 30619 -2482 30671
rect -2572 30610 -2482 30619
rect -2388 30656 -2342 30694
rect -2230 30838 -2224 30850
rect -2190 30850 -2162 30859
rect -2072 30910 -2066 30944
rect -2032 30910 -2026 30944
rect -1914 30944 -1868 30959
rect -1914 30920 -1908 30944
rect -2072 30872 -2026 30910
rect -2190 30838 -2184 30850
rect -2230 30800 -2184 30838
rect -2230 30766 -2224 30800
rect -2190 30766 -2184 30800
rect -2230 30728 -2184 30766
rect -2230 30694 -2224 30728
rect -2190 30694 -2184 30728
rect -2230 30680 -2184 30694
rect -2072 30838 -2066 30872
rect -2032 30838 -2026 30872
rect -1942 30911 -1908 30920
rect -1874 30920 -1868 30944
rect -1756 30944 -1710 30959
rect -1874 30911 -1852 30920
rect -1942 30859 -1923 30911
rect -1871 30859 -1852 30911
rect -1942 30850 -1908 30859
rect -2072 30800 -2026 30838
rect -2072 30766 -2066 30800
rect -2032 30766 -2026 30800
rect -2072 30728 -2026 30766
rect -2072 30694 -2066 30728
rect -2032 30694 -2026 30728
rect -2388 30622 -2382 30656
rect -2348 30622 -2342 30656
rect -2704 30550 -2698 30584
rect -2664 30550 -2658 30584
rect -2704 30512 -2658 30550
rect -2704 30478 -2698 30512
rect -2664 30478 -2658 30512
rect -2704 30440 -2658 30478
rect -2704 30406 -2698 30440
rect -2664 30406 -2658 30440
rect -2704 30368 -2658 30406
rect -2704 30334 -2698 30368
rect -2664 30334 -2658 30368
rect -2704 30310 -2658 30334
rect -2546 30584 -2500 30610
rect -2546 30550 -2540 30584
rect -2506 30550 -2500 30584
rect -2546 30512 -2500 30550
rect -2546 30478 -2540 30512
rect -2506 30478 -2500 30512
rect -2546 30440 -2500 30478
rect -2546 30406 -2540 30440
rect -2506 30406 -2500 30440
rect -2546 30368 -2500 30406
rect -2546 30334 -2540 30368
rect -2506 30334 -2500 30368
rect -2862 30262 -2856 30296
rect -2822 30262 -2816 30296
rect -3178 30190 -3172 30224
rect -3138 30190 -3132 30224
rect -3178 30152 -3132 30190
rect -3178 30118 -3172 30152
rect -3138 30118 -3132 30152
rect -3178 30080 -3132 30118
rect -3178 30046 -3172 30080
rect -3138 30046 -3132 30080
rect -3020 30224 -2974 30240
rect -3020 30190 -3014 30224
rect -2980 30190 -2974 30224
rect -3020 30152 -2974 30190
rect -3020 30118 -3014 30152
rect -2980 30118 -2974 30152
rect -3020 30080 -2974 30118
rect -3020 30070 -3014 30080
rect -3178 30008 -3132 30046
rect -3178 29974 -3172 30008
rect -3138 29974 -3132 30008
rect -3042 30061 -3014 30070
rect -2980 30070 -2974 30080
rect -2862 30224 -2816 30262
rect -2732 30301 -2642 30310
rect -2732 30249 -2713 30301
rect -2661 30249 -2642 30301
rect -2732 30240 -2642 30249
rect -2546 30296 -2500 30334
rect -2388 30584 -2342 30622
rect -2252 30671 -2162 30680
rect -2252 30619 -2233 30671
rect -2181 30619 -2162 30671
rect -2252 30610 -2162 30619
rect -2072 30656 -2026 30694
rect -1914 30838 -1908 30850
rect -1874 30850 -1852 30859
rect -1756 30910 -1750 30944
rect -1716 30910 -1710 30944
rect -1598 30944 -1552 30959
rect -1598 30920 -1592 30944
rect -1756 30872 -1710 30910
rect -1874 30838 -1868 30850
rect -1914 30800 -1868 30838
rect -1914 30766 -1908 30800
rect -1874 30766 -1868 30800
rect -1914 30728 -1868 30766
rect -1914 30694 -1908 30728
rect -1874 30694 -1868 30728
rect -1914 30680 -1868 30694
rect -1756 30838 -1750 30872
rect -1716 30838 -1710 30872
rect -1622 30911 -1592 30920
rect -1558 30920 -1552 30944
rect -1440 30944 -1394 30959
rect -1558 30911 -1532 30920
rect -1622 30859 -1603 30911
rect -1551 30859 -1532 30911
rect -1622 30850 -1592 30859
rect -1756 30800 -1710 30838
rect -1756 30766 -1750 30800
rect -1716 30766 -1710 30800
rect -1756 30728 -1710 30766
rect -1756 30694 -1750 30728
rect -1716 30694 -1710 30728
rect -2072 30622 -2066 30656
rect -2032 30622 -2026 30656
rect -2388 30550 -2382 30584
rect -2348 30550 -2342 30584
rect -2388 30512 -2342 30550
rect -2388 30478 -2382 30512
rect -2348 30478 -2342 30512
rect -2388 30440 -2342 30478
rect -2388 30406 -2382 30440
rect -2348 30406 -2342 30440
rect -2388 30368 -2342 30406
rect -2388 30334 -2382 30368
rect -2348 30334 -2342 30368
rect -2388 30310 -2342 30334
rect -2230 30584 -2184 30610
rect -2230 30550 -2224 30584
rect -2190 30550 -2184 30584
rect -2230 30512 -2184 30550
rect -2230 30478 -2224 30512
rect -2190 30478 -2184 30512
rect -2230 30440 -2184 30478
rect -2230 30406 -2224 30440
rect -2190 30406 -2184 30440
rect -2230 30368 -2184 30406
rect -2230 30334 -2224 30368
rect -2190 30334 -2184 30368
rect -2546 30262 -2540 30296
rect -2506 30262 -2500 30296
rect -2862 30190 -2856 30224
rect -2822 30190 -2816 30224
rect -2862 30152 -2816 30190
rect -2862 30118 -2856 30152
rect -2822 30118 -2816 30152
rect -2862 30080 -2816 30118
rect -2980 30061 -2952 30070
rect -3042 30009 -3023 30061
rect -2971 30009 -2952 30061
rect -3042 30008 -2952 30009
rect -3042 30000 -3014 30008
rect -3178 29959 -3132 29974
rect -3020 29974 -3014 30000
rect -2980 30000 -2952 30008
rect -2862 30046 -2856 30080
rect -2822 30046 -2816 30080
rect -2704 30224 -2658 30240
rect -2704 30190 -2698 30224
rect -2664 30190 -2658 30224
rect -2704 30152 -2658 30190
rect -2704 30118 -2698 30152
rect -2664 30118 -2658 30152
rect -2704 30080 -2658 30118
rect -2704 30070 -2698 30080
rect -2862 30008 -2816 30046
rect -2980 29974 -2974 30000
rect -3020 29959 -2974 29974
rect -2862 29974 -2856 30008
rect -2822 29974 -2816 30008
rect -2732 30061 -2698 30070
rect -2664 30070 -2658 30080
rect -2546 30224 -2500 30262
rect -2412 30301 -2322 30310
rect -2412 30249 -2393 30301
rect -2341 30249 -2322 30301
rect -2412 30240 -2322 30249
rect -2230 30296 -2184 30334
rect -2072 30584 -2026 30622
rect -1942 30671 -1852 30680
rect -1942 30619 -1923 30671
rect -1871 30619 -1852 30671
rect -1942 30610 -1852 30619
rect -1756 30656 -1710 30694
rect -1598 30838 -1592 30850
rect -1558 30850 -1532 30859
rect -1440 30910 -1434 30944
rect -1400 30910 -1394 30944
rect -1282 30944 -1236 30959
rect -1282 30920 -1276 30944
rect -1440 30872 -1394 30910
rect -1558 30838 -1552 30850
rect -1598 30800 -1552 30838
rect -1598 30766 -1592 30800
rect -1558 30766 -1552 30800
rect -1598 30728 -1552 30766
rect -1598 30694 -1592 30728
rect -1558 30694 -1552 30728
rect -1598 30680 -1552 30694
rect -1440 30838 -1434 30872
rect -1400 30838 -1394 30872
rect -1302 30911 -1276 30920
rect -1242 30920 -1236 30944
rect -1124 30944 -1078 30959
rect -1242 30911 -1212 30920
rect -1302 30859 -1283 30911
rect -1231 30859 -1212 30911
rect -1302 30850 -1276 30859
rect -1440 30800 -1394 30838
rect -1440 30766 -1434 30800
rect -1400 30766 -1394 30800
rect -1440 30728 -1394 30766
rect -1440 30694 -1434 30728
rect -1400 30694 -1394 30728
rect -1756 30622 -1750 30656
rect -1716 30622 -1710 30656
rect -2072 30550 -2066 30584
rect -2032 30550 -2026 30584
rect -2072 30512 -2026 30550
rect -2072 30478 -2066 30512
rect -2032 30478 -2026 30512
rect -2072 30440 -2026 30478
rect -2072 30406 -2066 30440
rect -2032 30406 -2026 30440
rect -2072 30368 -2026 30406
rect -2072 30334 -2066 30368
rect -2032 30334 -2026 30368
rect -2072 30310 -2026 30334
rect -1914 30584 -1868 30610
rect -1914 30550 -1908 30584
rect -1874 30550 -1868 30584
rect -1914 30512 -1868 30550
rect -1914 30478 -1908 30512
rect -1874 30478 -1868 30512
rect -1914 30440 -1868 30478
rect -1914 30406 -1908 30440
rect -1874 30406 -1868 30440
rect -1914 30368 -1868 30406
rect -1914 30334 -1908 30368
rect -1874 30334 -1868 30368
rect -2230 30262 -2224 30296
rect -2190 30262 -2184 30296
rect -2546 30190 -2540 30224
rect -2506 30190 -2500 30224
rect -2546 30152 -2500 30190
rect -2546 30118 -2540 30152
rect -2506 30118 -2500 30152
rect -2546 30080 -2500 30118
rect -2664 30061 -2642 30070
rect -2732 30009 -2713 30061
rect -2661 30009 -2642 30061
rect -2732 30008 -2642 30009
rect -2732 30000 -2698 30008
rect -2862 29959 -2816 29974
rect -2704 29974 -2698 30000
rect -2664 30000 -2642 30008
rect -2546 30046 -2540 30080
rect -2506 30046 -2500 30080
rect -2388 30224 -2342 30240
rect -2388 30190 -2382 30224
rect -2348 30190 -2342 30224
rect -2388 30152 -2342 30190
rect -2388 30118 -2382 30152
rect -2348 30118 -2342 30152
rect -2388 30080 -2342 30118
rect -2388 30070 -2382 30080
rect -2546 30008 -2500 30046
rect -2664 29974 -2658 30000
rect -2704 29959 -2658 29974
rect -2546 29974 -2540 30008
rect -2506 29974 -2500 30008
rect -2412 30061 -2382 30070
rect -2348 30070 -2342 30080
rect -2230 30224 -2184 30262
rect -2092 30301 -2002 30310
rect -2092 30249 -2073 30301
rect -2021 30249 -2002 30301
rect -2092 30240 -2002 30249
rect -1914 30296 -1868 30334
rect -1756 30584 -1710 30622
rect -1622 30671 -1532 30680
rect -1622 30619 -1603 30671
rect -1551 30619 -1532 30671
rect -1622 30610 -1532 30619
rect -1440 30656 -1394 30694
rect -1282 30838 -1276 30850
rect -1242 30850 -1212 30859
rect -1124 30910 -1118 30944
rect -1084 30910 -1078 30944
rect -966 30944 -920 30959
rect -966 30920 -960 30944
rect -1124 30872 -1078 30910
rect -1242 30838 -1236 30850
rect -1282 30800 -1236 30838
rect -1282 30766 -1276 30800
rect -1242 30766 -1236 30800
rect -1282 30728 -1236 30766
rect -1282 30694 -1276 30728
rect -1242 30694 -1236 30728
rect -1282 30680 -1236 30694
rect -1124 30838 -1118 30872
rect -1084 30838 -1078 30872
rect -992 30911 -960 30920
rect -926 30920 -920 30944
rect -808 30944 -762 30959
rect -926 30911 -902 30920
rect -992 30859 -973 30911
rect -921 30859 -902 30911
rect -992 30850 -960 30859
rect -1124 30800 -1078 30838
rect -1124 30766 -1118 30800
rect -1084 30766 -1078 30800
rect -1124 30728 -1078 30766
rect -1124 30694 -1118 30728
rect -1084 30694 -1078 30728
rect -1440 30622 -1434 30656
rect -1400 30622 -1394 30656
rect -1756 30550 -1750 30584
rect -1716 30550 -1710 30584
rect -1756 30512 -1710 30550
rect -1756 30478 -1750 30512
rect -1716 30478 -1710 30512
rect -1756 30440 -1710 30478
rect -1756 30406 -1750 30440
rect -1716 30406 -1710 30440
rect -1756 30368 -1710 30406
rect -1756 30334 -1750 30368
rect -1716 30334 -1710 30368
rect -1756 30310 -1710 30334
rect -1598 30584 -1552 30610
rect -1598 30550 -1592 30584
rect -1558 30550 -1552 30584
rect -1598 30512 -1552 30550
rect -1598 30478 -1592 30512
rect -1558 30478 -1552 30512
rect -1598 30440 -1552 30478
rect -1598 30406 -1592 30440
rect -1558 30406 -1552 30440
rect -1598 30368 -1552 30406
rect -1598 30334 -1592 30368
rect -1558 30334 -1552 30368
rect -1914 30262 -1908 30296
rect -1874 30262 -1868 30296
rect -2230 30190 -2224 30224
rect -2190 30190 -2184 30224
rect -2230 30152 -2184 30190
rect -2230 30118 -2224 30152
rect -2190 30118 -2184 30152
rect -2230 30080 -2184 30118
rect -2348 30061 -2322 30070
rect -2412 30009 -2393 30061
rect -2341 30009 -2322 30061
rect -2412 30008 -2322 30009
rect -2412 30000 -2382 30008
rect -2546 29959 -2500 29974
rect -2388 29974 -2382 30000
rect -2348 30000 -2322 30008
rect -2230 30046 -2224 30080
rect -2190 30046 -2184 30080
rect -2072 30224 -2026 30240
rect -2072 30190 -2066 30224
rect -2032 30190 -2026 30224
rect -2072 30152 -2026 30190
rect -2072 30118 -2066 30152
rect -2032 30118 -2026 30152
rect -2072 30080 -2026 30118
rect -2072 30070 -2066 30080
rect -2230 30008 -2184 30046
rect -2348 29974 -2342 30000
rect -2388 29959 -2342 29974
rect -2230 29974 -2224 30008
rect -2190 29974 -2184 30008
rect -2092 30061 -2066 30070
rect -2032 30070 -2026 30080
rect -1914 30224 -1868 30262
rect -1782 30301 -1692 30310
rect -1782 30249 -1763 30301
rect -1711 30249 -1692 30301
rect -1782 30240 -1692 30249
rect -1598 30296 -1552 30334
rect -1440 30584 -1394 30622
rect -1302 30671 -1212 30680
rect -1302 30619 -1283 30671
rect -1231 30619 -1212 30671
rect -1302 30610 -1212 30619
rect -1124 30656 -1078 30694
rect -966 30838 -960 30850
rect -926 30850 -902 30859
rect -808 30910 -802 30944
rect -768 30910 -762 30944
rect -650 30944 -604 30959
rect -650 30920 -644 30944
rect -808 30872 -762 30910
rect -926 30838 -920 30850
rect -966 30800 -920 30838
rect -966 30766 -960 30800
rect -926 30766 -920 30800
rect -966 30728 -920 30766
rect -966 30694 -960 30728
rect -926 30694 -920 30728
rect -966 30680 -920 30694
rect -808 30838 -802 30872
rect -768 30838 -762 30872
rect -672 30911 -644 30920
rect -610 30920 -604 30944
rect -492 30944 -446 30959
rect -610 30911 -582 30920
rect -672 30859 -653 30911
rect -601 30859 -582 30911
rect -672 30850 -644 30859
rect -808 30800 -762 30838
rect -808 30766 -802 30800
rect -768 30766 -762 30800
rect -808 30728 -762 30766
rect -808 30694 -802 30728
rect -768 30694 -762 30728
rect -1124 30622 -1118 30656
rect -1084 30622 -1078 30656
rect -1440 30550 -1434 30584
rect -1400 30550 -1394 30584
rect -1440 30512 -1394 30550
rect -1440 30478 -1434 30512
rect -1400 30478 -1394 30512
rect -1440 30440 -1394 30478
rect -1440 30406 -1434 30440
rect -1400 30406 -1394 30440
rect -1440 30368 -1394 30406
rect -1440 30334 -1434 30368
rect -1400 30334 -1394 30368
rect -1440 30310 -1394 30334
rect -1282 30584 -1236 30610
rect -1282 30550 -1276 30584
rect -1242 30550 -1236 30584
rect -1282 30512 -1236 30550
rect -1282 30478 -1276 30512
rect -1242 30478 -1236 30512
rect -1282 30440 -1236 30478
rect -1282 30406 -1276 30440
rect -1242 30406 -1236 30440
rect -1282 30368 -1236 30406
rect -1282 30334 -1276 30368
rect -1242 30334 -1236 30368
rect -1598 30262 -1592 30296
rect -1558 30262 -1552 30296
rect -1914 30190 -1908 30224
rect -1874 30190 -1868 30224
rect -1914 30152 -1868 30190
rect -1914 30118 -1908 30152
rect -1874 30118 -1868 30152
rect -1914 30080 -1868 30118
rect -2032 30061 -2002 30070
rect -2092 30009 -2073 30061
rect -2021 30009 -2002 30061
rect -2092 30008 -2002 30009
rect -2092 30000 -2066 30008
rect -2230 29959 -2184 29974
rect -2072 29974 -2066 30000
rect -2032 30000 -2002 30008
rect -1914 30046 -1908 30080
rect -1874 30046 -1868 30080
rect -1756 30224 -1710 30240
rect -1756 30190 -1750 30224
rect -1716 30190 -1710 30224
rect -1756 30152 -1710 30190
rect -1756 30118 -1750 30152
rect -1716 30118 -1710 30152
rect -1756 30080 -1710 30118
rect -1756 30070 -1750 30080
rect -1914 30008 -1868 30046
rect -2032 29974 -2026 30000
rect -2072 29959 -2026 29974
rect -1914 29974 -1908 30008
rect -1874 29974 -1868 30008
rect -1782 30061 -1750 30070
rect -1716 30070 -1710 30080
rect -1598 30224 -1552 30262
rect -1462 30301 -1372 30310
rect -1462 30249 -1443 30301
rect -1391 30249 -1372 30301
rect -1462 30240 -1372 30249
rect -1282 30296 -1236 30334
rect -1124 30584 -1078 30622
rect -992 30671 -902 30680
rect -992 30619 -973 30671
rect -921 30619 -902 30671
rect -992 30610 -902 30619
rect -808 30656 -762 30694
rect -650 30838 -644 30850
rect -610 30850 -582 30859
rect -492 30910 -486 30944
rect -452 30910 -446 30944
rect -334 30944 -288 30959
rect -334 30920 -328 30944
rect -492 30872 -446 30910
rect -610 30838 -604 30850
rect -650 30800 -604 30838
rect -650 30766 -644 30800
rect -610 30766 -604 30800
rect -650 30728 -604 30766
rect -650 30694 -644 30728
rect -610 30694 -604 30728
rect -650 30680 -604 30694
rect -492 30838 -486 30872
rect -452 30838 -446 30872
rect -352 30911 -328 30920
rect -294 30920 -288 30944
rect -176 30944 -130 30959
rect -294 30911 -262 30920
rect -352 30859 -333 30911
rect -281 30859 -262 30911
rect -352 30850 -328 30859
rect -492 30800 -446 30838
rect -492 30766 -486 30800
rect -452 30766 -446 30800
rect -492 30728 -446 30766
rect -492 30694 -486 30728
rect -452 30694 -446 30728
rect -808 30622 -802 30656
rect -768 30622 -762 30656
rect -1124 30550 -1118 30584
rect -1084 30550 -1078 30584
rect -1124 30512 -1078 30550
rect -1124 30478 -1118 30512
rect -1084 30478 -1078 30512
rect -1124 30440 -1078 30478
rect -1124 30406 -1118 30440
rect -1084 30406 -1078 30440
rect -1124 30368 -1078 30406
rect -1124 30334 -1118 30368
rect -1084 30334 -1078 30368
rect -1124 30310 -1078 30334
rect -966 30584 -920 30610
rect -966 30550 -960 30584
rect -926 30550 -920 30584
rect -966 30512 -920 30550
rect -966 30478 -960 30512
rect -926 30478 -920 30512
rect -966 30440 -920 30478
rect -966 30406 -960 30440
rect -926 30406 -920 30440
rect -966 30368 -920 30406
rect -966 30334 -960 30368
rect -926 30334 -920 30368
rect -1282 30262 -1276 30296
rect -1242 30262 -1236 30296
rect -1598 30190 -1592 30224
rect -1558 30190 -1552 30224
rect -1598 30152 -1552 30190
rect -1598 30118 -1592 30152
rect -1558 30118 -1552 30152
rect -1598 30080 -1552 30118
rect -1716 30061 -1692 30070
rect -1782 30009 -1763 30061
rect -1711 30009 -1692 30061
rect -1782 30008 -1692 30009
rect -1782 30000 -1750 30008
rect -1914 29959 -1868 29974
rect -1756 29974 -1750 30000
rect -1716 30000 -1692 30008
rect -1598 30046 -1592 30080
rect -1558 30046 -1552 30080
rect -1440 30224 -1394 30240
rect -1440 30190 -1434 30224
rect -1400 30190 -1394 30224
rect -1440 30152 -1394 30190
rect -1440 30118 -1434 30152
rect -1400 30118 -1394 30152
rect -1440 30080 -1394 30118
rect -1440 30070 -1434 30080
rect -1598 30008 -1552 30046
rect -1716 29974 -1710 30000
rect -1756 29959 -1710 29974
rect -1598 29974 -1592 30008
rect -1558 29974 -1552 30008
rect -1462 30061 -1434 30070
rect -1400 30070 -1394 30080
rect -1282 30224 -1236 30262
rect -1152 30301 -1062 30310
rect -1152 30249 -1133 30301
rect -1081 30249 -1062 30301
rect -1152 30240 -1062 30249
rect -966 30296 -920 30334
rect -808 30584 -762 30622
rect -672 30671 -582 30680
rect -672 30619 -653 30671
rect -601 30619 -582 30671
rect -672 30610 -582 30619
rect -492 30656 -446 30694
rect -334 30838 -328 30850
rect -294 30850 -262 30859
rect -176 30910 -170 30944
rect -136 30910 -130 30944
rect -18 30944 28 30959
rect -18 30920 -12 30944
rect -176 30872 -130 30910
rect -294 30838 -288 30850
rect -334 30800 -288 30838
rect -334 30766 -328 30800
rect -294 30766 -288 30800
rect -334 30728 -288 30766
rect -334 30694 -328 30728
rect -294 30694 -288 30728
rect -334 30680 -288 30694
rect -176 30838 -170 30872
rect -136 30838 -130 30872
rect -42 30911 -12 30920
rect 22 30920 28 30944
rect 140 30944 186 30959
rect 22 30911 48 30920
rect -42 30859 -23 30911
rect 29 30859 48 30911
rect -42 30850 -12 30859
rect -176 30800 -130 30838
rect -176 30766 -170 30800
rect -136 30766 -130 30800
rect -176 30728 -130 30766
rect -176 30694 -170 30728
rect -136 30694 -130 30728
rect -492 30622 -486 30656
rect -452 30622 -446 30656
rect -808 30550 -802 30584
rect -768 30550 -762 30584
rect -808 30512 -762 30550
rect -808 30478 -802 30512
rect -768 30478 -762 30512
rect -808 30440 -762 30478
rect -808 30406 -802 30440
rect -768 30406 -762 30440
rect -808 30368 -762 30406
rect -808 30334 -802 30368
rect -768 30334 -762 30368
rect -808 30310 -762 30334
rect -650 30584 -604 30610
rect -650 30550 -644 30584
rect -610 30550 -604 30584
rect -650 30512 -604 30550
rect -650 30478 -644 30512
rect -610 30478 -604 30512
rect -650 30440 -604 30478
rect -650 30406 -644 30440
rect -610 30406 -604 30440
rect -650 30368 -604 30406
rect -650 30334 -644 30368
rect -610 30334 -604 30368
rect -966 30262 -960 30296
rect -926 30262 -920 30296
rect -1282 30190 -1276 30224
rect -1242 30190 -1236 30224
rect -1282 30152 -1236 30190
rect -1282 30118 -1276 30152
rect -1242 30118 -1236 30152
rect -1282 30080 -1236 30118
rect -1400 30061 -1372 30070
rect -1462 30009 -1443 30061
rect -1391 30009 -1372 30061
rect -1462 30008 -1372 30009
rect -1462 30000 -1434 30008
rect -1598 29959 -1552 29974
rect -1440 29974 -1434 30000
rect -1400 30000 -1372 30008
rect -1282 30046 -1276 30080
rect -1242 30046 -1236 30080
rect -1124 30224 -1078 30240
rect -1124 30190 -1118 30224
rect -1084 30190 -1078 30224
rect -1124 30152 -1078 30190
rect -1124 30118 -1118 30152
rect -1084 30118 -1078 30152
rect -1124 30080 -1078 30118
rect -1124 30070 -1118 30080
rect -1282 30008 -1236 30046
rect -1400 29974 -1394 30000
rect -1440 29959 -1394 29974
rect -1282 29974 -1276 30008
rect -1242 29974 -1236 30008
rect -1152 30061 -1118 30070
rect -1084 30070 -1078 30080
rect -966 30224 -920 30262
rect -832 30301 -742 30310
rect -832 30249 -813 30301
rect -761 30249 -742 30301
rect -832 30240 -742 30249
rect -650 30296 -604 30334
rect -492 30584 -446 30622
rect -352 30671 -262 30680
rect -352 30619 -333 30671
rect -281 30619 -262 30671
rect -352 30610 -262 30619
rect -176 30656 -130 30694
rect -18 30838 -12 30850
rect 22 30850 48 30859
rect 140 30910 146 30944
rect 180 30910 186 30944
rect 298 30944 344 30959
rect 298 30920 304 30944
rect 140 30872 186 30910
rect 22 30838 28 30850
rect -18 30800 28 30838
rect -18 30766 -12 30800
rect 22 30766 28 30800
rect -18 30728 28 30766
rect -18 30694 -12 30728
rect 22 30694 28 30728
rect -18 30680 28 30694
rect 140 30838 146 30872
rect 180 30838 186 30872
rect 278 30911 304 30920
rect 338 30920 344 30944
rect 456 30944 502 30959
rect 338 30911 368 30920
rect 278 30859 297 30911
rect 349 30859 368 30911
rect 278 30850 304 30859
rect 140 30800 186 30838
rect 140 30766 146 30800
rect 180 30766 186 30800
rect 140 30728 186 30766
rect 140 30694 146 30728
rect 180 30694 186 30728
rect -176 30622 -170 30656
rect -136 30622 -130 30656
rect -492 30550 -486 30584
rect -452 30550 -446 30584
rect -492 30512 -446 30550
rect -492 30478 -486 30512
rect -452 30478 -446 30512
rect -492 30440 -446 30478
rect -492 30406 -486 30440
rect -452 30406 -446 30440
rect -492 30368 -446 30406
rect -492 30334 -486 30368
rect -452 30334 -446 30368
rect -492 30310 -446 30334
rect -334 30584 -288 30610
rect -334 30550 -328 30584
rect -294 30550 -288 30584
rect -334 30512 -288 30550
rect -334 30478 -328 30512
rect -294 30478 -288 30512
rect -334 30440 -288 30478
rect -334 30406 -328 30440
rect -294 30406 -288 30440
rect -334 30368 -288 30406
rect -334 30334 -328 30368
rect -294 30334 -288 30368
rect -650 30262 -644 30296
rect -610 30262 -604 30296
rect -966 30190 -960 30224
rect -926 30190 -920 30224
rect -966 30152 -920 30190
rect -966 30118 -960 30152
rect -926 30118 -920 30152
rect -966 30080 -920 30118
rect -1084 30061 -1062 30070
rect -1152 30009 -1133 30061
rect -1081 30009 -1062 30061
rect -1152 30008 -1062 30009
rect -1152 30000 -1118 30008
rect -1282 29959 -1236 29974
rect -1124 29974 -1118 30000
rect -1084 30000 -1062 30008
rect -966 30046 -960 30080
rect -926 30046 -920 30080
rect -808 30224 -762 30240
rect -808 30190 -802 30224
rect -768 30190 -762 30224
rect -808 30152 -762 30190
rect -808 30118 -802 30152
rect -768 30118 -762 30152
rect -808 30080 -762 30118
rect -808 30070 -802 30080
rect -966 30008 -920 30046
rect -1084 29974 -1078 30000
rect -1124 29959 -1078 29974
rect -966 29974 -960 30008
rect -926 29974 -920 30008
rect -832 30061 -802 30070
rect -768 30070 -762 30080
rect -650 30224 -604 30262
rect -512 30301 -422 30310
rect -512 30249 -493 30301
rect -441 30249 -422 30301
rect -512 30240 -422 30249
rect -334 30296 -288 30334
rect -176 30584 -130 30622
rect -42 30671 48 30680
rect -42 30619 -23 30671
rect 29 30619 48 30671
rect -42 30610 48 30619
rect 140 30656 186 30694
rect 298 30838 304 30850
rect 338 30850 368 30859
rect 456 30910 462 30944
rect 496 30910 502 30944
rect 614 30944 660 30959
rect 614 30920 620 30944
rect 456 30872 502 30910
rect 338 30838 344 30850
rect 298 30800 344 30838
rect 298 30766 304 30800
rect 338 30766 344 30800
rect 298 30728 344 30766
rect 298 30694 304 30728
rect 338 30694 344 30728
rect 298 30680 344 30694
rect 456 30838 462 30872
rect 496 30838 502 30872
rect 588 30911 620 30920
rect 654 30920 660 30944
rect 772 30944 818 30959
rect 654 30911 678 30920
rect 588 30859 607 30911
rect 659 30859 678 30911
rect 588 30850 620 30859
rect 456 30800 502 30838
rect 456 30766 462 30800
rect 496 30766 502 30800
rect 456 30728 502 30766
rect 456 30694 462 30728
rect 496 30694 502 30728
rect 140 30622 146 30656
rect 180 30622 186 30656
rect -176 30550 -170 30584
rect -136 30550 -130 30584
rect -176 30512 -130 30550
rect -176 30478 -170 30512
rect -136 30478 -130 30512
rect -176 30440 -130 30478
rect -176 30406 -170 30440
rect -136 30406 -130 30440
rect -176 30368 -130 30406
rect -176 30334 -170 30368
rect -136 30334 -130 30368
rect -176 30310 -130 30334
rect -18 30584 28 30610
rect -18 30550 -12 30584
rect 22 30550 28 30584
rect -18 30512 28 30550
rect -18 30478 -12 30512
rect 22 30478 28 30512
rect -18 30440 28 30478
rect -18 30406 -12 30440
rect 22 30406 28 30440
rect -18 30368 28 30406
rect -18 30334 -12 30368
rect 22 30334 28 30368
rect -334 30262 -328 30296
rect -294 30262 -288 30296
rect -650 30190 -644 30224
rect -610 30190 -604 30224
rect -650 30152 -604 30190
rect -650 30118 -644 30152
rect -610 30118 -604 30152
rect -650 30080 -604 30118
rect -768 30061 -742 30070
rect -832 30009 -813 30061
rect -761 30009 -742 30061
rect -832 30008 -742 30009
rect -832 30000 -802 30008
rect -966 29959 -920 29974
rect -808 29974 -802 30000
rect -768 30000 -742 30008
rect -650 30046 -644 30080
rect -610 30046 -604 30080
rect -492 30224 -446 30240
rect -492 30190 -486 30224
rect -452 30190 -446 30224
rect -492 30152 -446 30190
rect -492 30118 -486 30152
rect -452 30118 -446 30152
rect -492 30080 -446 30118
rect -492 30070 -486 30080
rect -650 30008 -604 30046
rect -768 29974 -762 30000
rect -808 29959 -762 29974
rect -650 29974 -644 30008
rect -610 29974 -604 30008
rect -512 30061 -486 30070
rect -452 30070 -446 30080
rect -334 30224 -288 30262
rect -202 30301 -112 30310
rect -202 30249 -183 30301
rect -131 30249 -112 30301
rect -202 30240 -112 30249
rect -18 30296 28 30334
rect 140 30584 186 30622
rect 278 30671 368 30680
rect 278 30619 297 30671
rect 349 30619 368 30671
rect 278 30610 368 30619
rect 456 30656 502 30694
rect 614 30838 620 30850
rect 654 30850 678 30859
rect 772 30910 778 30944
rect 812 30910 818 30944
rect 930 30944 976 30959
rect 930 30920 936 30944
rect 772 30872 818 30910
rect 654 30838 660 30850
rect 614 30800 660 30838
rect 614 30766 620 30800
rect 654 30766 660 30800
rect 614 30728 660 30766
rect 614 30694 620 30728
rect 654 30694 660 30728
rect 614 30680 660 30694
rect 772 30838 778 30872
rect 812 30838 818 30872
rect 908 30911 936 30920
rect 970 30920 976 30944
rect 1088 30944 1134 30959
rect 970 30911 998 30920
rect 908 30859 927 30911
rect 979 30859 998 30911
rect 908 30850 936 30859
rect 772 30800 818 30838
rect 772 30766 778 30800
rect 812 30766 818 30800
rect 772 30728 818 30766
rect 772 30694 778 30728
rect 812 30694 818 30728
rect 456 30622 462 30656
rect 496 30622 502 30656
rect 140 30550 146 30584
rect 180 30550 186 30584
rect 140 30512 186 30550
rect 140 30478 146 30512
rect 180 30478 186 30512
rect 140 30440 186 30478
rect 140 30406 146 30440
rect 180 30406 186 30440
rect 140 30368 186 30406
rect 140 30334 146 30368
rect 180 30334 186 30368
rect 140 30310 186 30334
rect 298 30584 344 30610
rect 298 30550 304 30584
rect 338 30550 344 30584
rect 298 30512 344 30550
rect 298 30478 304 30512
rect 338 30478 344 30512
rect 298 30440 344 30478
rect 298 30406 304 30440
rect 338 30406 344 30440
rect 298 30368 344 30406
rect 298 30334 304 30368
rect 338 30334 344 30368
rect -18 30262 -12 30296
rect 22 30262 28 30296
rect -334 30190 -328 30224
rect -294 30190 -288 30224
rect -334 30152 -288 30190
rect -334 30118 -328 30152
rect -294 30118 -288 30152
rect -334 30080 -288 30118
rect -452 30061 -422 30070
rect -512 30009 -493 30061
rect -441 30009 -422 30061
rect -512 30008 -422 30009
rect -512 30000 -486 30008
rect -650 29959 -604 29974
rect -492 29974 -486 30000
rect -452 30000 -422 30008
rect -334 30046 -328 30080
rect -294 30046 -288 30080
rect -176 30224 -130 30240
rect -176 30190 -170 30224
rect -136 30190 -130 30224
rect -176 30152 -130 30190
rect -176 30118 -170 30152
rect -136 30118 -130 30152
rect -176 30080 -130 30118
rect -176 30070 -170 30080
rect -334 30008 -288 30046
rect -452 29974 -446 30000
rect -492 29959 -446 29974
rect -334 29974 -328 30008
rect -294 29974 -288 30008
rect -202 30061 -170 30070
rect -136 30070 -130 30080
rect -18 30224 28 30262
rect 118 30301 208 30310
rect 118 30249 137 30301
rect 189 30249 208 30301
rect 118 30240 208 30249
rect 298 30296 344 30334
rect 456 30584 502 30622
rect 588 30671 678 30680
rect 588 30619 607 30671
rect 659 30619 678 30671
rect 588 30610 678 30619
rect 772 30656 818 30694
rect 930 30838 936 30850
rect 970 30850 998 30859
rect 1088 30910 1094 30944
rect 1128 30910 1134 30944
rect 1246 30944 1292 30959
rect 1246 30920 1252 30944
rect 1088 30872 1134 30910
rect 970 30838 976 30850
rect 930 30800 976 30838
rect 930 30766 936 30800
rect 970 30766 976 30800
rect 930 30728 976 30766
rect 930 30694 936 30728
rect 970 30694 976 30728
rect 930 30680 976 30694
rect 1088 30838 1094 30872
rect 1128 30838 1134 30872
rect 1228 30911 1252 30920
rect 1286 30920 1292 30944
rect 1404 30944 1450 30959
rect 1286 30911 1318 30920
rect 1228 30859 1247 30911
rect 1299 30859 1318 30911
rect 1228 30850 1252 30859
rect 1088 30800 1134 30838
rect 1088 30766 1094 30800
rect 1128 30766 1134 30800
rect 1088 30728 1134 30766
rect 1088 30694 1094 30728
rect 1128 30694 1134 30728
rect 772 30622 778 30656
rect 812 30622 818 30656
rect 456 30550 462 30584
rect 496 30550 502 30584
rect 456 30512 502 30550
rect 456 30478 462 30512
rect 496 30478 502 30512
rect 456 30440 502 30478
rect 456 30406 462 30440
rect 496 30406 502 30440
rect 456 30368 502 30406
rect 456 30334 462 30368
rect 496 30334 502 30368
rect 456 30310 502 30334
rect 614 30584 660 30610
rect 614 30550 620 30584
rect 654 30550 660 30584
rect 614 30512 660 30550
rect 614 30478 620 30512
rect 654 30478 660 30512
rect 614 30440 660 30478
rect 614 30406 620 30440
rect 654 30406 660 30440
rect 614 30368 660 30406
rect 614 30334 620 30368
rect 654 30334 660 30368
rect 298 30262 304 30296
rect 338 30262 344 30296
rect -18 30190 -12 30224
rect 22 30190 28 30224
rect -18 30152 28 30190
rect -18 30118 -12 30152
rect 22 30118 28 30152
rect -18 30080 28 30118
rect -136 30061 -112 30070
rect -202 30009 -183 30061
rect -131 30009 -112 30061
rect -202 30008 -112 30009
rect -202 30000 -170 30008
rect -334 29959 -288 29974
rect -176 29974 -170 30000
rect -136 30000 -112 30008
rect -18 30046 -12 30080
rect 22 30046 28 30080
rect 140 30224 186 30240
rect 140 30190 146 30224
rect 180 30190 186 30224
rect 140 30152 186 30190
rect 140 30118 146 30152
rect 180 30118 186 30152
rect 140 30080 186 30118
rect 140 30070 146 30080
rect -18 30008 28 30046
rect -136 29974 -130 30000
rect -176 29959 -130 29974
rect -18 29974 -12 30008
rect 22 29974 28 30008
rect 118 30061 146 30070
rect 180 30070 186 30080
rect 298 30224 344 30262
rect 438 30301 528 30310
rect 438 30249 457 30301
rect 509 30249 528 30301
rect 438 30240 528 30249
rect 614 30296 660 30334
rect 772 30584 818 30622
rect 908 30671 998 30680
rect 908 30619 927 30671
rect 979 30619 998 30671
rect 908 30610 998 30619
rect 1088 30656 1134 30694
rect 1246 30838 1252 30850
rect 1286 30850 1318 30859
rect 1404 30910 1410 30944
rect 1444 30910 1450 30944
rect 1562 30944 1608 30959
rect 1562 30920 1568 30944
rect 1404 30872 1450 30910
rect 1286 30838 1292 30850
rect 1246 30800 1292 30838
rect 1246 30766 1252 30800
rect 1286 30766 1292 30800
rect 1246 30728 1292 30766
rect 1246 30694 1252 30728
rect 1286 30694 1292 30728
rect 1246 30680 1292 30694
rect 1404 30838 1410 30872
rect 1444 30838 1450 30872
rect 1538 30911 1568 30920
rect 1602 30920 1608 30944
rect 1720 30944 1766 30959
rect 1602 30911 1628 30920
rect 1538 30859 1557 30911
rect 1609 30859 1628 30911
rect 1538 30850 1568 30859
rect 1404 30800 1450 30838
rect 1404 30766 1410 30800
rect 1444 30766 1450 30800
rect 1404 30728 1450 30766
rect 1404 30694 1410 30728
rect 1444 30694 1450 30728
rect 1088 30622 1094 30656
rect 1128 30622 1134 30656
rect 772 30550 778 30584
rect 812 30550 818 30584
rect 772 30512 818 30550
rect 772 30478 778 30512
rect 812 30478 818 30512
rect 772 30440 818 30478
rect 772 30406 778 30440
rect 812 30406 818 30440
rect 772 30368 818 30406
rect 772 30334 778 30368
rect 812 30334 818 30368
rect 772 30310 818 30334
rect 930 30584 976 30610
rect 930 30550 936 30584
rect 970 30550 976 30584
rect 930 30512 976 30550
rect 930 30478 936 30512
rect 970 30478 976 30512
rect 930 30440 976 30478
rect 930 30406 936 30440
rect 970 30406 976 30440
rect 930 30368 976 30406
rect 930 30334 936 30368
rect 970 30334 976 30368
rect 614 30262 620 30296
rect 654 30262 660 30296
rect 298 30190 304 30224
rect 338 30190 344 30224
rect 298 30152 344 30190
rect 298 30118 304 30152
rect 338 30118 344 30152
rect 298 30080 344 30118
rect 180 30061 208 30070
rect 118 30009 137 30061
rect 189 30009 208 30061
rect 118 30008 208 30009
rect 118 30000 146 30008
rect -18 29959 28 29974
rect 140 29974 146 30000
rect 180 30000 208 30008
rect 298 30046 304 30080
rect 338 30046 344 30080
rect 456 30224 502 30240
rect 456 30190 462 30224
rect 496 30190 502 30224
rect 456 30152 502 30190
rect 456 30118 462 30152
rect 496 30118 502 30152
rect 456 30080 502 30118
rect 456 30070 462 30080
rect 298 30008 344 30046
rect 180 29974 186 30000
rect 140 29959 186 29974
rect 298 29974 304 30008
rect 338 29974 344 30008
rect 438 30061 462 30070
rect 496 30070 502 30080
rect 614 30224 660 30262
rect 748 30301 838 30310
rect 748 30249 767 30301
rect 819 30249 838 30301
rect 748 30240 838 30249
rect 930 30296 976 30334
rect 1088 30584 1134 30622
rect 1228 30671 1318 30680
rect 1228 30619 1247 30671
rect 1299 30619 1318 30671
rect 1228 30610 1318 30619
rect 1404 30656 1450 30694
rect 1562 30838 1568 30850
rect 1602 30850 1628 30859
rect 1720 30910 1726 30944
rect 1760 30910 1766 30944
rect 1878 30944 1924 30959
rect 1878 30920 1884 30944
rect 1720 30872 1766 30910
rect 1602 30838 1608 30850
rect 1562 30800 1608 30838
rect 1562 30766 1568 30800
rect 1602 30766 1608 30800
rect 1562 30728 1608 30766
rect 1562 30694 1568 30728
rect 1602 30694 1608 30728
rect 1562 30680 1608 30694
rect 1720 30838 1726 30872
rect 1760 30838 1766 30872
rect 1858 30911 1884 30920
rect 1918 30920 1924 30944
rect 2036 30944 2082 30959
rect 1918 30911 1948 30920
rect 1858 30859 1877 30911
rect 1929 30859 1948 30911
rect 1858 30850 1884 30859
rect 1720 30800 1766 30838
rect 1720 30766 1726 30800
rect 1760 30766 1766 30800
rect 1720 30728 1766 30766
rect 1720 30694 1726 30728
rect 1760 30694 1766 30728
rect 1404 30622 1410 30656
rect 1444 30622 1450 30656
rect 1088 30550 1094 30584
rect 1128 30550 1134 30584
rect 1088 30512 1134 30550
rect 1088 30478 1094 30512
rect 1128 30478 1134 30512
rect 1088 30440 1134 30478
rect 1088 30406 1094 30440
rect 1128 30406 1134 30440
rect 1088 30368 1134 30406
rect 1088 30334 1094 30368
rect 1128 30334 1134 30368
rect 1088 30310 1134 30334
rect 1246 30584 1292 30610
rect 1246 30550 1252 30584
rect 1286 30550 1292 30584
rect 1246 30512 1292 30550
rect 1246 30478 1252 30512
rect 1286 30478 1292 30512
rect 1246 30440 1292 30478
rect 1246 30406 1252 30440
rect 1286 30406 1292 30440
rect 1246 30368 1292 30406
rect 1246 30334 1252 30368
rect 1286 30334 1292 30368
rect 930 30262 936 30296
rect 970 30262 976 30296
rect 614 30190 620 30224
rect 654 30190 660 30224
rect 614 30152 660 30190
rect 614 30118 620 30152
rect 654 30118 660 30152
rect 614 30080 660 30118
rect 496 30061 528 30070
rect 438 30009 457 30061
rect 509 30009 528 30061
rect 438 30008 528 30009
rect 438 30000 462 30008
rect 298 29959 344 29974
rect 456 29974 462 30000
rect 496 30000 528 30008
rect 614 30046 620 30080
rect 654 30046 660 30080
rect 772 30224 818 30240
rect 772 30190 778 30224
rect 812 30190 818 30224
rect 772 30152 818 30190
rect 772 30118 778 30152
rect 812 30118 818 30152
rect 772 30080 818 30118
rect 772 30070 778 30080
rect 614 30008 660 30046
rect 496 29974 502 30000
rect 456 29959 502 29974
rect 614 29974 620 30008
rect 654 29974 660 30008
rect 748 30061 778 30070
rect 812 30070 818 30080
rect 930 30224 976 30262
rect 1068 30301 1158 30310
rect 1068 30249 1087 30301
rect 1139 30249 1158 30301
rect 1068 30240 1158 30249
rect 1246 30296 1292 30334
rect 1404 30584 1450 30622
rect 1538 30671 1628 30680
rect 1538 30619 1557 30671
rect 1609 30619 1628 30671
rect 1538 30610 1628 30619
rect 1720 30656 1766 30694
rect 1878 30838 1884 30850
rect 1918 30850 1948 30859
rect 2036 30910 2042 30944
rect 2076 30910 2082 30944
rect 2194 30944 2240 30959
rect 2194 30920 2200 30944
rect 2036 30872 2082 30910
rect 1918 30838 1924 30850
rect 1878 30800 1924 30838
rect 1878 30766 1884 30800
rect 1918 30766 1924 30800
rect 1878 30728 1924 30766
rect 1878 30694 1884 30728
rect 1918 30694 1924 30728
rect 1878 30680 1924 30694
rect 2036 30838 2042 30872
rect 2076 30838 2082 30872
rect 2168 30911 2200 30920
rect 2234 30920 2240 30944
rect 2352 30944 2398 30959
rect 2234 30911 2258 30920
rect 2168 30859 2187 30911
rect 2239 30859 2258 30911
rect 2168 30850 2200 30859
rect 2036 30800 2082 30838
rect 2036 30766 2042 30800
rect 2076 30766 2082 30800
rect 2036 30728 2082 30766
rect 2036 30694 2042 30728
rect 2076 30694 2082 30728
rect 1720 30622 1726 30656
rect 1760 30622 1766 30656
rect 1404 30550 1410 30584
rect 1444 30550 1450 30584
rect 1404 30512 1450 30550
rect 1404 30478 1410 30512
rect 1444 30478 1450 30512
rect 1404 30440 1450 30478
rect 1404 30406 1410 30440
rect 1444 30406 1450 30440
rect 1404 30368 1450 30406
rect 1404 30334 1410 30368
rect 1444 30334 1450 30368
rect 1404 30310 1450 30334
rect 1562 30584 1608 30610
rect 1562 30550 1568 30584
rect 1602 30550 1608 30584
rect 1562 30512 1608 30550
rect 1562 30478 1568 30512
rect 1602 30478 1608 30512
rect 1562 30440 1608 30478
rect 1562 30406 1568 30440
rect 1602 30406 1608 30440
rect 1562 30368 1608 30406
rect 1562 30334 1568 30368
rect 1602 30334 1608 30368
rect 1246 30262 1252 30296
rect 1286 30262 1292 30296
rect 930 30190 936 30224
rect 970 30190 976 30224
rect 930 30152 976 30190
rect 930 30118 936 30152
rect 970 30118 976 30152
rect 930 30080 976 30118
rect 812 30061 838 30070
rect 748 30009 767 30061
rect 819 30009 838 30061
rect 748 30008 838 30009
rect 748 30000 778 30008
rect 614 29959 660 29974
rect 772 29974 778 30000
rect 812 30000 838 30008
rect 930 30046 936 30080
rect 970 30046 976 30080
rect 1088 30224 1134 30240
rect 1088 30190 1094 30224
rect 1128 30190 1134 30224
rect 1088 30152 1134 30190
rect 1088 30118 1094 30152
rect 1128 30118 1134 30152
rect 1088 30080 1134 30118
rect 1088 30070 1094 30080
rect 930 30008 976 30046
rect 812 29974 818 30000
rect 772 29959 818 29974
rect 930 29974 936 30008
rect 970 29974 976 30008
rect 1068 30061 1094 30070
rect 1128 30070 1134 30080
rect 1246 30224 1292 30262
rect 1378 30301 1468 30310
rect 1378 30249 1397 30301
rect 1449 30249 1468 30301
rect 1378 30240 1468 30249
rect 1562 30296 1608 30334
rect 1720 30584 1766 30622
rect 1858 30671 1948 30680
rect 1858 30619 1877 30671
rect 1929 30619 1948 30671
rect 1858 30610 1948 30619
rect 2036 30656 2082 30694
rect 2194 30838 2200 30850
rect 2234 30850 2258 30859
rect 2352 30910 2358 30944
rect 2392 30910 2398 30944
rect 2510 30944 2556 30959
rect 2510 30920 2516 30944
rect 2352 30872 2398 30910
rect 2234 30838 2240 30850
rect 2194 30800 2240 30838
rect 2194 30766 2200 30800
rect 2234 30766 2240 30800
rect 2194 30728 2240 30766
rect 2194 30694 2200 30728
rect 2234 30694 2240 30728
rect 2194 30680 2240 30694
rect 2352 30838 2358 30872
rect 2392 30838 2398 30872
rect 2488 30911 2516 30920
rect 2550 30920 2556 30944
rect 2668 30944 2714 30959
rect 2550 30911 2578 30920
rect 2488 30859 2507 30911
rect 2559 30859 2578 30911
rect 2488 30850 2516 30859
rect 2352 30800 2398 30838
rect 2352 30766 2358 30800
rect 2392 30766 2398 30800
rect 2352 30728 2398 30766
rect 2352 30694 2358 30728
rect 2392 30694 2398 30728
rect 2036 30622 2042 30656
rect 2076 30622 2082 30656
rect 1720 30550 1726 30584
rect 1760 30550 1766 30584
rect 1720 30512 1766 30550
rect 1720 30478 1726 30512
rect 1760 30478 1766 30512
rect 1720 30440 1766 30478
rect 1720 30406 1726 30440
rect 1760 30406 1766 30440
rect 1720 30368 1766 30406
rect 1720 30334 1726 30368
rect 1760 30334 1766 30368
rect 1720 30310 1766 30334
rect 1878 30584 1924 30610
rect 1878 30550 1884 30584
rect 1918 30550 1924 30584
rect 1878 30512 1924 30550
rect 1878 30478 1884 30512
rect 1918 30478 1924 30512
rect 1878 30440 1924 30478
rect 1878 30406 1884 30440
rect 1918 30406 1924 30440
rect 1878 30368 1924 30406
rect 1878 30334 1884 30368
rect 1918 30334 1924 30368
rect 1562 30262 1568 30296
rect 1602 30262 1608 30296
rect 1246 30190 1252 30224
rect 1286 30190 1292 30224
rect 1246 30152 1292 30190
rect 1246 30118 1252 30152
rect 1286 30118 1292 30152
rect 1246 30080 1292 30118
rect 1128 30061 1158 30070
rect 1068 30009 1087 30061
rect 1139 30009 1158 30061
rect 1068 30008 1158 30009
rect 1068 30000 1094 30008
rect 930 29959 976 29974
rect 1088 29974 1094 30000
rect 1128 30000 1158 30008
rect 1246 30046 1252 30080
rect 1286 30046 1292 30080
rect 1404 30224 1450 30240
rect 1404 30190 1410 30224
rect 1444 30190 1450 30224
rect 1404 30152 1450 30190
rect 1404 30118 1410 30152
rect 1444 30118 1450 30152
rect 1404 30080 1450 30118
rect 1404 30070 1410 30080
rect 1246 30008 1292 30046
rect 1128 29974 1134 30000
rect 1088 29959 1134 29974
rect 1246 29974 1252 30008
rect 1286 29974 1292 30008
rect 1378 30061 1410 30070
rect 1444 30070 1450 30080
rect 1562 30224 1608 30262
rect 1698 30301 1788 30310
rect 1698 30249 1717 30301
rect 1769 30249 1788 30301
rect 1698 30240 1788 30249
rect 1878 30296 1924 30334
rect 2036 30584 2082 30622
rect 2168 30671 2258 30680
rect 2168 30619 2187 30671
rect 2239 30619 2258 30671
rect 2168 30610 2258 30619
rect 2352 30656 2398 30694
rect 2510 30838 2516 30850
rect 2550 30850 2578 30859
rect 2668 30910 2674 30944
rect 2708 30910 2714 30944
rect 2826 30944 2872 30959
rect 2826 30920 2832 30944
rect 2668 30872 2714 30910
rect 2550 30838 2556 30850
rect 2510 30800 2556 30838
rect 2510 30766 2516 30800
rect 2550 30766 2556 30800
rect 2510 30728 2556 30766
rect 2510 30694 2516 30728
rect 2550 30694 2556 30728
rect 2510 30680 2556 30694
rect 2668 30838 2674 30872
rect 2708 30838 2714 30872
rect 2808 30911 2832 30920
rect 2866 30920 2872 30944
rect 2984 30944 3030 30959
rect 2866 30911 2898 30920
rect 2808 30859 2827 30911
rect 2879 30859 2898 30911
rect 2808 30850 2832 30859
rect 2668 30800 2714 30838
rect 2668 30766 2674 30800
rect 2708 30766 2714 30800
rect 2668 30728 2714 30766
rect 2668 30694 2674 30728
rect 2708 30694 2714 30728
rect 2352 30622 2358 30656
rect 2392 30622 2398 30656
rect 2036 30550 2042 30584
rect 2076 30550 2082 30584
rect 2036 30512 2082 30550
rect 2036 30478 2042 30512
rect 2076 30478 2082 30512
rect 2036 30440 2082 30478
rect 2036 30406 2042 30440
rect 2076 30406 2082 30440
rect 2036 30368 2082 30406
rect 2036 30334 2042 30368
rect 2076 30334 2082 30368
rect 2036 30310 2082 30334
rect 2194 30584 2240 30610
rect 2194 30550 2200 30584
rect 2234 30550 2240 30584
rect 2194 30512 2240 30550
rect 2194 30478 2200 30512
rect 2234 30478 2240 30512
rect 2194 30440 2240 30478
rect 2194 30406 2200 30440
rect 2234 30406 2240 30440
rect 2194 30368 2240 30406
rect 2194 30334 2200 30368
rect 2234 30334 2240 30368
rect 1878 30262 1884 30296
rect 1918 30262 1924 30296
rect 1562 30190 1568 30224
rect 1602 30190 1608 30224
rect 1562 30152 1608 30190
rect 1562 30118 1568 30152
rect 1602 30118 1608 30152
rect 1562 30080 1608 30118
rect 1444 30061 1468 30070
rect 1378 30009 1397 30061
rect 1449 30009 1468 30061
rect 1378 30008 1468 30009
rect 1378 30000 1410 30008
rect 1246 29959 1292 29974
rect 1404 29974 1410 30000
rect 1444 30000 1468 30008
rect 1562 30046 1568 30080
rect 1602 30046 1608 30080
rect 1720 30224 1766 30240
rect 1720 30190 1726 30224
rect 1760 30190 1766 30224
rect 1720 30152 1766 30190
rect 1720 30118 1726 30152
rect 1760 30118 1766 30152
rect 1720 30080 1766 30118
rect 1720 30070 1726 30080
rect 1562 30008 1608 30046
rect 1444 29974 1450 30000
rect 1404 29959 1450 29974
rect 1562 29974 1568 30008
rect 1602 29974 1608 30008
rect 1698 30061 1726 30070
rect 1760 30070 1766 30080
rect 1878 30224 1924 30262
rect 2018 30301 2108 30310
rect 2018 30249 2037 30301
rect 2089 30249 2108 30301
rect 2018 30240 2108 30249
rect 2194 30296 2240 30334
rect 2352 30584 2398 30622
rect 2488 30671 2578 30680
rect 2488 30619 2507 30671
rect 2559 30619 2578 30671
rect 2488 30610 2578 30619
rect 2668 30656 2714 30694
rect 2826 30838 2832 30850
rect 2866 30850 2898 30859
rect 2984 30910 2990 30944
rect 3024 30910 3030 30944
rect 3142 30944 3188 30959
rect 3142 30920 3148 30944
rect 2984 30872 3030 30910
rect 2866 30838 2872 30850
rect 2826 30800 2872 30838
rect 2826 30766 2832 30800
rect 2866 30766 2872 30800
rect 2826 30728 2872 30766
rect 2826 30694 2832 30728
rect 2866 30694 2872 30728
rect 2826 30680 2872 30694
rect 2984 30838 2990 30872
rect 3024 30838 3030 30872
rect 3118 30911 3148 30920
rect 3182 30920 3188 30944
rect 3182 30911 3208 30920
rect 3118 30859 3137 30911
rect 3189 30859 3208 30911
rect 3118 30850 3148 30859
rect 2984 30800 3030 30838
rect 2984 30766 2990 30800
rect 3024 30766 3030 30800
rect 2984 30728 3030 30766
rect 2984 30694 2990 30728
rect 3024 30694 3030 30728
rect 2668 30622 2674 30656
rect 2708 30622 2714 30656
rect 2352 30550 2358 30584
rect 2392 30550 2398 30584
rect 2352 30512 2398 30550
rect 2352 30478 2358 30512
rect 2392 30478 2398 30512
rect 2352 30440 2398 30478
rect 2352 30406 2358 30440
rect 2392 30406 2398 30440
rect 2352 30368 2398 30406
rect 2352 30334 2358 30368
rect 2392 30334 2398 30368
rect 2352 30310 2398 30334
rect 2510 30584 2556 30610
rect 2510 30550 2516 30584
rect 2550 30550 2556 30584
rect 2510 30512 2556 30550
rect 2510 30478 2516 30512
rect 2550 30478 2556 30512
rect 2510 30440 2556 30478
rect 2510 30406 2516 30440
rect 2550 30406 2556 30440
rect 2510 30368 2556 30406
rect 2510 30334 2516 30368
rect 2550 30334 2556 30368
rect 2194 30262 2200 30296
rect 2234 30262 2240 30296
rect 1878 30190 1884 30224
rect 1918 30190 1924 30224
rect 1878 30152 1924 30190
rect 1878 30118 1884 30152
rect 1918 30118 1924 30152
rect 1878 30080 1924 30118
rect 1760 30061 1788 30070
rect 1698 30009 1717 30061
rect 1769 30009 1788 30061
rect 1698 30008 1788 30009
rect 1698 30000 1726 30008
rect 1562 29959 1608 29974
rect 1720 29974 1726 30000
rect 1760 30000 1788 30008
rect 1878 30046 1884 30080
rect 1918 30046 1924 30080
rect 2036 30224 2082 30240
rect 2036 30190 2042 30224
rect 2076 30190 2082 30224
rect 2036 30152 2082 30190
rect 2036 30118 2042 30152
rect 2076 30118 2082 30152
rect 2036 30080 2082 30118
rect 2036 30070 2042 30080
rect 1878 30008 1924 30046
rect 1760 29974 1766 30000
rect 1720 29959 1766 29974
rect 1878 29974 1884 30008
rect 1918 29974 1924 30008
rect 2018 30061 2042 30070
rect 2076 30070 2082 30080
rect 2194 30224 2240 30262
rect 2328 30301 2418 30310
rect 2328 30249 2347 30301
rect 2399 30249 2418 30301
rect 2328 30240 2418 30249
rect 2510 30296 2556 30334
rect 2668 30584 2714 30622
rect 2808 30671 2898 30680
rect 2808 30619 2827 30671
rect 2879 30619 2898 30671
rect 2808 30610 2898 30619
rect 2984 30656 3030 30694
rect 3142 30838 3148 30850
rect 3182 30850 3208 30859
rect 3182 30838 3188 30850
rect 3142 30800 3188 30838
rect 3142 30766 3148 30800
rect 3182 30766 3188 30800
rect 3142 30728 3188 30766
rect 3142 30694 3148 30728
rect 3182 30694 3188 30728
rect 3142 30680 3188 30694
rect 2984 30622 2990 30656
rect 3024 30622 3030 30656
rect 2668 30550 2674 30584
rect 2708 30550 2714 30584
rect 2668 30512 2714 30550
rect 2668 30478 2674 30512
rect 2708 30478 2714 30512
rect 2668 30440 2714 30478
rect 2668 30406 2674 30440
rect 2708 30406 2714 30440
rect 2668 30368 2714 30406
rect 2668 30334 2674 30368
rect 2708 30334 2714 30368
rect 2668 30310 2714 30334
rect 2826 30584 2872 30610
rect 2826 30550 2832 30584
rect 2866 30550 2872 30584
rect 2826 30512 2872 30550
rect 2826 30478 2832 30512
rect 2866 30478 2872 30512
rect 2826 30440 2872 30478
rect 2826 30406 2832 30440
rect 2866 30406 2872 30440
rect 2826 30368 2872 30406
rect 2826 30334 2832 30368
rect 2866 30334 2872 30368
rect 2510 30262 2516 30296
rect 2550 30262 2556 30296
rect 2194 30190 2200 30224
rect 2234 30190 2240 30224
rect 2194 30152 2240 30190
rect 2194 30118 2200 30152
rect 2234 30118 2240 30152
rect 2194 30080 2240 30118
rect 2076 30061 2108 30070
rect 2018 30009 2037 30061
rect 2089 30009 2108 30061
rect 2018 30008 2108 30009
rect 2018 30000 2042 30008
rect 1878 29959 1924 29974
rect 2036 29974 2042 30000
rect 2076 30000 2108 30008
rect 2194 30046 2200 30080
rect 2234 30046 2240 30080
rect 2352 30224 2398 30240
rect 2352 30190 2358 30224
rect 2392 30190 2398 30224
rect 2352 30152 2398 30190
rect 2352 30118 2358 30152
rect 2392 30118 2398 30152
rect 2352 30080 2398 30118
rect 2352 30070 2358 30080
rect 2194 30008 2240 30046
rect 2076 29974 2082 30000
rect 2036 29959 2082 29974
rect 2194 29974 2200 30008
rect 2234 29974 2240 30008
rect 2328 30061 2358 30070
rect 2392 30070 2398 30080
rect 2510 30224 2556 30262
rect 2648 30301 2738 30310
rect 2648 30249 2667 30301
rect 2719 30249 2738 30301
rect 2648 30240 2738 30249
rect 2826 30296 2872 30334
rect 2984 30584 3030 30622
rect 3118 30671 3208 30680
rect 3118 30619 3137 30671
rect 3189 30619 3208 30671
rect 3118 30610 3208 30619
rect 3258 30620 3338 31000
rect 4148 30782 4293 31896
rect 4687 30782 4698 31896
rect 4148 30620 4698 30782
rect 2984 30550 2990 30584
rect 3024 30550 3030 30584
rect 2984 30512 3030 30550
rect 2984 30478 2990 30512
rect 3024 30478 3030 30512
rect 2984 30440 3030 30478
rect 2984 30406 2990 30440
rect 3024 30406 3030 30440
rect 2984 30368 3030 30406
rect 2984 30334 2990 30368
rect 3024 30334 3030 30368
rect 2984 30310 3030 30334
rect 3142 30584 3188 30610
rect 3142 30550 3148 30584
rect 3182 30550 3188 30584
rect 3142 30512 3188 30550
rect 3142 30478 3148 30512
rect 3182 30478 3188 30512
rect 3142 30440 3188 30478
rect 3142 30406 3148 30440
rect 3182 30406 3188 30440
rect 3142 30368 3188 30406
rect 3142 30334 3148 30368
rect 3182 30334 3188 30368
rect 2826 30262 2832 30296
rect 2866 30262 2872 30296
rect 2510 30190 2516 30224
rect 2550 30190 2556 30224
rect 2510 30152 2556 30190
rect 2510 30118 2516 30152
rect 2550 30118 2556 30152
rect 2510 30080 2556 30118
rect 2392 30061 2418 30070
rect 2328 30009 2347 30061
rect 2399 30009 2418 30061
rect 2328 30008 2418 30009
rect 2328 30000 2358 30008
rect 2194 29959 2240 29974
rect 2352 29974 2358 30000
rect 2392 30000 2418 30008
rect 2510 30046 2516 30080
rect 2550 30046 2556 30080
rect 2668 30224 2714 30240
rect 2668 30190 2674 30224
rect 2708 30190 2714 30224
rect 2668 30152 2714 30190
rect 2668 30118 2674 30152
rect 2708 30118 2714 30152
rect 2668 30080 2714 30118
rect 2668 30070 2674 30080
rect 2510 30008 2556 30046
rect 2392 29974 2398 30000
rect 2352 29959 2398 29974
rect 2510 29974 2516 30008
rect 2550 29974 2556 30008
rect 2648 30061 2674 30070
rect 2708 30070 2714 30080
rect 2826 30224 2872 30262
rect 2968 30301 3058 30310
rect 2968 30249 2987 30301
rect 3039 30249 3058 30301
rect 2968 30240 3058 30249
rect 3142 30296 3188 30334
rect 3142 30262 3148 30296
rect 3182 30262 3188 30296
rect 2826 30190 2832 30224
rect 2866 30190 2872 30224
rect 2826 30152 2872 30190
rect 2826 30118 2832 30152
rect 2866 30118 2872 30152
rect 2826 30080 2872 30118
rect 2708 30061 2738 30070
rect 2648 30009 2667 30061
rect 2719 30009 2738 30061
rect 2648 30008 2738 30009
rect 2648 30000 2674 30008
rect 2510 29959 2556 29974
rect 2668 29974 2674 30000
rect 2708 30000 2738 30008
rect 2826 30046 2832 30080
rect 2866 30046 2872 30080
rect 2984 30224 3030 30240
rect 2984 30190 2990 30224
rect 3024 30190 3030 30224
rect 2984 30152 3030 30190
rect 2984 30118 2990 30152
rect 3024 30118 3030 30152
rect 2984 30080 3030 30118
rect 2984 30070 2990 30080
rect 2826 30008 2872 30046
rect 2708 29974 2714 30000
rect 2668 29959 2714 29974
rect 2826 29974 2832 30008
rect 2866 29974 2872 30008
rect 2968 30061 2990 30070
rect 3024 30070 3030 30080
rect 3142 30224 3188 30262
rect 3142 30190 3148 30224
rect 3182 30190 3188 30224
rect 3142 30152 3188 30190
rect 3142 30118 3148 30152
rect 3182 30118 3188 30152
rect 3142 30080 3188 30118
rect 3024 30061 3058 30070
rect 2968 30009 2987 30061
rect 3039 30009 3058 30061
rect 2968 30008 3058 30009
rect 2968 30000 2990 30008
rect 2826 29959 2872 29974
rect 2984 29974 2990 30000
rect 3024 30000 3058 30008
rect 3142 30046 3148 30080
rect 3182 30046 3188 30080
rect 3142 30008 3188 30046
rect 3024 29974 3030 30000
rect 2984 29959 3030 29974
rect 3142 29974 3148 30008
rect 3182 29974 3188 30008
rect 3142 29959 3188 29974
rect 3258 30416 4698 30620
rect 3258 30330 4293 30416
rect 3258 29920 3338 30330
rect -3322 29912 3338 29920
rect -3322 29878 -3093 29912
rect -3059 29878 -2935 29912
rect -2901 29878 -2777 29912
rect -2743 29878 -2619 29912
rect -2585 29878 -2461 29912
rect -2427 29878 -2303 29912
rect -2269 29878 -2145 29912
rect -2111 29886 -1987 29912
rect -2111 29878 -2058 29886
rect -3322 29870 -2058 29878
rect -2112 29834 -2058 29870
rect -2006 29878 -1987 29886
rect -1953 29878 -1829 29912
rect -1795 29878 -1671 29912
rect -1637 29878 -1513 29912
rect -1479 29878 -1355 29912
rect -1321 29878 -1197 29912
rect -1163 29878 -1039 29912
rect -1005 29878 -881 29912
rect -847 29878 -723 29912
rect -689 29878 -565 29912
rect -531 29878 -407 29912
rect -373 29878 -249 29912
rect -215 29878 -91 29912
rect -57 29878 67 29912
rect 101 29878 225 29912
rect 259 29878 383 29912
rect 417 29878 541 29912
rect 575 29878 699 29912
rect 733 29878 857 29912
rect 891 29878 1015 29912
rect 1049 29878 1173 29912
rect 1207 29878 1331 29912
rect 1365 29878 1489 29912
rect 1523 29878 1647 29912
rect 1681 29878 1805 29912
rect 1839 29878 1963 29912
rect 1997 29886 2121 29912
rect 1997 29878 2002 29886
rect -2006 29870 2002 29878
rect -2006 29834 -1952 29870
rect -2112 29810 -1952 29834
rect 1948 29834 2002 29870
rect 2054 29878 2121 29886
rect 2155 29878 2279 29912
rect 2313 29878 2437 29912
rect 2471 29878 2595 29912
rect 2629 29878 2753 29912
rect 2787 29878 2911 29912
rect 2945 29878 3069 29912
rect 3103 29878 3338 29912
rect 2054 29870 3338 29878
rect 2054 29834 2108 29870
rect -892 29816 898 29820
rect -1635 29810 1645 29816
rect 1948 29810 2108 29834
rect -1635 29776 -1596 29810
rect -1562 29776 -1524 29810
rect -1490 29776 -1452 29810
rect -1418 29776 -1380 29810
rect -1346 29776 -1308 29810
rect -1274 29776 -1236 29810
rect -1202 29776 -1164 29810
rect -1130 29776 -1092 29810
rect -1058 29776 -1020 29810
rect -986 29776 -948 29810
rect -914 29776 -876 29810
rect -842 29776 -804 29810
rect -770 29776 -732 29810
rect -698 29776 -660 29810
rect -626 29776 -588 29810
rect -554 29776 -516 29810
rect -482 29776 -444 29810
rect -410 29776 -372 29810
rect -338 29776 -300 29810
rect -266 29776 -228 29810
rect -194 29776 -156 29810
rect -122 29776 -84 29810
rect -50 29776 -12 29810
rect 22 29776 60 29810
rect 94 29776 132 29810
rect 166 29776 204 29810
rect 238 29776 276 29810
rect 310 29776 348 29810
rect 382 29776 420 29810
rect 454 29776 492 29810
rect 526 29776 564 29810
rect 598 29776 636 29810
rect 670 29776 708 29810
rect 742 29776 780 29810
rect 814 29776 852 29810
rect 886 29776 924 29810
rect 958 29776 996 29810
rect 1030 29776 1068 29810
rect 1102 29776 1140 29810
rect 1174 29776 1212 29810
rect 1246 29776 1284 29810
rect 1318 29776 1356 29810
rect 1390 29776 1428 29810
rect 1462 29776 1500 29810
rect 1534 29776 1572 29810
rect 1606 29776 1645 29810
rect -1635 29770 1645 29776
rect -892 29747 898 29770
rect -892 29503 -629 29747
rect -385 29503 421 29747
rect 665 29503 898 29747
rect -892 29472 898 29503
rect -892 29438 -841 29472
rect -807 29438 -769 29472
rect -735 29438 -697 29472
rect -663 29438 -625 29472
rect -591 29438 -553 29472
rect -519 29438 -481 29472
rect -447 29438 -409 29472
rect -375 29438 -337 29472
rect -303 29438 -265 29472
rect -231 29438 -193 29472
rect -159 29438 -121 29472
rect -87 29438 -49 29472
rect -15 29438 23 29472
rect 57 29438 95 29472
rect 129 29438 167 29472
rect 201 29438 239 29472
rect 273 29438 311 29472
rect 345 29438 383 29472
rect 417 29438 455 29472
rect 489 29438 527 29472
rect 561 29438 599 29472
rect 633 29438 671 29472
rect 705 29438 743 29472
rect 777 29438 815 29472
rect 849 29438 898 29472
rect -892 29430 898 29438
rect -4710 29300 -4270 29312
rect -1822 29370 1828 29380
rect -1822 29336 -1593 29370
rect -1559 29336 -1435 29370
rect -1401 29336 -1277 29370
rect -1243 29336 -1119 29370
rect -1085 29336 -961 29370
rect -927 29336 -803 29370
rect -769 29336 -645 29370
rect -611 29336 -487 29370
rect -453 29336 -329 29370
rect -295 29336 -171 29370
rect -137 29336 -13 29370
rect 21 29336 145 29370
rect 179 29336 303 29370
rect 337 29336 461 29370
rect 495 29336 619 29370
rect 653 29336 777 29370
rect 811 29336 935 29370
rect 969 29336 1093 29370
rect 1127 29336 1251 29370
rect 1285 29336 1409 29370
rect 1443 29336 1567 29370
rect 1601 29336 1828 29370
rect -1822 29330 1828 29336
rect -6370 29190 -5440 29200
rect -6370 29140 -6350 29190
rect -6190 29140 -6000 29190
rect -5840 29140 -5630 29190
rect -5470 29140 -5440 29190
rect -6370 21760 -5440 29140
rect -1822 28250 -1742 29330
rect -1678 29274 -1632 29289
rect -1678 29250 -1672 29274
rect -1702 29241 -1672 29250
rect -1638 29250 -1632 29274
rect -1520 29274 -1474 29289
rect -1638 29241 -1612 29250
rect -1702 29189 -1683 29241
rect -1631 29189 -1612 29241
rect -1702 29180 -1672 29189
rect -1678 29168 -1672 29180
rect -1638 29180 -1612 29189
rect -1520 29240 -1514 29274
rect -1480 29240 -1474 29274
rect -1362 29274 -1316 29289
rect -1362 29250 -1356 29274
rect -1520 29202 -1474 29240
rect -1638 29168 -1632 29180
rect -1678 29130 -1632 29168
rect -1678 29096 -1672 29130
rect -1638 29096 -1632 29130
rect -1678 29058 -1632 29096
rect -1678 29040 -1672 29058
rect -1702 29031 -1672 29040
rect -1638 29040 -1632 29058
rect -1520 29168 -1514 29202
rect -1480 29168 -1474 29202
rect -1382 29241 -1356 29250
rect -1322 29250 -1316 29274
rect -1204 29274 -1158 29289
rect -1322 29241 -1292 29250
rect -1382 29189 -1363 29241
rect -1311 29189 -1292 29241
rect -1382 29180 -1356 29189
rect -1520 29130 -1474 29168
rect -1520 29096 -1514 29130
rect -1480 29096 -1474 29130
rect -1520 29058 -1474 29096
rect -1638 29031 -1612 29040
rect -1702 28979 -1683 29031
rect -1631 28979 -1612 29031
rect -1702 28970 -1672 28979
rect -1678 28952 -1672 28970
rect -1638 28970 -1612 28979
rect -1520 29024 -1514 29058
rect -1480 29024 -1474 29058
rect -1362 29168 -1356 29180
rect -1322 29180 -1292 29189
rect -1204 29240 -1198 29274
rect -1164 29240 -1158 29274
rect -1046 29274 -1000 29289
rect -1046 29250 -1040 29274
rect -1204 29202 -1158 29240
rect -1322 29168 -1316 29180
rect -1362 29130 -1316 29168
rect -1362 29096 -1356 29130
rect -1322 29096 -1316 29130
rect -1362 29058 -1316 29096
rect -1362 29040 -1356 29058
rect -1520 28986 -1474 29024
rect -1638 28952 -1632 28970
rect -1678 28914 -1632 28952
rect -1678 28880 -1672 28914
rect -1638 28880 -1632 28914
rect -1678 28842 -1632 28880
rect -1678 28808 -1672 28842
rect -1638 28808 -1632 28842
rect -1678 28770 -1632 28808
rect -1678 28736 -1672 28770
rect -1638 28736 -1632 28770
rect -1678 28698 -1632 28736
rect -1678 28664 -1672 28698
rect -1638 28664 -1632 28698
rect -1678 28626 -1632 28664
rect -1678 28592 -1672 28626
rect -1638 28592 -1632 28626
rect -1520 28952 -1514 28986
rect -1480 28952 -1474 28986
rect -1382 29031 -1356 29040
rect -1322 29040 -1316 29058
rect -1204 29168 -1198 29202
rect -1164 29168 -1158 29202
rect -1072 29241 -1040 29250
rect -1006 29250 -1000 29274
rect -888 29274 -842 29289
rect -1006 29241 -982 29250
rect -1072 29189 -1053 29241
rect -1001 29189 -982 29241
rect -1072 29180 -1040 29189
rect -1204 29130 -1158 29168
rect -1204 29096 -1198 29130
rect -1164 29096 -1158 29130
rect -1204 29058 -1158 29096
rect -1322 29031 -1292 29040
rect -1382 28979 -1363 29031
rect -1311 28979 -1292 29031
rect -1382 28970 -1356 28979
rect -1520 28914 -1474 28952
rect -1520 28880 -1514 28914
rect -1480 28880 -1474 28914
rect -1520 28842 -1474 28880
rect -1520 28808 -1514 28842
rect -1480 28808 -1474 28842
rect -1520 28770 -1474 28808
rect -1520 28736 -1514 28770
rect -1480 28736 -1474 28770
rect -1520 28698 -1474 28736
rect -1520 28664 -1514 28698
rect -1480 28664 -1474 28698
rect -1520 28626 -1474 28664
rect -1520 28610 -1514 28626
rect -1678 28554 -1632 28592
rect -1678 28520 -1672 28554
rect -1638 28520 -1632 28554
rect -1542 28601 -1514 28610
rect -1480 28610 -1474 28626
rect -1362 28952 -1356 28970
rect -1322 28970 -1292 28979
rect -1204 29024 -1198 29058
rect -1164 29024 -1158 29058
rect -1046 29168 -1040 29180
rect -1006 29180 -982 29189
rect -888 29240 -882 29274
rect -848 29240 -842 29274
rect -730 29274 -684 29289
rect -730 29250 -724 29274
rect -888 29202 -842 29240
rect -1006 29168 -1000 29180
rect -1046 29130 -1000 29168
rect -1046 29096 -1040 29130
rect -1006 29096 -1000 29130
rect -1046 29058 -1000 29096
rect -1046 29040 -1040 29058
rect -1204 28986 -1158 29024
rect -1322 28952 -1316 28970
rect -1362 28914 -1316 28952
rect -1362 28880 -1356 28914
rect -1322 28880 -1316 28914
rect -1362 28842 -1316 28880
rect -1362 28808 -1356 28842
rect -1322 28808 -1316 28842
rect -1362 28770 -1316 28808
rect -1362 28736 -1356 28770
rect -1322 28736 -1316 28770
rect -1362 28698 -1316 28736
rect -1362 28664 -1356 28698
rect -1322 28664 -1316 28698
rect -1362 28626 -1316 28664
rect -1480 28601 -1452 28610
rect -1542 28549 -1523 28601
rect -1471 28549 -1452 28601
rect -1542 28540 -1514 28549
rect -1678 28482 -1632 28520
rect -1678 28448 -1672 28482
rect -1638 28448 -1632 28482
rect -1678 28410 -1632 28448
rect -1678 28376 -1672 28410
rect -1638 28376 -1632 28410
rect -1520 28520 -1514 28540
rect -1480 28540 -1452 28549
rect -1362 28592 -1356 28626
rect -1322 28592 -1316 28626
rect -1204 28952 -1198 28986
rect -1164 28952 -1158 28986
rect -1072 29031 -1040 29040
rect -1006 29040 -1000 29058
rect -888 29168 -882 29202
rect -848 29168 -842 29202
rect -752 29241 -724 29250
rect -690 29250 -684 29274
rect -572 29274 -526 29289
rect -690 29241 -662 29250
rect -752 29189 -733 29241
rect -681 29189 -662 29241
rect -752 29180 -724 29189
rect -888 29130 -842 29168
rect -888 29096 -882 29130
rect -848 29096 -842 29130
rect -888 29058 -842 29096
rect -1006 29031 -982 29040
rect -1072 28979 -1053 29031
rect -1001 28979 -982 29031
rect -1072 28970 -1040 28979
rect -1204 28914 -1158 28952
rect -1204 28880 -1198 28914
rect -1164 28880 -1158 28914
rect -1204 28842 -1158 28880
rect -1204 28808 -1198 28842
rect -1164 28808 -1158 28842
rect -1204 28770 -1158 28808
rect -1204 28736 -1198 28770
rect -1164 28736 -1158 28770
rect -1204 28698 -1158 28736
rect -1204 28664 -1198 28698
rect -1164 28664 -1158 28698
rect -1204 28626 -1158 28664
rect -1204 28610 -1198 28626
rect -1362 28554 -1316 28592
rect -1480 28520 -1474 28540
rect -1520 28482 -1474 28520
rect -1520 28448 -1514 28482
rect -1480 28448 -1474 28482
rect -1520 28410 -1474 28448
rect -1520 28400 -1514 28410
rect -1678 28338 -1632 28376
rect -1678 28304 -1672 28338
rect -1638 28304 -1632 28338
rect -1542 28391 -1514 28400
rect -1480 28400 -1474 28410
rect -1362 28520 -1356 28554
rect -1322 28520 -1316 28554
rect -1222 28601 -1198 28610
rect -1164 28610 -1158 28626
rect -1046 28952 -1040 28970
rect -1006 28970 -982 28979
rect -888 29024 -882 29058
rect -848 29024 -842 29058
rect -730 29168 -724 29180
rect -690 29180 -662 29189
rect -572 29240 -566 29274
rect -532 29240 -526 29274
rect -414 29274 -368 29289
rect -414 29250 -408 29274
rect -572 29202 -526 29240
rect -690 29168 -684 29180
rect -730 29130 -684 29168
rect -730 29096 -724 29130
rect -690 29096 -684 29130
rect -730 29058 -684 29096
rect -730 29040 -724 29058
rect -888 28986 -842 29024
rect -1006 28952 -1000 28970
rect -1046 28914 -1000 28952
rect -1046 28880 -1040 28914
rect -1006 28880 -1000 28914
rect -1046 28842 -1000 28880
rect -1046 28808 -1040 28842
rect -1006 28808 -1000 28842
rect -1046 28770 -1000 28808
rect -1046 28736 -1040 28770
rect -1006 28736 -1000 28770
rect -1046 28698 -1000 28736
rect -1046 28664 -1040 28698
rect -1006 28664 -1000 28698
rect -1046 28626 -1000 28664
rect -1164 28601 -1132 28610
rect -1222 28549 -1203 28601
rect -1151 28549 -1132 28601
rect -1222 28540 -1198 28549
rect -1362 28482 -1316 28520
rect -1362 28448 -1356 28482
rect -1322 28448 -1316 28482
rect -1362 28410 -1316 28448
rect -1480 28391 -1452 28400
rect -1542 28339 -1523 28391
rect -1471 28339 -1452 28391
rect -1542 28338 -1452 28339
rect -1542 28330 -1514 28338
rect -1678 28289 -1632 28304
rect -1520 28304 -1514 28330
rect -1480 28330 -1452 28338
rect -1362 28376 -1356 28410
rect -1322 28376 -1316 28410
rect -1204 28520 -1198 28540
rect -1164 28540 -1132 28549
rect -1046 28592 -1040 28626
rect -1006 28592 -1000 28626
rect -888 28952 -882 28986
rect -848 28952 -842 28986
rect -752 29031 -724 29040
rect -690 29040 -684 29058
rect -572 29168 -566 29202
rect -532 29168 -526 29202
rect -432 29241 -408 29250
rect -374 29250 -368 29274
rect -256 29274 -210 29289
rect -374 29241 -342 29250
rect -432 29189 -413 29241
rect -361 29189 -342 29241
rect -432 29180 -408 29189
rect -572 29130 -526 29168
rect -572 29096 -566 29130
rect -532 29096 -526 29130
rect -572 29058 -526 29096
rect -690 29031 -662 29040
rect -752 28979 -733 29031
rect -681 28979 -662 29031
rect -752 28970 -724 28979
rect -888 28914 -842 28952
rect -888 28880 -882 28914
rect -848 28880 -842 28914
rect -888 28842 -842 28880
rect -888 28808 -882 28842
rect -848 28808 -842 28842
rect -888 28770 -842 28808
rect -888 28736 -882 28770
rect -848 28736 -842 28770
rect -888 28698 -842 28736
rect -888 28664 -882 28698
rect -848 28664 -842 28698
rect -888 28626 -842 28664
rect -888 28610 -882 28626
rect -1046 28554 -1000 28592
rect -1164 28520 -1158 28540
rect -1204 28482 -1158 28520
rect -1204 28448 -1198 28482
rect -1164 28448 -1158 28482
rect -1204 28410 -1158 28448
rect -1204 28400 -1198 28410
rect -1362 28338 -1316 28376
rect -1480 28304 -1474 28330
rect -1520 28289 -1474 28304
rect -1362 28304 -1356 28338
rect -1322 28304 -1316 28338
rect -1222 28391 -1198 28400
rect -1164 28400 -1158 28410
rect -1046 28520 -1040 28554
rect -1006 28520 -1000 28554
rect -912 28601 -882 28610
rect -848 28610 -842 28626
rect -730 28952 -724 28970
rect -690 28970 -662 28979
rect -572 29024 -566 29058
rect -532 29024 -526 29058
rect -414 29168 -408 29180
rect -374 29180 -342 29189
rect -256 29240 -250 29274
rect -216 29240 -210 29274
rect -98 29274 -52 29289
rect -98 29250 -92 29274
rect -256 29202 -210 29240
rect -374 29168 -368 29180
rect -414 29130 -368 29168
rect -414 29096 -408 29130
rect -374 29096 -368 29130
rect -414 29058 -368 29096
rect -414 29040 -408 29058
rect -572 28986 -526 29024
rect -690 28952 -684 28970
rect -730 28914 -684 28952
rect -730 28880 -724 28914
rect -690 28880 -684 28914
rect -730 28842 -684 28880
rect -730 28808 -724 28842
rect -690 28808 -684 28842
rect -730 28770 -684 28808
rect -730 28736 -724 28770
rect -690 28736 -684 28770
rect -730 28698 -684 28736
rect -730 28664 -724 28698
rect -690 28664 -684 28698
rect -730 28626 -684 28664
rect -848 28601 -822 28610
rect -912 28549 -893 28601
rect -841 28549 -822 28601
rect -912 28540 -882 28549
rect -1046 28482 -1000 28520
rect -1046 28448 -1040 28482
rect -1006 28448 -1000 28482
rect -1046 28410 -1000 28448
rect -1164 28391 -1132 28400
rect -1222 28339 -1203 28391
rect -1151 28339 -1132 28391
rect -1222 28338 -1132 28339
rect -1222 28330 -1198 28338
rect -1362 28289 -1316 28304
rect -1204 28304 -1198 28330
rect -1164 28330 -1132 28338
rect -1046 28376 -1040 28410
rect -1006 28376 -1000 28410
rect -888 28520 -882 28540
rect -848 28540 -822 28549
rect -730 28592 -724 28626
rect -690 28592 -684 28626
rect -572 28952 -566 28986
rect -532 28952 -526 28986
rect -432 29031 -408 29040
rect -374 29040 -368 29058
rect -256 29168 -250 29202
rect -216 29168 -210 29202
rect -122 29241 -92 29250
rect -58 29250 -52 29274
rect 60 29274 106 29289
rect -58 29241 -32 29250
rect -122 29189 -103 29241
rect -51 29189 -32 29241
rect -122 29180 -92 29189
rect -256 29130 -210 29168
rect -256 29096 -250 29130
rect -216 29096 -210 29130
rect -256 29058 -210 29096
rect -374 29031 -342 29040
rect -432 28979 -413 29031
rect -361 28979 -342 29031
rect -432 28970 -408 28979
rect -572 28914 -526 28952
rect -572 28880 -566 28914
rect -532 28880 -526 28914
rect -572 28842 -526 28880
rect -572 28808 -566 28842
rect -532 28808 -526 28842
rect -572 28770 -526 28808
rect -572 28736 -566 28770
rect -532 28736 -526 28770
rect -572 28698 -526 28736
rect -572 28664 -566 28698
rect -532 28664 -526 28698
rect -572 28626 -526 28664
rect -572 28610 -566 28626
rect -730 28554 -684 28592
rect -848 28520 -842 28540
rect -888 28482 -842 28520
rect -888 28448 -882 28482
rect -848 28448 -842 28482
rect -888 28410 -842 28448
rect -888 28400 -882 28410
rect -1046 28338 -1000 28376
rect -1164 28304 -1158 28330
rect -1204 28289 -1158 28304
rect -1046 28304 -1040 28338
rect -1006 28304 -1000 28338
rect -912 28391 -882 28400
rect -848 28400 -842 28410
rect -730 28520 -724 28554
rect -690 28520 -684 28554
rect -592 28601 -566 28610
rect -532 28610 -526 28626
rect -414 28952 -408 28970
rect -374 28970 -342 28979
rect -256 29024 -250 29058
rect -216 29024 -210 29058
rect -98 29168 -92 29180
rect -58 29180 -32 29189
rect 60 29240 66 29274
rect 100 29240 106 29274
rect 218 29274 264 29289
rect 218 29250 224 29274
rect 60 29202 106 29240
rect -58 29168 -52 29180
rect -98 29130 -52 29168
rect -98 29096 -92 29130
rect -58 29096 -52 29130
rect -98 29058 -52 29096
rect -98 29040 -92 29058
rect -256 28986 -210 29024
rect -374 28952 -368 28970
rect -414 28914 -368 28952
rect -414 28880 -408 28914
rect -374 28880 -368 28914
rect -414 28842 -368 28880
rect -414 28808 -408 28842
rect -374 28808 -368 28842
rect -414 28770 -368 28808
rect -414 28736 -408 28770
rect -374 28736 -368 28770
rect -414 28698 -368 28736
rect -414 28664 -408 28698
rect -374 28664 -368 28698
rect -414 28626 -368 28664
rect -532 28601 -502 28610
rect -592 28549 -573 28601
rect -521 28549 -502 28601
rect -592 28540 -566 28549
rect -730 28482 -684 28520
rect -730 28448 -724 28482
rect -690 28448 -684 28482
rect -730 28410 -684 28448
rect -848 28391 -822 28400
rect -912 28339 -893 28391
rect -841 28339 -822 28391
rect -912 28338 -822 28339
rect -912 28330 -882 28338
rect -1046 28289 -1000 28304
rect -888 28304 -882 28330
rect -848 28330 -822 28338
rect -730 28376 -724 28410
rect -690 28376 -684 28410
rect -572 28520 -566 28540
rect -532 28540 -502 28549
rect -414 28592 -408 28626
rect -374 28592 -368 28626
rect -256 28952 -250 28986
rect -216 28952 -210 28986
rect -122 29031 -92 29040
rect -58 29040 -52 29058
rect 60 29168 66 29202
rect 100 29168 106 29202
rect 198 29241 224 29250
rect 258 29250 264 29274
rect 376 29274 422 29289
rect 258 29241 288 29250
rect 198 29189 217 29241
rect 269 29189 288 29241
rect 198 29180 224 29189
rect 60 29130 106 29168
rect 60 29096 66 29130
rect 100 29096 106 29130
rect 60 29058 106 29096
rect -58 29031 -32 29040
rect -122 28979 -103 29031
rect -51 28979 -32 29031
rect -122 28970 -92 28979
rect -256 28914 -210 28952
rect -256 28880 -250 28914
rect -216 28880 -210 28914
rect -256 28842 -210 28880
rect -256 28808 -250 28842
rect -216 28808 -210 28842
rect -256 28770 -210 28808
rect -256 28736 -250 28770
rect -216 28736 -210 28770
rect -256 28698 -210 28736
rect -256 28664 -250 28698
rect -216 28664 -210 28698
rect -256 28626 -210 28664
rect -256 28610 -250 28626
rect -414 28554 -368 28592
rect -532 28520 -526 28540
rect -572 28482 -526 28520
rect -572 28448 -566 28482
rect -532 28448 -526 28482
rect -572 28410 -526 28448
rect -572 28400 -566 28410
rect -730 28338 -684 28376
rect -848 28304 -842 28330
rect -888 28289 -842 28304
rect -730 28304 -724 28338
rect -690 28304 -684 28338
rect -592 28391 -566 28400
rect -532 28400 -526 28410
rect -414 28520 -408 28554
rect -374 28520 -368 28554
rect -272 28601 -250 28610
rect -216 28610 -210 28626
rect -98 28952 -92 28970
rect -58 28970 -32 28979
rect 60 29024 66 29058
rect 100 29024 106 29058
rect 218 29168 224 29180
rect 258 29180 288 29189
rect 376 29240 382 29274
rect 416 29240 422 29274
rect 534 29274 580 29289
rect 534 29250 540 29274
rect 376 29202 422 29240
rect 258 29168 264 29180
rect 218 29130 264 29168
rect 218 29096 224 29130
rect 258 29096 264 29130
rect 218 29058 264 29096
rect 218 29040 224 29058
rect 60 28986 106 29024
rect -58 28952 -52 28970
rect -98 28914 -52 28952
rect -98 28880 -92 28914
rect -58 28880 -52 28914
rect -98 28842 -52 28880
rect -98 28808 -92 28842
rect -58 28808 -52 28842
rect -98 28770 -52 28808
rect -98 28736 -92 28770
rect -58 28736 -52 28770
rect -98 28698 -52 28736
rect -98 28664 -92 28698
rect -58 28664 -52 28698
rect -98 28626 -52 28664
rect -216 28601 -182 28610
rect -272 28549 -253 28601
rect -201 28549 -182 28601
rect -272 28540 -250 28549
rect -414 28482 -368 28520
rect -414 28448 -408 28482
rect -374 28448 -368 28482
rect -414 28410 -368 28448
rect -532 28391 -502 28400
rect -592 28339 -573 28391
rect -521 28339 -502 28391
rect -592 28338 -502 28339
rect -592 28330 -566 28338
rect -730 28289 -684 28304
rect -572 28304 -566 28330
rect -532 28330 -502 28338
rect -414 28376 -408 28410
rect -374 28376 -368 28410
rect -256 28520 -250 28540
rect -216 28540 -182 28549
rect -98 28592 -92 28626
rect -58 28592 -52 28626
rect 60 28952 66 28986
rect 100 28952 106 28986
rect 198 29031 224 29040
rect 258 29040 264 29058
rect 376 29168 382 29202
rect 416 29168 422 29202
rect 518 29241 540 29250
rect 574 29250 580 29274
rect 692 29274 738 29289
rect 574 29241 608 29250
rect 518 29189 537 29241
rect 589 29189 608 29241
rect 518 29180 540 29189
rect 376 29130 422 29168
rect 376 29096 382 29130
rect 416 29096 422 29130
rect 376 29058 422 29096
rect 258 29031 288 29040
rect 198 28979 217 29031
rect 269 28979 288 29031
rect 198 28970 224 28979
rect 60 28914 106 28952
rect 60 28880 66 28914
rect 100 28880 106 28914
rect 60 28842 106 28880
rect 60 28808 66 28842
rect 100 28808 106 28842
rect 60 28770 106 28808
rect 60 28736 66 28770
rect 100 28736 106 28770
rect 60 28698 106 28736
rect 60 28664 66 28698
rect 100 28664 106 28698
rect 60 28626 106 28664
rect 60 28610 66 28626
rect -98 28554 -52 28592
rect -216 28520 -210 28540
rect -256 28482 -210 28520
rect -256 28448 -250 28482
rect -216 28448 -210 28482
rect -256 28410 -210 28448
rect -256 28400 -250 28410
rect -414 28338 -368 28376
rect -532 28304 -526 28330
rect -572 28289 -526 28304
rect -414 28304 -408 28338
rect -374 28304 -368 28338
rect -272 28391 -250 28400
rect -216 28400 -210 28410
rect -98 28520 -92 28554
rect -58 28520 -52 28554
rect 38 28601 66 28610
rect 100 28610 106 28626
rect 218 28952 224 28970
rect 258 28970 288 28979
rect 376 29024 382 29058
rect 416 29024 422 29058
rect 534 29168 540 29180
rect 574 29180 608 29189
rect 692 29240 698 29274
rect 732 29240 738 29274
rect 850 29274 896 29289
rect 850 29250 856 29274
rect 692 29202 738 29240
rect 574 29168 580 29180
rect 534 29130 580 29168
rect 534 29096 540 29130
rect 574 29096 580 29130
rect 534 29058 580 29096
rect 534 29040 540 29058
rect 376 28986 422 29024
rect 258 28952 264 28970
rect 218 28914 264 28952
rect 218 28880 224 28914
rect 258 28880 264 28914
rect 218 28842 264 28880
rect 218 28808 224 28842
rect 258 28808 264 28842
rect 218 28770 264 28808
rect 218 28736 224 28770
rect 258 28736 264 28770
rect 218 28698 264 28736
rect 218 28664 224 28698
rect 258 28664 264 28698
rect 218 28626 264 28664
rect 100 28601 128 28610
rect 38 28549 57 28601
rect 109 28549 128 28601
rect 38 28540 66 28549
rect -98 28482 -52 28520
rect -98 28448 -92 28482
rect -58 28448 -52 28482
rect -98 28410 -52 28448
rect -216 28391 -182 28400
rect -272 28339 -253 28391
rect -201 28339 -182 28391
rect -272 28338 -182 28339
rect -272 28330 -250 28338
rect -414 28289 -368 28304
rect -256 28304 -250 28330
rect -216 28330 -182 28338
rect -98 28376 -92 28410
rect -58 28376 -52 28410
rect 60 28520 66 28540
rect 100 28540 128 28549
rect 218 28592 224 28626
rect 258 28592 264 28626
rect 376 28952 382 28986
rect 416 28952 422 28986
rect 518 29031 540 29040
rect 574 29040 580 29058
rect 692 29168 698 29202
rect 732 29168 738 29202
rect 828 29241 856 29250
rect 890 29250 896 29274
rect 1008 29274 1054 29289
rect 890 29241 918 29250
rect 828 29189 847 29241
rect 899 29189 918 29241
rect 828 29180 856 29189
rect 692 29130 738 29168
rect 692 29096 698 29130
rect 732 29096 738 29130
rect 692 29058 738 29096
rect 574 29031 608 29040
rect 518 28979 537 29031
rect 589 28979 608 29031
rect 518 28970 540 28979
rect 376 28914 422 28952
rect 376 28880 382 28914
rect 416 28880 422 28914
rect 376 28842 422 28880
rect 376 28808 382 28842
rect 416 28808 422 28842
rect 376 28770 422 28808
rect 376 28736 382 28770
rect 416 28736 422 28770
rect 376 28698 422 28736
rect 376 28664 382 28698
rect 416 28664 422 28698
rect 376 28626 422 28664
rect 376 28610 382 28626
rect 218 28554 264 28592
rect 100 28520 106 28540
rect 60 28482 106 28520
rect 60 28448 66 28482
rect 100 28448 106 28482
rect 60 28410 106 28448
rect 60 28400 66 28410
rect -98 28338 -52 28376
rect -216 28304 -210 28330
rect -256 28289 -210 28304
rect -98 28304 -92 28338
rect -58 28304 -52 28338
rect 38 28391 66 28400
rect 100 28400 106 28410
rect 218 28520 224 28554
rect 258 28520 264 28554
rect 358 28601 382 28610
rect 416 28610 422 28626
rect 534 28952 540 28970
rect 574 28970 608 28979
rect 692 29024 698 29058
rect 732 29024 738 29058
rect 850 29168 856 29180
rect 890 29180 918 29189
rect 1008 29240 1014 29274
rect 1048 29240 1054 29274
rect 1166 29274 1212 29289
rect 1166 29250 1172 29274
rect 1008 29202 1054 29240
rect 890 29168 896 29180
rect 850 29130 896 29168
rect 850 29096 856 29130
rect 890 29096 896 29130
rect 850 29058 896 29096
rect 850 29040 856 29058
rect 692 28986 738 29024
rect 574 28952 580 28970
rect 534 28914 580 28952
rect 534 28880 540 28914
rect 574 28880 580 28914
rect 534 28842 580 28880
rect 534 28808 540 28842
rect 574 28808 580 28842
rect 534 28770 580 28808
rect 534 28736 540 28770
rect 574 28736 580 28770
rect 534 28698 580 28736
rect 534 28664 540 28698
rect 574 28664 580 28698
rect 534 28626 580 28664
rect 416 28601 448 28610
rect 358 28549 377 28601
rect 429 28549 448 28601
rect 358 28540 382 28549
rect 218 28482 264 28520
rect 218 28448 224 28482
rect 258 28448 264 28482
rect 218 28410 264 28448
rect 100 28391 128 28400
rect 38 28339 57 28391
rect 109 28339 128 28391
rect 38 28338 128 28339
rect 38 28330 66 28338
rect -98 28289 -52 28304
rect 60 28304 66 28330
rect 100 28330 128 28338
rect 218 28376 224 28410
rect 258 28376 264 28410
rect 376 28520 382 28540
rect 416 28540 448 28549
rect 534 28592 540 28626
rect 574 28592 580 28626
rect 692 28952 698 28986
rect 732 28952 738 28986
rect 828 29031 856 29040
rect 890 29040 896 29058
rect 1008 29168 1014 29202
rect 1048 29168 1054 29202
rect 1148 29241 1172 29250
rect 1206 29250 1212 29274
rect 1324 29274 1370 29289
rect 1206 29241 1238 29250
rect 1148 29189 1167 29241
rect 1219 29189 1238 29241
rect 1148 29180 1172 29189
rect 1008 29130 1054 29168
rect 1008 29096 1014 29130
rect 1048 29096 1054 29130
rect 1008 29058 1054 29096
rect 890 29031 918 29040
rect 828 28979 847 29031
rect 899 28979 918 29031
rect 828 28970 856 28979
rect 692 28914 738 28952
rect 692 28880 698 28914
rect 732 28880 738 28914
rect 692 28842 738 28880
rect 692 28808 698 28842
rect 732 28808 738 28842
rect 692 28770 738 28808
rect 692 28736 698 28770
rect 732 28736 738 28770
rect 692 28698 738 28736
rect 692 28664 698 28698
rect 732 28664 738 28698
rect 692 28626 738 28664
rect 692 28610 698 28626
rect 534 28554 580 28592
rect 416 28520 422 28540
rect 376 28482 422 28520
rect 376 28448 382 28482
rect 416 28448 422 28482
rect 376 28410 422 28448
rect 376 28400 382 28410
rect 218 28338 264 28376
rect 100 28304 106 28330
rect 60 28289 106 28304
rect 218 28304 224 28338
rect 258 28304 264 28338
rect 358 28391 382 28400
rect 416 28400 422 28410
rect 534 28520 540 28554
rect 574 28520 580 28554
rect 668 28601 698 28610
rect 732 28610 738 28626
rect 850 28952 856 28970
rect 890 28970 918 28979
rect 1008 29024 1014 29058
rect 1048 29024 1054 29058
rect 1166 29168 1172 29180
rect 1206 29180 1238 29189
rect 1324 29240 1330 29274
rect 1364 29240 1370 29274
rect 1482 29274 1528 29289
rect 1482 29250 1488 29274
rect 1324 29202 1370 29240
rect 1206 29168 1212 29180
rect 1166 29130 1212 29168
rect 1166 29096 1172 29130
rect 1206 29096 1212 29130
rect 1166 29058 1212 29096
rect 1166 29040 1172 29058
rect 1008 28986 1054 29024
rect 890 28952 896 28970
rect 850 28914 896 28952
rect 850 28880 856 28914
rect 890 28880 896 28914
rect 850 28842 896 28880
rect 850 28808 856 28842
rect 890 28808 896 28842
rect 850 28770 896 28808
rect 850 28736 856 28770
rect 890 28736 896 28770
rect 850 28698 896 28736
rect 850 28664 856 28698
rect 890 28664 896 28698
rect 850 28626 896 28664
rect 732 28601 758 28610
rect 668 28549 687 28601
rect 739 28549 758 28601
rect 668 28540 698 28549
rect 534 28482 580 28520
rect 534 28448 540 28482
rect 574 28448 580 28482
rect 534 28410 580 28448
rect 416 28391 448 28400
rect 358 28339 377 28391
rect 429 28339 448 28391
rect 358 28338 448 28339
rect 358 28330 382 28338
rect 218 28289 264 28304
rect 376 28304 382 28330
rect 416 28330 448 28338
rect 534 28376 540 28410
rect 574 28376 580 28410
rect 692 28520 698 28540
rect 732 28540 758 28549
rect 850 28592 856 28626
rect 890 28592 896 28626
rect 1008 28952 1014 28986
rect 1048 28952 1054 28986
rect 1148 29031 1172 29040
rect 1206 29040 1212 29058
rect 1324 29168 1330 29202
rect 1364 29168 1370 29202
rect 1458 29241 1488 29250
rect 1522 29250 1528 29274
rect 1640 29274 1686 29289
rect 1522 29241 1548 29250
rect 1458 29189 1477 29241
rect 1529 29189 1548 29241
rect 1458 29180 1488 29189
rect 1324 29130 1370 29168
rect 1324 29096 1330 29130
rect 1364 29096 1370 29130
rect 1324 29058 1370 29096
rect 1206 29031 1238 29040
rect 1148 28979 1167 29031
rect 1219 28979 1238 29031
rect 1148 28970 1172 28979
rect 1008 28914 1054 28952
rect 1008 28880 1014 28914
rect 1048 28880 1054 28914
rect 1008 28842 1054 28880
rect 1008 28808 1014 28842
rect 1048 28808 1054 28842
rect 1008 28770 1054 28808
rect 1008 28736 1014 28770
rect 1048 28736 1054 28770
rect 1008 28698 1054 28736
rect 1008 28664 1014 28698
rect 1048 28664 1054 28698
rect 1008 28626 1054 28664
rect 1008 28610 1014 28626
rect 850 28554 896 28592
rect 732 28520 738 28540
rect 692 28482 738 28520
rect 692 28448 698 28482
rect 732 28448 738 28482
rect 692 28410 738 28448
rect 692 28400 698 28410
rect 534 28338 580 28376
rect 416 28304 422 28330
rect 376 28289 422 28304
rect 534 28304 540 28338
rect 574 28304 580 28338
rect 668 28391 698 28400
rect 732 28400 738 28410
rect 850 28520 856 28554
rect 890 28520 896 28554
rect 988 28601 1014 28610
rect 1048 28610 1054 28626
rect 1166 28952 1172 28970
rect 1206 28970 1238 28979
rect 1324 29024 1330 29058
rect 1364 29024 1370 29058
rect 1482 29168 1488 29180
rect 1522 29180 1548 29189
rect 1640 29240 1646 29274
rect 1680 29240 1686 29274
rect 1640 29202 1686 29240
rect 1522 29168 1528 29180
rect 1482 29130 1528 29168
rect 1482 29096 1488 29130
rect 1522 29096 1528 29130
rect 1482 29058 1528 29096
rect 1482 29040 1488 29058
rect 1324 28986 1370 29024
rect 1206 28952 1212 28970
rect 1166 28914 1212 28952
rect 1166 28880 1172 28914
rect 1206 28880 1212 28914
rect 1166 28842 1212 28880
rect 1166 28808 1172 28842
rect 1206 28808 1212 28842
rect 1166 28770 1212 28808
rect 1166 28736 1172 28770
rect 1206 28736 1212 28770
rect 1166 28698 1212 28736
rect 1166 28664 1172 28698
rect 1206 28664 1212 28698
rect 1166 28626 1212 28664
rect 1048 28601 1078 28610
rect 988 28549 1007 28601
rect 1059 28549 1078 28601
rect 988 28540 1014 28549
rect 850 28482 896 28520
rect 850 28448 856 28482
rect 890 28448 896 28482
rect 850 28410 896 28448
rect 732 28391 758 28400
rect 668 28339 687 28391
rect 739 28339 758 28391
rect 668 28338 758 28339
rect 668 28330 698 28338
rect 534 28289 580 28304
rect 692 28304 698 28330
rect 732 28330 758 28338
rect 850 28376 856 28410
rect 890 28376 896 28410
rect 1008 28520 1014 28540
rect 1048 28540 1078 28549
rect 1166 28592 1172 28626
rect 1206 28592 1212 28626
rect 1324 28952 1330 28986
rect 1364 28952 1370 28986
rect 1458 29031 1488 29040
rect 1522 29040 1528 29058
rect 1640 29168 1646 29202
rect 1680 29168 1686 29202
rect 1640 29130 1686 29168
rect 1640 29096 1646 29130
rect 1680 29096 1686 29130
rect 1640 29058 1686 29096
rect 1522 29031 1548 29040
rect 1458 28979 1477 29031
rect 1529 28979 1548 29031
rect 1458 28970 1488 28979
rect 1324 28914 1370 28952
rect 1324 28880 1330 28914
rect 1364 28880 1370 28914
rect 1324 28842 1370 28880
rect 1324 28808 1330 28842
rect 1364 28808 1370 28842
rect 1324 28770 1370 28808
rect 1324 28736 1330 28770
rect 1364 28736 1370 28770
rect 1324 28698 1370 28736
rect 1324 28664 1330 28698
rect 1364 28664 1370 28698
rect 1324 28626 1370 28664
rect 1324 28610 1330 28626
rect 1166 28554 1212 28592
rect 1048 28520 1054 28540
rect 1008 28482 1054 28520
rect 1008 28448 1014 28482
rect 1048 28448 1054 28482
rect 1008 28410 1054 28448
rect 1008 28400 1014 28410
rect 850 28338 896 28376
rect 732 28304 738 28330
rect 692 28289 738 28304
rect 850 28304 856 28338
rect 890 28304 896 28338
rect 988 28391 1014 28400
rect 1048 28400 1054 28410
rect 1166 28520 1172 28554
rect 1206 28520 1212 28554
rect 1308 28601 1330 28610
rect 1364 28610 1370 28626
rect 1482 28952 1488 28970
rect 1522 28970 1548 28979
rect 1640 29024 1646 29058
rect 1680 29024 1686 29058
rect 1640 28986 1686 29024
rect 1522 28952 1528 28970
rect 1482 28914 1528 28952
rect 1482 28880 1488 28914
rect 1522 28880 1528 28914
rect 1482 28842 1528 28880
rect 1482 28808 1488 28842
rect 1522 28808 1528 28842
rect 1482 28770 1528 28808
rect 1482 28736 1488 28770
rect 1522 28736 1528 28770
rect 1482 28698 1528 28736
rect 1482 28664 1488 28698
rect 1522 28664 1528 28698
rect 1482 28626 1528 28664
rect 1364 28601 1398 28610
rect 1308 28549 1327 28601
rect 1379 28549 1398 28601
rect 1308 28540 1330 28549
rect 1166 28482 1212 28520
rect 1166 28448 1172 28482
rect 1206 28448 1212 28482
rect 1166 28410 1212 28448
rect 1048 28391 1078 28400
rect 988 28339 1007 28391
rect 1059 28339 1078 28391
rect 988 28338 1078 28339
rect 988 28330 1014 28338
rect 850 28289 896 28304
rect 1008 28304 1014 28330
rect 1048 28330 1078 28338
rect 1166 28376 1172 28410
rect 1206 28376 1212 28410
rect 1324 28520 1330 28540
rect 1364 28540 1398 28549
rect 1482 28592 1488 28626
rect 1522 28592 1528 28626
rect 1640 28952 1646 28986
rect 1680 28952 1686 28986
rect 1640 28914 1686 28952
rect 1640 28880 1646 28914
rect 1680 28880 1686 28914
rect 1640 28842 1686 28880
rect 1640 28808 1646 28842
rect 1680 28808 1686 28842
rect 1640 28770 1686 28808
rect 1640 28736 1646 28770
rect 1680 28736 1686 28770
rect 1640 28698 1686 28736
rect 1640 28664 1646 28698
rect 1680 28664 1686 28698
rect 1640 28626 1686 28664
rect 1640 28610 1646 28626
rect 1482 28554 1528 28592
rect 1364 28520 1370 28540
rect 1324 28482 1370 28520
rect 1324 28448 1330 28482
rect 1364 28448 1370 28482
rect 1324 28410 1370 28448
rect 1324 28400 1330 28410
rect 1166 28338 1212 28376
rect 1048 28304 1054 28330
rect 1008 28289 1054 28304
rect 1166 28304 1172 28338
rect 1206 28304 1212 28338
rect 1308 28391 1330 28400
rect 1364 28400 1370 28410
rect 1482 28520 1488 28554
rect 1522 28520 1528 28554
rect 1618 28601 1646 28610
rect 1680 28610 1686 28626
rect 1680 28601 1708 28610
rect 1618 28549 1637 28601
rect 1689 28549 1708 28601
rect 1618 28540 1646 28549
rect 1482 28482 1528 28520
rect 1482 28448 1488 28482
rect 1522 28448 1528 28482
rect 1482 28410 1528 28448
rect 1364 28391 1398 28400
rect 1308 28339 1327 28391
rect 1379 28339 1398 28391
rect 1308 28338 1398 28339
rect 1308 28330 1330 28338
rect 1166 28289 1212 28304
rect 1324 28304 1330 28330
rect 1364 28330 1398 28338
rect 1482 28376 1488 28410
rect 1522 28376 1528 28410
rect 1640 28520 1646 28540
rect 1680 28540 1708 28549
rect 1680 28520 1686 28540
rect 1640 28482 1686 28520
rect 1640 28448 1646 28482
rect 1680 28448 1686 28482
rect 1640 28410 1686 28448
rect 1640 28400 1646 28410
rect 1482 28338 1528 28376
rect 1364 28304 1370 28330
rect 1324 28289 1370 28304
rect 1482 28304 1488 28338
rect 1522 28304 1528 28338
rect 1618 28391 1646 28400
rect 1680 28400 1686 28410
rect 1680 28391 1708 28400
rect 1618 28339 1637 28391
rect 1689 28339 1708 28391
rect 1618 28338 1708 28339
rect 1618 28330 1646 28338
rect 1482 28289 1528 28304
rect 1640 28304 1646 28330
rect 1680 28330 1708 28338
rect 1680 28304 1686 28330
rect 1640 28289 1686 28304
rect 1748 28250 1828 29330
rect 4148 29302 4293 30330
rect 4687 29302 4698 30416
rect 4148 29270 4698 29302
rect 6708 31896 7138 31920
rect 6708 30782 6724 31896
rect 7118 30782 7138 31896
rect 6708 30670 7138 30782
rect 6708 30616 8188 30670
rect 6708 30564 8002 30616
rect 8054 30564 8112 30616
rect 8164 30564 8188 30616
rect 6708 30530 8188 30564
rect 6708 30416 7138 30530
rect 6708 29302 6724 30416
rect 7118 29302 7138 30416
rect 6708 29280 7138 29302
rect -1822 28242 1828 28250
rect -1822 28208 -1593 28242
rect -1559 28208 -1435 28242
rect -1401 28208 -1277 28242
rect -1243 28208 -1119 28242
rect -1085 28208 -961 28242
rect -927 28208 -803 28242
rect -769 28208 -645 28242
rect -611 28208 -487 28242
rect -453 28208 -329 28242
rect -295 28208 -171 28242
rect -137 28208 -13 28242
rect 21 28208 145 28242
rect 179 28208 303 28242
rect 337 28208 461 28242
rect 495 28208 619 28242
rect 653 28208 777 28242
rect 811 28208 935 28242
rect 969 28208 1093 28242
rect 1127 28208 1251 28242
rect 1285 28208 1409 28242
rect 1443 28208 1567 28242
rect 1601 28208 1828 28242
rect -1822 28200 1828 28208
rect 5418 29180 6328 29210
rect 5418 29120 5438 29180
rect 5638 29120 6098 29180
rect 6298 29120 6328 29180
rect -1632 27840 -1362 28200
rect -882 28146 -602 28150
rect -1024 28142 -430 28146
rect -1024 28109 -864 28142
rect -620 28109 -430 28142
rect -1024 27931 -996 28109
rect -458 27931 -430 28109
rect -1024 27898 -864 27931
rect -620 27898 -430 27931
rect -1024 27894 -430 27898
rect -882 27890 -602 27894
rect -132 27840 138 28200
rect 618 28146 898 28150
rect 446 28142 1040 28146
rect 446 28109 636 28142
rect 880 28109 1040 28142
rect 446 27931 474 28109
rect 1012 27931 1040 28109
rect 446 27898 636 27931
rect 880 27898 1040 27931
rect 446 27894 1040 27898
rect 618 27890 898 27894
rect 1368 27840 1638 28200
rect -1632 27830 1638 27840
rect -1632 27796 -1593 27830
rect -1559 27796 -1435 27830
rect -1401 27796 -1277 27830
rect -1243 27796 -1119 27830
rect -1085 27796 -961 27830
rect -927 27796 -803 27830
rect -769 27796 -645 27830
rect -611 27796 -487 27830
rect -453 27796 -329 27830
rect -295 27796 -171 27830
rect -137 27796 -13 27830
rect 21 27796 145 27830
rect 179 27796 303 27830
rect 337 27796 461 27830
rect 495 27796 619 27830
rect 653 27796 777 27830
rect 811 27796 935 27830
rect 969 27796 1093 27830
rect 1127 27796 1251 27830
rect 1285 27796 1409 27830
rect 1443 27796 1567 27830
rect 1601 27796 1638 27830
rect -1632 27790 1638 27796
rect -1678 27734 -1632 27749
rect -1678 27700 -1672 27734
rect -1638 27700 -1632 27734
rect -1520 27734 -1474 27749
rect -1520 27700 -1514 27734
rect -1480 27700 -1474 27734
rect -1362 27734 -1316 27749
rect -1362 27700 -1356 27734
rect -1322 27700 -1316 27734
rect -1212 27734 -1152 27790
rect -1212 27700 -1198 27734
rect -1164 27700 -1152 27734
rect -1046 27734 -1000 27749
rect -1046 27700 -1040 27734
rect -1006 27700 -1000 27734
rect -892 27734 -832 27790
rect -892 27700 -882 27734
rect -848 27700 -832 27734
rect -730 27734 -684 27749
rect -730 27700 -724 27734
rect -690 27700 -684 27734
rect -572 27734 -526 27749
rect -572 27700 -566 27734
rect -532 27700 -526 27734
rect -414 27734 -368 27749
rect -414 27700 -408 27734
rect -374 27700 -368 27734
rect -256 27734 -210 27749
rect -256 27700 -250 27734
rect -216 27700 -210 27734
rect -98 27734 -52 27749
rect -98 27700 -92 27734
rect -58 27700 -52 27734
rect 60 27734 106 27749
rect 60 27700 66 27734
rect 100 27700 106 27734
rect 218 27734 264 27749
rect 218 27700 224 27734
rect 258 27700 264 27734
rect 376 27734 422 27749
rect 376 27700 382 27734
rect 416 27700 422 27734
rect 534 27734 580 27749
rect 534 27700 540 27734
rect 574 27700 580 27734
rect 692 27734 738 27749
rect 692 27700 698 27734
rect 732 27700 738 27734
rect 850 27734 896 27749
rect 850 27700 856 27734
rect 890 27700 896 27734
rect 998 27734 1058 27790
rect 998 27700 1014 27734
rect 1048 27700 1058 27734
rect 1166 27734 1212 27749
rect 1166 27700 1172 27734
rect 1206 27700 1212 27734
rect 1318 27734 1378 27790
rect 1318 27700 1330 27734
rect 1364 27700 1378 27734
rect 1482 27734 1528 27749
rect 1482 27700 1488 27734
rect 1522 27700 1528 27734
rect 1640 27734 1686 27749
rect 1640 27700 1646 27734
rect 1680 27700 1686 27734
rect -1702 27691 -1612 27700
rect -1702 27639 -1683 27691
rect -1631 27639 -1612 27691
rect -1702 27630 -1672 27639
rect -1678 27628 -1672 27630
rect -1638 27630 -1612 27639
rect -1520 27662 -1474 27700
rect -1638 27628 -1632 27630
rect -1678 27590 -1632 27628
rect -1678 27556 -1672 27590
rect -1638 27556 -1632 27590
rect -1678 27518 -1632 27556
rect -1678 27490 -1672 27518
rect -1702 27484 -1672 27490
rect -1638 27490 -1632 27518
rect -1520 27628 -1514 27662
rect -1480 27628 -1474 27662
rect -1382 27691 -1292 27700
rect -1382 27639 -1363 27691
rect -1311 27639 -1292 27691
rect -1382 27630 -1356 27639
rect -1520 27590 -1474 27628
rect -1520 27556 -1514 27590
rect -1480 27556 -1474 27590
rect -1520 27518 -1474 27556
rect -1638 27484 -1612 27490
rect -1702 27481 -1612 27484
rect -1702 27429 -1683 27481
rect -1631 27429 -1612 27481
rect -1702 27420 -1672 27429
rect -1678 27412 -1672 27420
rect -1638 27420 -1612 27429
rect -1520 27484 -1514 27518
rect -1480 27484 -1474 27518
rect -1362 27628 -1356 27630
rect -1322 27630 -1292 27639
rect -1212 27662 -1152 27700
rect -1322 27628 -1316 27630
rect -1362 27590 -1316 27628
rect -1362 27556 -1356 27590
rect -1322 27556 -1316 27590
rect -1362 27518 -1316 27556
rect -1362 27490 -1356 27518
rect -1520 27446 -1474 27484
rect -1638 27412 -1632 27420
rect -1678 27374 -1632 27412
rect -1678 27340 -1672 27374
rect -1638 27340 -1632 27374
rect -1678 27302 -1632 27340
rect -1678 27268 -1672 27302
rect -1638 27268 -1632 27302
rect -1678 27230 -1632 27268
rect -1678 27196 -1672 27230
rect -1638 27196 -1632 27230
rect -1678 27158 -1632 27196
rect -1678 27124 -1672 27158
rect -1638 27124 -1632 27158
rect -1678 27086 -1632 27124
rect -1678 27052 -1672 27086
rect -1638 27052 -1632 27086
rect -1520 27412 -1514 27446
rect -1480 27412 -1474 27446
rect -1382 27484 -1356 27490
rect -1322 27490 -1316 27518
rect -1212 27628 -1198 27662
rect -1164 27628 -1152 27662
rect -1072 27691 -982 27700
rect -1072 27639 -1053 27691
rect -1001 27639 -982 27691
rect -1072 27630 -1040 27639
rect -1212 27590 -1152 27628
rect -1212 27556 -1198 27590
rect -1164 27556 -1152 27590
rect -1212 27518 -1152 27556
rect -1322 27484 -1292 27490
rect -1382 27481 -1292 27484
rect -1382 27429 -1363 27481
rect -1311 27429 -1292 27481
rect -1382 27420 -1356 27429
rect -1520 27374 -1474 27412
rect -1520 27340 -1514 27374
rect -1480 27340 -1474 27374
rect -1520 27302 -1474 27340
rect -1520 27268 -1514 27302
rect -1480 27268 -1474 27302
rect -1520 27230 -1474 27268
rect -1520 27196 -1514 27230
rect -1480 27196 -1474 27230
rect -1520 27158 -1474 27196
rect -1520 27124 -1514 27158
rect -1480 27124 -1474 27158
rect -1520 27086 -1474 27124
rect -1520 27070 -1514 27086
rect -1678 27014 -1632 27052
rect -1678 26980 -1672 27014
rect -1638 26980 -1632 27014
rect -1542 27061 -1514 27070
rect -1480 27070 -1474 27086
rect -1362 27412 -1356 27420
rect -1322 27420 -1292 27429
rect -1212 27484 -1198 27518
rect -1164 27484 -1152 27518
rect -1046 27628 -1040 27630
rect -1006 27630 -982 27639
rect -892 27662 -832 27700
rect -1006 27628 -1000 27630
rect -1046 27590 -1000 27628
rect -1046 27556 -1040 27590
rect -1006 27556 -1000 27590
rect -1046 27518 -1000 27556
rect -1046 27490 -1040 27518
rect -1212 27446 -1152 27484
rect -1322 27412 -1316 27420
rect -1362 27374 -1316 27412
rect -1362 27340 -1356 27374
rect -1322 27340 -1316 27374
rect -1362 27302 -1316 27340
rect -1362 27268 -1356 27302
rect -1322 27268 -1316 27302
rect -1362 27230 -1316 27268
rect -1362 27196 -1356 27230
rect -1322 27196 -1316 27230
rect -1362 27158 -1316 27196
rect -1362 27124 -1356 27158
rect -1322 27124 -1316 27158
rect -1362 27086 -1316 27124
rect -1480 27061 -1452 27070
rect -1542 27009 -1523 27061
rect -1471 27009 -1452 27061
rect -1542 27000 -1514 27009
rect -1678 26942 -1632 26980
rect -1678 26908 -1672 26942
rect -1638 26908 -1632 26942
rect -1678 26870 -1632 26908
rect -1678 26836 -1672 26870
rect -1638 26836 -1632 26870
rect -1520 26980 -1514 27000
rect -1480 27000 -1452 27009
rect -1362 27052 -1356 27086
rect -1322 27052 -1316 27086
rect -1212 27412 -1198 27446
rect -1164 27412 -1152 27446
rect -1072 27484 -1040 27490
rect -1006 27490 -1000 27518
rect -892 27628 -882 27662
rect -848 27628 -832 27662
rect -752 27691 -662 27700
rect -752 27639 -733 27691
rect -681 27639 -662 27691
rect -752 27630 -724 27639
rect -892 27590 -832 27628
rect -892 27556 -882 27590
rect -848 27556 -832 27590
rect -892 27518 -832 27556
rect -1006 27484 -982 27490
rect -1072 27481 -982 27484
rect -1072 27429 -1053 27481
rect -1001 27429 -982 27481
rect -1072 27420 -1040 27429
rect -1212 27374 -1152 27412
rect -1212 27340 -1198 27374
rect -1164 27340 -1152 27374
rect -1212 27302 -1152 27340
rect -1212 27268 -1198 27302
rect -1164 27268 -1152 27302
rect -1212 27230 -1152 27268
rect -1212 27196 -1198 27230
rect -1164 27196 -1152 27230
rect -1212 27158 -1152 27196
rect -1212 27124 -1198 27158
rect -1164 27124 -1152 27158
rect -1212 27086 -1152 27124
rect -1212 27070 -1198 27086
rect -1362 27014 -1316 27052
rect -1480 26980 -1474 27000
rect -1520 26942 -1474 26980
rect -1520 26908 -1514 26942
rect -1480 26908 -1474 26942
rect -1520 26870 -1474 26908
rect -1520 26860 -1514 26870
rect -1678 26798 -1632 26836
rect -1678 26764 -1672 26798
rect -1638 26764 -1632 26798
rect -1542 26851 -1514 26860
rect -1480 26860 -1474 26870
rect -1362 26980 -1356 27014
rect -1322 26980 -1316 27014
rect -1222 27061 -1198 27070
rect -1164 27070 -1152 27086
rect -1046 27412 -1040 27420
rect -1006 27420 -982 27429
rect -892 27484 -882 27518
rect -848 27484 -832 27518
rect -730 27628 -724 27630
rect -690 27630 -662 27639
rect -572 27662 -526 27700
rect -690 27628 -684 27630
rect -730 27590 -684 27628
rect -730 27556 -724 27590
rect -690 27556 -684 27590
rect -730 27518 -684 27556
rect -730 27490 -724 27518
rect -892 27446 -832 27484
rect -1006 27412 -1000 27420
rect -1046 27374 -1000 27412
rect -1046 27340 -1040 27374
rect -1006 27340 -1000 27374
rect -1046 27302 -1000 27340
rect -1046 27268 -1040 27302
rect -1006 27268 -1000 27302
rect -1046 27230 -1000 27268
rect -1046 27196 -1040 27230
rect -1006 27196 -1000 27230
rect -1046 27158 -1000 27196
rect -1046 27124 -1040 27158
rect -1006 27124 -1000 27158
rect -1046 27086 -1000 27124
rect -1164 27061 -1132 27070
rect -1222 27009 -1203 27061
rect -1151 27009 -1132 27061
rect -1222 27000 -1198 27009
rect -1362 26942 -1316 26980
rect -1362 26908 -1356 26942
rect -1322 26908 -1316 26942
rect -1362 26870 -1316 26908
rect -1480 26851 -1452 26860
rect -1542 26799 -1523 26851
rect -1471 26799 -1452 26851
rect -1542 26798 -1452 26799
rect -1542 26790 -1514 26798
rect -1678 26749 -1632 26764
rect -1520 26764 -1514 26790
rect -1480 26790 -1452 26798
rect -1362 26836 -1356 26870
rect -1322 26836 -1316 26870
rect -1212 26980 -1198 27000
rect -1164 27000 -1132 27009
rect -1046 27052 -1040 27086
rect -1006 27052 -1000 27086
rect -892 27412 -882 27446
rect -848 27412 -832 27446
rect -752 27484 -724 27490
rect -690 27490 -684 27518
rect -572 27628 -566 27662
rect -532 27628 -526 27662
rect -432 27691 -342 27700
rect -432 27639 -413 27691
rect -361 27639 -342 27691
rect -432 27630 -408 27639
rect -572 27590 -526 27628
rect -572 27556 -566 27590
rect -532 27556 -526 27590
rect -572 27518 -526 27556
rect -690 27484 -662 27490
rect -752 27481 -662 27484
rect -752 27429 -733 27481
rect -681 27429 -662 27481
rect -752 27420 -724 27429
rect -892 27374 -832 27412
rect -892 27340 -882 27374
rect -848 27340 -832 27374
rect -892 27302 -832 27340
rect -892 27268 -882 27302
rect -848 27268 -832 27302
rect -892 27230 -832 27268
rect -892 27196 -882 27230
rect -848 27196 -832 27230
rect -892 27158 -832 27196
rect -892 27124 -882 27158
rect -848 27124 -832 27158
rect -892 27086 -832 27124
rect -892 27070 -882 27086
rect -1046 27014 -1000 27052
rect -1164 26980 -1152 27000
rect -1212 26942 -1152 26980
rect -1212 26908 -1198 26942
rect -1164 26908 -1152 26942
rect -1212 26870 -1152 26908
rect -1212 26860 -1198 26870
rect -1362 26798 -1316 26836
rect -1480 26764 -1474 26790
rect -1520 26749 -1474 26764
rect -1362 26764 -1356 26798
rect -1322 26764 -1316 26798
rect -1222 26851 -1198 26860
rect -1164 26860 -1152 26870
rect -1046 26980 -1040 27014
rect -1006 26980 -1000 27014
rect -912 27061 -882 27070
rect -848 27070 -832 27086
rect -730 27412 -724 27420
rect -690 27420 -662 27429
rect -572 27484 -566 27518
rect -532 27484 -526 27518
rect -414 27628 -408 27630
rect -374 27630 -342 27639
rect -256 27662 -210 27700
rect -374 27628 -368 27630
rect -414 27590 -368 27628
rect -414 27556 -408 27590
rect -374 27556 -368 27590
rect -414 27518 -368 27556
rect -414 27490 -408 27518
rect -572 27446 -526 27484
rect -690 27412 -684 27420
rect -730 27374 -684 27412
rect -730 27340 -724 27374
rect -690 27340 -684 27374
rect -730 27302 -684 27340
rect -730 27268 -724 27302
rect -690 27268 -684 27302
rect -730 27230 -684 27268
rect -730 27196 -724 27230
rect -690 27196 -684 27230
rect -730 27158 -684 27196
rect -730 27124 -724 27158
rect -690 27124 -684 27158
rect -730 27086 -684 27124
rect -848 27061 -822 27070
rect -912 27009 -893 27061
rect -841 27009 -822 27061
rect -912 27000 -882 27009
rect -1046 26942 -1000 26980
rect -1046 26908 -1040 26942
rect -1006 26908 -1000 26942
rect -1046 26870 -1000 26908
rect -1164 26851 -1132 26860
rect -1222 26799 -1203 26851
rect -1151 26799 -1132 26851
rect -1222 26798 -1132 26799
rect -1222 26790 -1198 26798
rect -1362 26749 -1316 26764
rect -1212 26764 -1198 26790
rect -1164 26790 -1132 26798
rect -1046 26836 -1040 26870
rect -1006 26836 -1000 26870
rect -892 26980 -882 27000
rect -848 27000 -822 27009
rect -730 27052 -724 27086
rect -690 27052 -684 27086
rect -572 27412 -566 27446
rect -532 27412 -526 27446
rect -432 27484 -408 27490
rect -374 27490 -368 27518
rect -256 27628 -250 27662
rect -216 27628 -210 27662
rect -122 27691 -32 27700
rect -122 27639 -103 27691
rect -51 27639 -32 27691
rect -122 27630 -92 27639
rect -256 27590 -210 27628
rect -256 27556 -250 27590
rect -216 27556 -210 27590
rect -256 27518 -210 27556
rect -374 27484 -342 27490
rect -432 27481 -342 27484
rect -432 27429 -413 27481
rect -361 27429 -342 27481
rect -432 27420 -408 27429
rect -572 27374 -526 27412
rect -572 27340 -566 27374
rect -532 27340 -526 27374
rect -572 27302 -526 27340
rect -572 27268 -566 27302
rect -532 27268 -526 27302
rect -572 27230 -526 27268
rect -572 27196 -566 27230
rect -532 27196 -526 27230
rect -572 27158 -526 27196
rect -572 27124 -566 27158
rect -532 27124 -526 27158
rect -572 27086 -526 27124
rect -572 27070 -566 27086
rect -730 27014 -684 27052
rect -848 26980 -832 27000
rect -892 26942 -832 26980
rect -892 26908 -882 26942
rect -848 26908 -832 26942
rect -892 26870 -832 26908
rect -892 26860 -882 26870
rect -1046 26798 -1000 26836
rect -1164 26764 -1152 26790
rect -1212 26710 -1152 26764
rect -1046 26764 -1040 26798
rect -1006 26764 -1000 26798
rect -912 26851 -882 26860
rect -848 26860 -832 26870
rect -730 26980 -724 27014
rect -690 26980 -684 27014
rect -592 27061 -566 27070
rect -532 27070 -526 27086
rect -414 27412 -408 27420
rect -374 27420 -342 27429
rect -256 27484 -250 27518
rect -216 27484 -210 27518
rect -98 27628 -92 27630
rect -58 27630 -32 27639
rect 60 27662 106 27700
rect -58 27628 -52 27630
rect -98 27590 -52 27628
rect -98 27556 -92 27590
rect -58 27556 -52 27590
rect -98 27518 -52 27556
rect -98 27490 -92 27518
rect -256 27446 -210 27484
rect -374 27412 -368 27420
rect -414 27374 -368 27412
rect -414 27340 -408 27374
rect -374 27340 -368 27374
rect -414 27302 -368 27340
rect -414 27268 -408 27302
rect -374 27268 -368 27302
rect -414 27230 -368 27268
rect -414 27196 -408 27230
rect -374 27196 -368 27230
rect -414 27158 -368 27196
rect -414 27124 -408 27158
rect -374 27124 -368 27158
rect -414 27086 -368 27124
rect -532 27061 -502 27070
rect -592 27009 -573 27061
rect -521 27009 -502 27061
rect -592 27000 -566 27009
rect -730 26942 -684 26980
rect -730 26908 -724 26942
rect -690 26908 -684 26942
rect -730 26870 -684 26908
rect -848 26851 -822 26860
rect -912 26799 -893 26851
rect -841 26799 -822 26851
rect -912 26798 -822 26799
rect -912 26790 -882 26798
rect -1046 26749 -1000 26764
rect -892 26764 -882 26790
rect -848 26790 -822 26798
rect -730 26836 -724 26870
rect -690 26836 -684 26870
rect -572 26980 -566 27000
rect -532 27000 -502 27009
rect -414 27052 -408 27086
rect -374 27052 -368 27086
rect -256 27412 -250 27446
rect -216 27412 -210 27446
rect -122 27484 -92 27490
rect -58 27490 -52 27518
rect 60 27628 66 27662
rect 100 27628 106 27662
rect 198 27691 288 27700
rect 198 27639 217 27691
rect 269 27639 288 27691
rect 198 27630 224 27639
rect 60 27590 106 27628
rect 60 27556 66 27590
rect 100 27556 106 27590
rect 60 27518 106 27556
rect -58 27484 -32 27490
rect -122 27481 -32 27484
rect -122 27429 -103 27481
rect -51 27429 -32 27481
rect -122 27420 -92 27429
rect -256 27374 -210 27412
rect -256 27340 -250 27374
rect -216 27340 -210 27374
rect -256 27302 -210 27340
rect -256 27268 -250 27302
rect -216 27268 -210 27302
rect -256 27230 -210 27268
rect -256 27196 -250 27230
rect -216 27196 -210 27230
rect -256 27158 -210 27196
rect -256 27124 -250 27158
rect -216 27124 -210 27158
rect -256 27086 -210 27124
rect -256 27070 -250 27086
rect -414 27014 -368 27052
rect -532 26980 -526 27000
rect -572 26942 -526 26980
rect -572 26908 -566 26942
rect -532 26908 -526 26942
rect -572 26870 -526 26908
rect -572 26860 -566 26870
rect -730 26798 -684 26836
rect -848 26764 -832 26790
rect -892 26710 -832 26764
rect -730 26764 -724 26798
rect -690 26764 -684 26798
rect -592 26851 -566 26860
rect -532 26860 -526 26870
rect -414 26980 -408 27014
rect -374 26980 -368 27014
rect -282 27061 -250 27070
rect -216 27070 -210 27086
rect -98 27412 -92 27420
rect -58 27420 -32 27429
rect 60 27484 66 27518
rect 100 27484 106 27518
rect 218 27628 224 27630
rect 258 27630 288 27639
rect 376 27662 422 27700
rect 258 27628 264 27630
rect 218 27590 264 27628
rect 218 27556 224 27590
rect 258 27556 264 27590
rect 218 27518 264 27556
rect 218 27490 224 27518
rect 60 27446 106 27484
rect -58 27412 -52 27420
rect -98 27374 -52 27412
rect -98 27340 -92 27374
rect -58 27340 -52 27374
rect -98 27302 -52 27340
rect -98 27268 -92 27302
rect -58 27268 -52 27302
rect -98 27230 -52 27268
rect -98 27196 -92 27230
rect -58 27196 -52 27230
rect -98 27158 -52 27196
rect -98 27124 -92 27158
rect -58 27124 -52 27158
rect -98 27086 -52 27124
rect -216 27061 -192 27070
rect -282 27009 -263 27061
rect -211 27009 -192 27061
rect -282 27000 -250 27009
rect -414 26942 -368 26980
rect -414 26908 -408 26942
rect -374 26908 -368 26942
rect -414 26870 -368 26908
rect -532 26851 -502 26860
rect -592 26799 -573 26851
rect -521 26799 -502 26851
rect -592 26798 -502 26799
rect -592 26790 -566 26798
rect -730 26749 -684 26764
rect -572 26764 -566 26790
rect -532 26790 -502 26798
rect -414 26836 -408 26870
rect -374 26836 -368 26870
rect -256 26980 -250 27000
rect -216 27000 -192 27009
rect -98 27052 -92 27086
rect -58 27052 -52 27086
rect 60 27412 66 27446
rect 100 27412 106 27446
rect 198 27484 224 27490
rect 258 27490 264 27518
rect 376 27628 382 27662
rect 416 27628 422 27662
rect 508 27691 598 27700
rect 508 27639 527 27691
rect 579 27639 598 27691
rect 508 27630 540 27639
rect 376 27590 422 27628
rect 376 27556 382 27590
rect 416 27556 422 27590
rect 376 27518 422 27556
rect 258 27484 288 27490
rect 198 27481 288 27484
rect 198 27429 217 27481
rect 269 27429 288 27481
rect 198 27420 224 27429
rect 60 27374 106 27412
rect 60 27340 66 27374
rect 100 27340 106 27374
rect 60 27302 106 27340
rect 60 27268 66 27302
rect 100 27268 106 27302
rect 60 27230 106 27268
rect 60 27196 66 27230
rect 100 27196 106 27230
rect 60 27158 106 27196
rect 60 27124 66 27158
rect 100 27124 106 27158
rect 60 27086 106 27124
rect 60 27070 66 27086
rect -98 27014 -52 27052
rect -216 26980 -210 27000
rect -256 26942 -210 26980
rect -256 26908 -250 26942
rect -216 26908 -210 26942
rect -256 26870 -210 26908
rect -256 26860 -250 26870
rect -414 26798 -368 26836
rect -532 26764 -526 26790
rect -572 26749 -526 26764
rect -414 26764 -408 26798
rect -374 26764 -368 26798
rect -282 26851 -250 26860
rect -216 26860 -210 26870
rect -98 26980 -92 27014
rect -58 26980 -52 27014
rect 38 27061 66 27070
rect 100 27070 106 27086
rect 218 27412 224 27420
rect 258 27420 288 27429
rect 376 27484 382 27518
rect 416 27484 422 27518
rect 534 27628 540 27630
rect 574 27630 598 27639
rect 692 27662 738 27700
rect 574 27628 580 27630
rect 534 27590 580 27628
rect 534 27556 540 27590
rect 574 27556 580 27590
rect 534 27518 580 27556
rect 534 27490 540 27518
rect 376 27446 422 27484
rect 258 27412 264 27420
rect 218 27374 264 27412
rect 218 27340 224 27374
rect 258 27340 264 27374
rect 218 27302 264 27340
rect 218 27268 224 27302
rect 258 27268 264 27302
rect 218 27230 264 27268
rect 218 27196 224 27230
rect 258 27196 264 27230
rect 218 27158 264 27196
rect 218 27124 224 27158
rect 258 27124 264 27158
rect 218 27086 264 27124
rect 100 27061 128 27070
rect 38 27009 57 27061
rect 109 27009 128 27061
rect 38 27000 66 27009
rect -98 26942 -52 26980
rect -98 26908 -92 26942
rect -58 26908 -52 26942
rect -98 26870 -52 26908
rect -216 26851 -192 26860
rect -282 26799 -263 26851
rect -211 26799 -192 26851
rect -282 26798 -192 26799
rect -282 26790 -250 26798
rect -414 26749 -368 26764
rect -256 26764 -250 26790
rect -216 26790 -192 26798
rect -98 26836 -92 26870
rect -58 26836 -52 26870
rect 60 26980 66 27000
rect 100 27000 128 27009
rect 218 27052 224 27086
rect 258 27052 264 27086
rect 376 27412 382 27446
rect 416 27412 422 27446
rect 508 27484 540 27490
rect 574 27490 580 27518
rect 692 27628 698 27662
rect 732 27628 738 27662
rect 828 27691 918 27700
rect 828 27639 847 27691
rect 899 27639 918 27691
rect 828 27630 856 27639
rect 692 27590 738 27628
rect 692 27556 698 27590
rect 732 27556 738 27590
rect 692 27518 738 27556
rect 574 27484 598 27490
rect 508 27481 598 27484
rect 508 27429 527 27481
rect 579 27429 598 27481
rect 508 27420 540 27429
rect 376 27374 422 27412
rect 376 27340 382 27374
rect 416 27340 422 27374
rect 376 27302 422 27340
rect 376 27268 382 27302
rect 416 27268 422 27302
rect 376 27230 422 27268
rect 376 27196 382 27230
rect 416 27196 422 27230
rect 376 27158 422 27196
rect 376 27124 382 27158
rect 416 27124 422 27158
rect 376 27086 422 27124
rect 376 27070 382 27086
rect 218 27014 264 27052
rect 100 26980 106 27000
rect 60 26942 106 26980
rect 60 26908 66 26942
rect 100 26908 106 26942
rect 60 26870 106 26908
rect 60 26860 66 26870
rect -98 26798 -52 26836
rect -216 26764 -210 26790
rect -256 26749 -210 26764
rect -98 26764 -92 26798
rect -58 26764 -52 26798
rect 38 26851 66 26860
rect 100 26860 106 26870
rect 218 26980 224 27014
rect 258 26980 264 27014
rect 358 27061 382 27070
rect 416 27070 422 27086
rect 534 27412 540 27420
rect 574 27420 598 27429
rect 692 27484 698 27518
rect 732 27484 738 27518
rect 850 27628 856 27630
rect 890 27630 918 27639
rect 998 27662 1058 27700
rect 890 27628 896 27630
rect 850 27590 896 27628
rect 850 27556 856 27590
rect 890 27556 896 27590
rect 850 27518 896 27556
rect 850 27490 856 27518
rect 692 27446 738 27484
rect 574 27412 580 27420
rect 534 27374 580 27412
rect 534 27340 540 27374
rect 574 27340 580 27374
rect 534 27302 580 27340
rect 534 27268 540 27302
rect 574 27268 580 27302
rect 534 27230 580 27268
rect 534 27196 540 27230
rect 574 27196 580 27230
rect 534 27158 580 27196
rect 534 27124 540 27158
rect 574 27124 580 27158
rect 534 27086 580 27124
rect 416 27061 448 27070
rect 358 27009 377 27061
rect 429 27009 448 27061
rect 358 27000 382 27009
rect 218 26942 264 26980
rect 218 26908 224 26942
rect 258 26908 264 26942
rect 218 26870 264 26908
rect 100 26851 128 26860
rect 38 26799 57 26851
rect 109 26799 128 26851
rect 38 26798 128 26799
rect 38 26790 66 26798
rect -98 26749 -52 26764
rect 60 26764 66 26790
rect 100 26790 128 26798
rect 218 26836 224 26870
rect 258 26836 264 26870
rect 376 26980 382 27000
rect 416 27000 448 27009
rect 534 27052 540 27086
rect 574 27052 580 27086
rect 692 27412 698 27446
rect 732 27412 738 27446
rect 828 27484 856 27490
rect 890 27490 896 27518
rect 998 27628 1014 27662
rect 1048 27628 1058 27662
rect 1148 27691 1238 27700
rect 1148 27639 1167 27691
rect 1219 27639 1238 27691
rect 1148 27630 1172 27639
rect 998 27590 1058 27628
rect 998 27556 1014 27590
rect 1048 27556 1058 27590
rect 998 27518 1058 27556
rect 890 27484 918 27490
rect 828 27481 918 27484
rect 828 27429 847 27481
rect 899 27429 918 27481
rect 828 27420 856 27429
rect 692 27374 738 27412
rect 692 27340 698 27374
rect 732 27340 738 27374
rect 692 27302 738 27340
rect 692 27268 698 27302
rect 732 27268 738 27302
rect 692 27230 738 27268
rect 692 27196 698 27230
rect 732 27196 738 27230
rect 692 27158 738 27196
rect 692 27124 698 27158
rect 732 27124 738 27158
rect 692 27086 738 27124
rect 692 27070 698 27086
rect 534 27014 580 27052
rect 416 26980 422 27000
rect 376 26942 422 26980
rect 376 26908 382 26942
rect 416 26908 422 26942
rect 376 26870 422 26908
rect 376 26860 382 26870
rect 218 26798 264 26836
rect 100 26764 106 26790
rect 60 26749 106 26764
rect 218 26764 224 26798
rect 258 26764 264 26798
rect 358 26851 382 26860
rect 416 26860 422 26870
rect 534 26980 540 27014
rect 574 26980 580 27014
rect 668 27061 698 27070
rect 732 27070 738 27086
rect 850 27412 856 27420
rect 890 27420 918 27429
rect 998 27484 1014 27518
rect 1048 27484 1058 27518
rect 1166 27628 1172 27630
rect 1206 27630 1238 27639
rect 1318 27662 1378 27700
rect 1206 27628 1212 27630
rect 1166 27590 1212 27628
rect 1166 27556 1172 27590
rect 1206 27556 1212 27590
rect 1166 27518 1212 27556
rect 1166 27490 1172 27518
rect 998 27446 1058 27484
rect 890 27412 896 27420
rect 850 27374 896 27412
rect 850 27340 856 27374
rect 890 27340 896 27374
rect 850 27302 896 27340
rect 850 27268 856 27302
rect 890 27268 896 27302
rect 850 27230 896 27268
rect 850 27196 856 27230
rect 890 27196 896 27230
rect 850 27158 896 27196
rect 850 27124 856 27158
rect 890 27124 896 27158
rect 850 27086 896 27124
rect 732 27061 758 27070
rect 668 27009 687 27061
rect 739 27009 758 27061
rect 668 27000 698 27009
rect 534 26942 580 26980
rect 534 26908 540 26942
rect 574 26908 580 26942
rect 534 26870 580 26908
rect 416 26851 448 26860
rect 358 26799 377 26851
rect 429 26799 448 26851
rect 358 26798 448 26799
rect 358 26790 382 26798
rect 218 26749 264 26764
rect 376 26764 382 26790
rect 416 26790 448 26798
rect 534 26836 540 26870
rect 574 26836 580 26870
rect 692 26980 698 27000
rect 732 27000 758 27009
rect 850 27052 856 27086
rect 890 27052 896 27086
rect 998 27412 1014 27446
rect 1048 27412 1058 27446
rect 1148 27484 1172 27490
rect 1206 27490 1212 27518
rect 1318 27628 1330 27662
rect 1364 27628 1378 27662
rect 1458 27691 1548 27700
rect 1458 27639 1477 27691
rect 1529 27639 1548 27691
rect 1458 27630 1488 27639
rect 1318 27590 1378 27628
rect 1318 27556 1330 27590
rect 1364 27556 1378 27590
rect 1318 27518 1378 27556
rect 1206 27484 1238 27490
rect 1148 27481 1238 27484
rect 1148 27429 1167 27481
rect 1219 27429 1238 27481
rect 1148 27420 1172 27429
rect 998 27374 1058 27412
rect 998 27340 1014 27374
rect 1048 27340 1058 27374
rect 998 27302 1058 27340
rect 998 27268 1014 27302
rect 1048 27268 1058 27302
rect 998 27230 1058 27268
rect 998 27196 1014 27230
rect 1048 27196 1058 27230
rect 998 27158 1058 27196
rect 998 27124 1014 27158
rect 1048 27124 1058 27158
rect 998 27086 1058 27124
rect 998 27070 1014 27086
rect 850 27014 896 27052
rect 732 26980 738 27000
rect 692 26942 738 26980
rect 692 26908 698 26942
rect 732 26908 738 26942
rect 692 26870 738 26908
rect 692 26860 698 26870
rect 534 26798 580 26836
rect 416 26764 422 26790
rect 376 26749 422 26764
rect 534 26764 540 26798
rect 574 26764 580 26798
rect 668 26851 698 26860
rect 732 26860 738 26870
rect 850 26980 856 27014
rect 890 26980 896 27014
rect 988 27061 1014 27070
rect 1048 27070 1058 27086
rect 1166 27412 1172 27420
rect 1206 27420 1238 27429
rect 1318 27484 1330 27518
rect 1364 27484 1378 27518
rect 1482 27628 1488 27630
rect 1522 27630 1548 27639
rect 1640 27662 1686 27700
rect 1522 27628 1528 27630
rect 1482 27590 1528 27628
rect 1482 27556 1488 27590
rect 1522 27556 1528 27590
rect 1482 27518 1528 27556
rect 1482 27490 1488 27518
rect 1318 27446 1378 27484
rect 1206 27412 1212 27420
rect 1166 27374 1212 27412
rect 1166 27340 1172 27374
rect 1206 27340 1212 27374
rect 1166 27302 1212 27340
rect 1166 27268 1172 27302
rect 1206 27268 1212 27302
rect 1166 27230 1212 27268
rect 1166 27196 1172 27230
rect 1206 27196 1212 27230
rect 1166 27158 1212 27196
rect 1166 27124 1172 27158
rect 1206 27124 1212 27158
rect 1166 27086 1212 27124
rect 1048 27061 1078 27070
rect 988 27009 1007 27061
rect 1059 27009 1078 27061
rect 988 27000 1014 27009
rect 850 26942 896 26980
rect 850 26908 856 26942
rect 890 26908 896 26942
rect 850 26870 896 26908
rect 732 26851 758 26860
rect 668 26799 687 26851
rect 739 26799 758 26851
rect 668 26798 758 26799
rect 668 26790 698 26798
rect 534 26749 580 26764
rect 692 26764 698 26790
rect 732 26790 758 26798
rect 850 26836 856 26870
rect 890 26836 896 26870
rect 998 26980 1014 27000
rect 1048 27000 1078 27009
rect 1166 27052 1172 27086
rect 1206 27052 1212 27086
rect 1318 27412 1330 27446
rect 1364 27412 1378 27446
rect 1458 27484 1488 27490
rect 1522 27490 1528 27518
rect 1640 27628 1646 27662
rect 1680 27628 1686 27662
rect 1640 27590 1686 27628
rect 1640 27556 1646 27590
rect 1680 27556 1686 27590
rect 1640 27518 1686 27556
rect 1522 27484 1548 27490
rect 1458 27481 1548 27484
rect 1458 27429 1477 27481
rect 1529 27429 1548 27481
rect 1458 27420 1488 27429
rect 1318 27374 1378 27412
rect 1318 27340 1330 27374
rect 1364 27340 1378 27374
rect 1318 27302 1378 27340
rect 1318 27268 1330 27302
rect 1364 27268 1378 27302
rect 1318 27230 1378 27268
rect 1318 27196 1330 27230
rect 1364 27196 1378 27230
rect 1318 27158 1378 27196
rect 1318 27124 1330 27158
rect 1364 27124 1378 27158
rect 1318 27086 1378 27124
rect 1318 27070 1330 27086
rect 1166 27014 1212 27052
rect 1048 26980 1058 27000
rect 998 26942 1058 26980
rect 998 26908 1014 26942
rect 1048 26908 1058 26942
rect 998 26870 1058 26908
rect 998 26860 1014 26870
rect 850 26798 896 26836
rect 732 26764 738 26790
rect 692 26749 738 26764
rect 850 26764 856 26798
rect 890 26764 896 26798
rect 988 26851 1014 26860
rect 1048 26860 1058 26870
rect 1166 26980 1172 27014
rect 1206 26980 1212 27014
rect 1298 27061 1330 27070
rect 1364 27070 1378 27086
rect 1482 27412 1488 27420
rect 1522 27420 1548 27429
rect 1640 27484 1646 27518
rect 1680 27484 1686 27518
rect 1640 27446 1686 27484
rect 1522 27412 1528 27420
rect 1482 27374 1528 27412
rect 1482 27340 1488 27374
rect 1522 27340 1528 27374
rect 1482 27302 1528 27340
rect 1482 27268 1488 27302
rect 1522 27268 1528 27302
rect 1482 27230 1528 27268
rect 1482 27196 1488 27230
rect 1522 27196 1528 27230
rect 1482 27158 1528 27196
rect 1482 27124 1488 27158
rect 1522 27124 1528 27158
rect 1482 27086 1528 27124
rect 1364 27061 1388 27070
rect 1298 27009 1317 27061
rect 1369 27009 1388 27061
rect 1298 27000 1330 27009
rect 1166 26942 1212 26980
rect 1166 26908 1172 26942
rect 1206 26908 1212 26942
rect 1166 26870 1212 26908
rect 1048 26851 1078 26860
rect 988 26799 1007 26851
rect 1059 26799 1078 26851
rect 988 26798 1078 26799
rect 988 26790 1014 26798
rect 850 26749 896 26764
rect 998 26764 1014 26790
rect 1048 26790 1078 26798
rect 1166 26836 1172 26870
rect 1206 26836 1212 26870
rect 1318 26980 1330 27000
rect 1364 27000 1388 27009
rect 1482 27052 1488 27086
rect 1522 27052 1528 27086
rect 1640 27412 1646 27446
rect 1680 27412 1686 27446
rect 1640 27374 1686 27412
rect 1640 27340 1646 27374
rect 1680 27340 1686 27374
rect 1640 27302 1686 27340
rect 1640 27268 1646 27302
rect 1680 27268 1686 27302
rect 1640 27230 1686 27268
rect 1640 27196 1646 27230
rect 1680 27196 1686 27230
rect 1640 27158 1686 27196
rect 1640 27124 1646 27158
rect 1680 27124 1686 27158
rect 1640 27086 1686 27124
rect 1640 27070 1646 27086
rect 1482 27014 1528 27052
rect 1364 26980 1378 27000
rect 1318 26942 1378 26980
rect 1318 26908 1330 26942
rect 1364 26908 1378 26942
rect 1318 26870 1378 26908
rect 1318 26860 1330 26870
rect 1166 26798 1212 26836
rect 1048 26764 1058 26790
rect 998 26710 1058 26764
rect 1166 26764 1172 26798
rect 1206 26764 1212 26798
rect 1298 26851 1330 26860
rect 1364 26860 1378 26870
rect 1482 26980 1488 27014
rect 1522 26980 1528 27014
rect 1618 27061 1646 27070
rect 1680 27070 1686 27086
rect 1680 27061 1708 27070
rect 1618 27009 1637 27061
rect 1689 27009 1708 27061
rect 1618 27000 1646 27009
rect 1482 26942 1528 26980
rect 1482 26908 1488 26942
rect 1522 26908 1528 26942
rect 1482 26870 1528 26908
rect 1364 26851 1388 26860
rect 1298 26799 1317 26851
rect 1369 26799 1388 26851
rect 1298 26798 1388 26799
rect 1298 26790 1330 26798
rect 1166 26749 1212 26764
rect 1318 26764 1330 26790
rect 1364 26790 1388 26798
rect 1482 26836 1488 26870
rect 1522 26836 1528 26870
rect 1640 26980 1646 27000
rect 1680 27000 1708 27009
rect 1680 26980 1686 27000
rect 1640 26942 1686 26980
rect 1640 26908 1646 26942
rect 1680 26908 1686 26942
rect 1640 26870 1686 26908
rect 1640 26860 1646 26870
rect 1482 26798 1528 26836
rect 1364 26764 1378 26790
rect 1318 26710 1378 26764
rect 1482 26764 1488 26798
rect 1522 26764 1528 26798
rect 1618 26851 1646 26860
rect 1680 26860 1686 26870
rect 1680 26851 1708 26860
rect 1618 26799 1637 26851
rect 1689 26799 1708 26851
rect 1618 26798 1708 26799
rect 1618 26790 1646 26798
rect 1482 26749 1528 26764
rect 1640 26764 1646 26790
rect 1680 26790 1708 26798
rect 1680 26764 1686 26790
rect 1640 26749 1686 26764
rect -1632 26702 1638 26710
rect -1632 26668 -1593 26702
rect -1559 26668 -1435 26702
rect -1401 26668 -1277 26702
rect -1243 26668 -1119 26702
rect -1085 26668 -961 26702
rect -927 26668 -803 26702
rect -769 26668 -645 26702
rect -611 26668 -487 26702
rect -453 26668 -329 26702
rect -295 26668 -171 26702
rect -137 26668 -13 26702
rect 21 26668 145 26702
rect 179 26668 303 26702
rect 337 26668 461 26702
rect 495 26668 619 26702
rect 653 26668 777 26702
rect 811 26668 935 26702
rect 969 26668 1093 26702
rect 1127 26668 1251 26702
rect 1285 26668 1409 26702
rect 1443 26668 1567 26702
rect 1601 26668 1638 26702
rect -1632 26660 1638 26668
rect -338 26355 336 26361
rect -338 26321 -306 26355
rect -272 26321 -234 26355
rect -200 26321 -162 26355
rect -128 26321 -90 26355
rect -56 26321 -18 26355
rect 16 26321 54 26355
rect 88 26321 126 26355
rect 160 26321 198 26355
rect 232 26321 270 26355
rect 304 26321 336 26355
rect -338 26315 336 26321
rect -782 26253 778 26260
rect -782 26219 -492 26253
rect -458 26219 -334 26253
rect -300 26219 -176 26253
rect -142 26219 -18 26253
rect 16 26219 140 26253
rect 174 26219 298 26253
rect 332 26219 456 26253
rect 490 26219 778 26253
rect -782 26210 778 26219
rect -782 25150 -702 26210
rect -577 26166 -531 26181
rect -577 26140 -571 26166
rect -602 26132 -571 26140
rect -537 26140 -531 26166
rect -419 26166 -373 26181
rect -537 26132 -512 26140
rect -602 26131 -512 26132
rect -602 26079 -583 26131
rect -531 26079 -512 26131
rect -602 26070 -571 26079
rect -577 26060 -571 26070
rect -537 26070 -512 26079
rect -419 26132 -413 26166
rect -379 26132 -373 26166
rect -261 26166 -215 26181
rect -261 26140 -255 26166
rect -419 26094 -373 26132
rect -537 26060 -531 26070
rect -577 26022 -531 26060
rect -577 25988 -571 26022
rect -537 25988 -531 26022
rect -577 25950 -531 25988
rect -577 25916 -571 25950
rect -537 25916 -531 25950
rect -577 25878 -531 25916
rect -577 25850 -571 25878
rect -602 25844 -571 25850
rect -537 25850 -531 25878
rect -419 26060 -413 26094
rect -379 26060 -373 26094
rect -282 26132 -255 26140
rect -221 26140 -215 26166
rect -103 26166 -57 26181
rect -221 26132 -192 26140
rect -282 26131 -192 26132
rect -282 26079 -263 26131
rect -211 26079 -192 26131
rect -282 26070 -255 26079
rect -419 26022 -373 26060
rect -419 25988 -413 26022
rect -379 25988 -373 26022
rect -419 25950 -373 25988
rect -419 25916 -413 25950
rect -379 25916 -373 25950
rect -419 25878 -373 25916
rect -537 25844 -512 25850
rect -602 25841 -512 25844
rect -602 25789 -583 25841
rect -531 25789 -512 25841
rect -602 25780 -571 25789
rect -577 25772 -571 25780
rect -537 25780 -512 25789
rect -419 25844 -413 25878
rect -379 25844 -373 25878
rect -261 26060 -255 26070
rect -221 26070 -192 26079
rect -103 26132 -97 26166
rect -63 26132 -57 26166
rect 55 26166 101 26181
rect 55 26140 61 26166
rect -103 26094 -57 26132
rect -221 26060 -215 26070
rect -261 26022 -215 26060
rect -261 25988 -255 26022
rect -221 25988 -215 26022
rect -261 25950 -215 25988
rect -261 25916 -255 25950
rect -221 25916 -215 25950
rect -261 25878 -215 25916
rect -261 25850 -255 25878
rect -419 25806 -373 25844
rect -537 25772 -531 25780
rect -577 25734 -531 25772
rect -577 25700 -571 25734
rect -537 25700 -531 25734
rect -577 25662 -531 25700
rect -577 25628 -571 25662
rect -537 25628 -531 25662
rect -577 25590 -531 25628
rect -577 25556 -571 25590
rect -537 25556 -531 25590
rect -419 25772 -413 25806
rect -379 25772 -373 25806
rect -282 25844 -255 25850
rect -221 25850 -215 25878
rect -103 26060 -97 26094
rect -63 26060 -57 26094
rect 28 26132 61 26140
rect 95 26140 101 26166
rect 213 26166 259 26181
rect 95 26132 118 26140
rect 28 26131 118 26132
rect 28 26079 47 26131
rect 99 26079 118 26131
rect 28 26070 61 26079
rect -103 26022 -57 26060
rect -103 25988 -97 26022
rect -63 25988 -57 26022
rect -103 25950 -57 25988
rect -103 25916 -97 25950
rect -63 25916 -57 25950
rect -103 25878 -57 25916
rect -221 25844 -192 25850
rect -282 25841 -192 25844
rect -282 25789 -263 25841
rect -211 25789 -192 25841
rect -282 25780 -255 25789
rect -419 25734 -373 25772
rect -419 25700 -413 25734
rect -379 25700 -373 25734
rect -419 25662 -373 25700
rect -419 25628 -413 25662
rect -379 25628 -373 25662
rect -419 25590 -373 25628
rect -419 25580 -413 25590
rect -577 25518 -531 25556
rect -577 25484 -571 25518
rect -537 25484 -531 25518
rect -442 25571 -413 25580
rect -379 25580 -373 25590
rect -261 25772 -255 25780
rect -221 25780 -192 25789
rect -103 25844 -97 25878
rect -63 25844 -57 25878
rect 55 26060 61 26070
rect 95 26070 118 26079
rect 213 26132 219 26166
rect 253 26132 259 26166
rect 371 26166 417 26181
rect 371 26140 377 26166
rect 213 26094 259 26132
rect 95 26060 101 26070
rect 55 26022 101 26060
rect 55 25988 61 26022
rect 95 25988 101 26022
rect 55 25950 101 25988
rect 55 25916 61 25950
rect 95 25916 101 25950
rect 55 25878 101 25916
rect 55 25850 61 25878
rect -103 25806 -57 25844
rect -221 25772 -215 25780
rect -261 25734 -215 25772
rect -261 25700 -255 25734
rect -221 25700 -215 25734
rect -261 25662 -215 25700
rect -261 25628 -255 25662
rect -221 25628 -215 25662
rect -261 25590 -215 25628
rect -379 25571 -352 25580
rect -442 25519 -423 25571
rect -371 25519 -352 25571
rect -442 25518 -352 25519
rect -442 25510 -413 25518
rect -577 25446 -531 25484
rect -577 25412 -571 25446
rect -537 25412 -531 25446
rect -577 25374 -531 25412
rect -577 25340 -571 25374
rect -537 25340 -531 25374
rect -577 25302 -531 25340
rect -577 25268 -571 25302
rect -537 25268 -531 25302
rect -419 25484 -413 25510
rect -379 25510 -352 25518
rect -261 25556 -255 25590
rect -221 25556 -215 25590
rect -103 25772 -97 25806
rect -63 25772 -57 25806
rect 28 25844 61 25850
rect 95 25850 101 25878
rect 213 26060 219 26094
rect 253 26060 259 26094
rect 348 26132 377 26140
rect 411 26140 417 26166
rect 529 26166 575 26181
rect 411 26132 438 26140
rect 348 26131 438 26132
rect 348 26079 367 26131
rect 419 26079 438 26131
rect 348 26070 377 26079
rect 213 26022 259 26060
rect 213 25988 219 26022
rect 253 25988 259 26022
rect 213 25950 259 25988
rect 213 25916 219 25950
rect 253 25916 259 25950
rect 213 25878 259 25916
rect 95 25844 118 25850
rect 28 25841 118 25844
rect 28 25789 47 25841
rect 99 25789 118 25841
rect 28 25780 61 25789
rect -103 25734 -57 25772
rect -103 25700 -97 25734
rect -63 25700 -57 25734
rect -103 25662 -57 25700
rect -103 25628 -97 25662
rect -63 25628 -57 25662
rect -103 25590 -57 25628
rect -103 25580 -97 25590
rect -261 25518 -215 25556
rect -379 25484 -373 25510
rect -419 25446 -373 25484
rect -419 25412 -413 25446
rect -379 25412 -373 25446
rect -419 25374 -373 25412
rect -419 25340 -413 25374
rect -379 25340 -373 25374
rect -419 25302 -373 25340
rect -419 25290 -413 25302
rect -577 25230 -531 25268
rect -577 25196 -571 25230
rect -537 25196 -531 25230
rect -442 25281 -413 25290
rect -379 25290 -373 25302
rect -261 25484 -255 25518
rect -221 25484 -215 25518
rect -132 25571 -97 25580
rect -63 25580 -57 25590
rect 55 25772 61 25780
rect 95 25780 118 25789
rect 213 25844 219 25878
rect 253 25844 259 25878
rect 371 26060 377 26070
rect 411 26070 438 26079
rect 529 26132 535 26166
rect 569 26132 575 26166
rect 529 26094 575 26132
rect 411 26060 417 26070
rect 371 26022 417 26060
rect 371 25988 377 26022
rect 411 25988 417 26022
rect 371 25950 417 25988
rect 371 25916 377 25950
rect 411 25916 417 25950
rect 371 25878 417 25916
rect 371 25850 377 25878
rect 213 25806 259 25844
rect 95 25772 101 25780
rect 55 25734 101 25772
rect 55 25700 61 25734
rect 95 25700 101 25734
rect 55 25662 101 25700
rect 55 25628 61 25662
rect 95 25628 101 25662
rect 55 25590 101 25628
rect -63 25571 -42 25580
rect -132 25519 -113 25571
rect -61 25519 -42 25571
rect -132 25518 -42 25519
rect -132 25510 -97 25518
rect -261 25446 -215 25484
rect -261 25412 -255 25446
rect -221 25412 -215 25446
rect -261 25374 -215 25412
rect -261 25340 -255 25374
rect -221 25340 -215 25374
rect -261 25302 -215 25340
rect -379 25281 -352 25290
rect -442 25229 -423 25281
rect -371 25229 -352 25281
rect -442 25220 -413 25229
rect -577 25181 -531 25196
rect -419 25196 -413 25220
rect -379 25220 -352 25229
rect -261 25268 -255 25302
rect -221 25268 -215 25302
rect -103 25484 -97 25510
rect -63 25510 -42 25518
rect 55 25556 61 25590
rect 95 25556 101 25590
rect 213 25772 219 25806
rect 253 25772 259 25806
rect 348 25844 377 25850
rect 411 25850 417 25878
rect 529 26060 535 26094
rect 569 26060 575 26094
rect 529 26022 575 26060
rect 529 25988 535 26022
rect 569 25988 575 26022
rect 529 25950 575 25988
rect 529 25916 535 25950
rect 569 25916 575 25950
rect 529 25878 575 25916
rect 411 25844 438 25850
rect 348 25841 438 25844
rect 348 25789 367 25841
rect 419 25789 438 25841
rect 348 25780 377 25789
rect 213 25734 259 25772
rect 213 25700 219 25734
rect 253 25700 259 25734
rect 213 25662 259 25700
rect 213 25628 219 25662
rect 253 25628 259 25662
rect 213 25590 259 25628
rect 213 25580 219 25590
rect 55 25518 101 25556
rect -63 25484 -57 25510
rect -103 25446 -57 25484
rect -103 25412 -97 25446
rect -63 25412 -57 25446
rect -103 25374 -57 25412
rect -103 25340 -97 25374
rect -63 25340 -57 25374
rect -103 25302 -57 25340
rect -103 25290 -97 25302
rect -261 25230 -215 25268
rect -379 25196 -373 25220
rect -419 25181 -373 25196
rect -261 25196 -255 25230
rect -221 25196 -215 25230
rect -132 25281 -97 25290
rect -63 25290 -57 25302
rect 55 25484 61 25518
rect 95 25484 101 25518
rect 188 25571 219 25580
rect 253 25580 259 25590
rect 371 25772 377 25780
rect 411 25780 438 25789
rect 529 25844 535 25878
rect 569 25844 575 25878
rect 529 25806 575 25844
rect 411 25772 417 25780
rect 371 25734 417 25772
rect 371 25700 377 25734
rect 411 25700 417 25734
rect 371 25662 417 25700
rect 371 25628 377 25662
rect 411 25628 417 25662
rect 371 25590 417 25628
rect 253 25571 278 25580
rect 188 25519 207 25571
rect 259 25519 278 25571
rect 188 25518 278 25519
rect 188 25510 219 25518
rect 55 25446 101 25484
rect 55 25412 61 25446
rect 95 25412 101 25446
rect 55 25374 101 25412
rect 55 25340 61 25374
rect 95 25340 101 25374
rect 55 25302 101 25340
rect -63 25281 -42 25290
rect -132 25229 -113 25281
rect -61 25229 -42 25281
rect -132 25220 -97 25229
rect -261 25181 -215 25196
rect -103 25196 -97 25220
rect -63 25220 -42 25229
rect 55 25268 61 25302
rect 95 25268 101 25302
rect 213 25484 219 25510
rect 253 25510 278 25518
rect 371 25556 377 25590
rect 411 25556 417 25590
rect 529 25772 535 25806
rect 569 25772 575 25806
rect 529 25734 575 25772
rect 529 25700 535 25734
rect 569 25700 575 25734
rect 529 25662 575 25700
rect 529 25628 535 25662
rect 569 25628 575 25662
rect 529 25590 575 25628
rect 529 25580 535 25590
rect 371 25518 417 25556
rect 253 25484 259 25510
rect 213 25446 259 25484
rect 213 25412 219 25446
rect 253 25412 259 25446
rect 213 25374 259 25412
rect 213 25340 219 25374
rect 253 25340 259 25374
rect 213 25302 259 25340
rect 213 25290 219 25302
rect 55 25230 101 25268
rect -63 25196 -57 25220
rect -103 25181 -57 25196
rect 55 25196 61 25230
rect 95 25196 101 25230
rect 188 25281 219 25290
rect 253 25290 259 25302
rect 371 25484 377 25518
rect 411 25484 417 25518
rect 508 25571 535 25580
rect 569 25580 575 25590
rect 569 25571 598 25580
rect 508 25519 527 25571
rect 579 25519 598 25571
rect 508 25518 598 25519
rect 508 25510 535 25518
rect 371 25446 417 25484
rect 371 25412 377 25446
rect 411 25412 417 25446
rect 371 25374 417 25412
rect 371 25340 377 25374
rect 411 25340 417 25374
rect 371 25302 417 25340
rect 253 25281 278 25290
rect 188 25229 207 25281
rect 259 25229 278 25281
rect 188 25220 219 25229
rect 55 25181 101 25196
rect 213 25196 219 25220
rect 253 25220 278 25229
rect 371 25268 377 25302
rect 411 25268 417 25302
rect 529 25484 535 25510
rect 569 25510 598 25518
rect 569 25484 575 25510
rect 529 25446 575 25484
rect 529 25412 535 25446
rect 569 25412 575 25446
rect 529 25374 575 25412
rect 529 25340 535 25374
rect 569 25340 575 25374
rect 529 25302 575 25340
rect 529 25290 535 25302
rect 371 25230 417 25268
rect 253 25196 259 25220
rect 213 25181 259 25196
rect 371 25196 377 25230
rect 411 25196 417 25230
rect 508 25281 535 25290
rect 569 25290 575 25302
rect 569 25281 598 25290
rect 508 25229 527 25281
rect 579 25229 598 25281
rect 508 25220 535 25229
rect 371 25181 417 25196
rect 529 25196 535 25220
rect 569 25220 598 25229
rect 569 25196 575 25220
rect 529 25181 575 25196
rect 698 25150 778 26210
rect -782 25143 778 25150
rect -782 25109 -492 25143
rect -458 25109 -334 25143
rect -300 25109 -176 25143
rect -142 25109 -18 25143
rect 16 25109 140 25143
rect 174 25109 298 25143
rect 332 25109 456 25143
rect 490 25109 778 25143
rect -782 25100 778 25109
rect -142 25047 138 25050
rect -338 25042 336 25047
rect -338 25041 -124 25042
rect 120 25041 336 25042
rect -338 25007 -306 25041
rect -272 25007 -234 25041
rect -200 25007 -162 25041
rect -128 25007 -124 25041
rect 120 25007 126 25041
rect 160 25007 198 25041
rect 232 25007 270 25041
rect 304 25007 336 25041
rect -338 25001 -124 25007
rect -142 24841 -124 25001
rect -338 24835 -124 24841
rect 120 25001 336 25007
rect 120 24841 138 25001
rect 120 24835 336 24841
rect -338 24801 -306 24835
rect -272 24801 -234 24835
rect -200 24801 -162 24835
rect -128 24801 -124 24835
rect 120 24801 126 24835
rect 160 24801 198 24835
rect 232 24801 270 24835
rect 304 24801 336 24835
rect -338 24798 -124 24801
rect 120 24798 336 24801
rect -338 24795 336 24798
rect -142 24790 138 24795
rect -782 24733 778 24740
rect -782 24699 -492 24733
rect -458 24699 -334 24733
rect -300 24699 -176 24733
rect -142 24699 -18 24733
rect 16 24699 140 24733
rect 174 24699 298 24733
rect 332 24699 456 24733
rect 490 24699 778 24733
rect -782 24690 778 24699
rect -782 23630 -702 24690
rect -577 24646 -531 24661
rect -577 24620 -571 24646
rect -602 24612 -571 24620
rect -537 24620 -531 24646
rect -419 24646 -373 24661
rect -537 24612 -512 24620
rect -602 24611 -512 24612
rect -602 24559 -583 24611
rect -531 24559 -512 24611
rect -602 24550 -571 24559
rect -577 24540 -571 24550
rect -537 24550 -512 24559
rect -419 24612 -413 24646
rect -379 24612 -373 24646
rect -261 24646 -215 24661
rect -261 24620 -255 24646
rect -419 24574 -373 24612
rect -537 24540 -531 24550
rect -577 24502 -531 24540
rect -577 24468 -571 24502
rect -537 24468 -531 24502
rect -577 24430 -531 24468
rect -577 24396 -571 24430
rect -537 24396 -531 24430
rect -577 24358 -531 24396
rect -577 24330 -571 24358
rect -602 24324 -571 24330
rect -537 24330 -531 24358
rect -419 24540 -413 24574
rect -379 24540 -373 24574
rect -282 24612 -255 24620
rect -221 24620 -215 24646
rect -103 24646 -57 24661
rect -221 24612 -192 24620
rect -282 24611 -192 24612
rect -282 24559 -263 24611
rect -211 24559 -192 24611
rect -282 24550 -255 24559
rect -419 24502 -373 24540
rect -419 24468 -413 24502
rect -379 24468 -373 24502
rect -419 24430 -373 24468
rect -419 24396 -413 24430
rect -379 24396 -373 24430
rect -419 24358 -373 24396
rect -537 24324 -512 24330
rect -602 24321 -512 24324
rect -602 24269 -583 24321
rect -531 24269 -512 24321
rect -602 24260 -571 24269
rect -577 24252 -571 24260
rect -537 24260 -512 24269
rect -419 24324 -413 24358
rect -379 24324 -373 24358
rect -261 24540 -255 24550
rect -221 24550 -192 24559
rect -103 24612 -97 24646
rect -63 24612 -57 24646
rect 55 24646 101 24661
rect 55 24620 61 24646
rect -103 24574 -57 24612
rect -221 24540 -215 24550
rect -261 24502 -215 24540
rect -261 24468 -255 24502
rect -221 24468 -215 24502
rect -261 24430 -215 24468
rect -261 24396 -255 24430
rect -221 24396 -215 24430
rect -261 24358 -215 24396
rect -261 24330 -255 24358
rect -419 24286 -373 24324
rect -537 24252 -531 24260
rect -577 24214 -531 24252
rect -577 24180 -571 24214
rect -537 24180 -531 24214
rect -577 24142 -531 24180
rect -577 24108 -571 24142
rect -537 24108 -531 24142
rect -577 24070 -531 24108
rect -577 24036 -571 24070
rect -537 24036 -531 24070
rect -419 24252 -413 24286
rect -379 24252 -373 24286
rect -282 24324 -255 24330
rect -221 24330 -215 24358
rect -103 24540 -97 24574
rect -63 24540 -57 24574
rect 28 24612 61 24620
rect 95 24620 101 24646
rect 213 24646 259 24661
rect 95 24612 118 24620
rect 28 24611 118 24612
rect 28 24559 47 24611
rect 99 24559 118 24611
rect 28 24550 61 24559
rect -103 24502 -57 24540
rect -103 24468 -97 24502
rect -63 24468 -57 24502
rect -103 24430 -57 24468
rect -103 24396 -97 24430
rect -63 24396 -57 24430
rect -103 24358 -57 24396
rect -221 24324 -192 24330
rect -282 24321 -192 24324
rect -282 24269 -263 24321
rect -211 24269 -192 24321
rect -282 24260 -255 24269
rect -419 24214 -373 24252
rect -419 24180 -413 24214
rect -379 24180 -373 24214
rect -419 24142 -373 24180
rect -419 24108 -413 24142
rect -379 24108 -373 24142
rect -419 24070 -373 24108
rect -419 24060 -413 24070
rect -577 23998 -531 24036
rect -577 23964 -571 23998
rect -537 23964 -531 23998
rect -442 24051 -413 24060
rect -379 24060 -373 24070
rect -261 24252 -255 24260
rect -221 24260 -192 24269
rect -103 24324 -97 24358
rect -63 24324 -57 24358
rect 55 24540 61 24550
rect 95 24550 118 24559
rect 213 24612 219 24646
rect 253 24612 259 24646
rect 371 24646 417 24661
rect 371 24620 377 24646
rect 213 24574 259 24612
rect 95 24540 101 24550
rect 55 24502 101 24540
rect 55 24468 61 24502
rect 95 24468 101 24502
rect 55 24430 101 24468
rect 55 24396 61 24430
rect 95 24396 101 24430
rect 55 24358 101 24396
rect 55 24330 61 24358
rect -103 24286 -57 24324
rect -221 24252 -215 24260
rect -261 24214 -215 24252
rect -261 24180 -255 24214
rect -221 24180 -215 24214
rect -261 24142 -215 24180
rect -261 24108 -255 24142
rect -221 24108 -215 24142
rect -261 24070 -215 24108
rect -379 24051 -352 24060
rect -442 23999 -423 24051
rect -371 23999 -352 24051
rect -442 23998 -352 23999
rect -442 23990 -413 23998
rect -577 23926 -531 23964
rect -577 23892 -571 23926
rect -537 23892 -531 23926
rect -577 23854 -531 23892
rect -577 23820 -571 23854
rect -537 23820 -531 23854
rect -577 23782 -531 23820
rect -577 23748 -571 23782
rect -537 23748 -531 23782
rect -419 23964 -413 23990
rect -379 23990 -352 23998
rect -261 24036 -255 24070
rect -221 24036 -215 24070
rect -103 24252 -97 24286
rect -63 24252 -57 24286
rect 28 24324 61 24330
rect 95 24330 101 24358
rect 213 24540 219 24574
rect 253 24540 259 24574
rect 348 24612 377 24620
rect 411 24620 417 24646
rect 529 24646 575 24661
rect 411 24612 438 24620
rect 348 24611 438 24612
rect 348 24559 367 24611
rect 419 24559 438 24611
rect 348 24550 377 24559
rect 213 24502 259 24540
rect 213 24468 219 24502
rect 253 24468 259 24502
rect 213 24430 259 24468
rect 213 24396 219 24430
rect 253 24396 259 24430
rect 213 24358 259 24396
rect 95 24324 118 24330
rect 28 24321 118 24324
rect 28 24269 47 24321
rect 99 24269 118 24321
rect 28 24260 61 24269
rect -103 24214 -57 24252
rect -103 24180 -97 24214
rect -63 24180 -57 24214
rect -103 24142 -57 24180
rect -103 24108 -97 24142
rect -63 24108 -57 24142
rect -103 24070 -57 24108
rect -103 24060 -97 24070
rect -261 23998 -215 24036
rect -379 23964 -373 23990
rect -419 23926 -373 23964
rect -419 23892 -413 23926
rect -379 23892 -373 23926
rect -419 23854 -373 23892
rect -419 23820 -413 23854
rect -379 23820 -373 23854
rect -419 23782 -373 23820
rect -419 23770 -413 23782
rect -577 23710 -531 23748
rect -577 23676 -571 23710
rect -537 23676 -531 23710
rect -442 23761 -413 23770
rect -379 23770 -373 23782
rect -261 23964 -255 23998
rect -221 23964 -215 23998
rect -132 24051 -97 24060
rect -63 24060 -57 24070
rect 55 24252 61 24260
rect 95 24260 118 24269
rect 213 24324 219 24358
rect 253 24324 259 24358
rect 371 24540 377 24550
rect 411 24550 438 24559
rect 529 24612 535 24646
rect 569 24612 575 24646
rect 529 24574 575 24612
rect 411 24540 417 24550
rect 371 24502 417 24540
rect 371 24468 377 24502
rect 411 24468 417 24502
rect 371 24430 417 24468
rect 371 24396 377 24430
rect 411 24396 417 24430
rect 371 24358 417 24396
rect 371 24330 377 24358
rect 213 24286 259 24324
rect 95 24252 101 24260
rect 55 24214 101 24252
rect 55 24180 61 24214
rect 95 24180 101 24214
rect 55 24142 101 24180
rect 55 24108 61 24142
rect 95 24108 101 24142
rect 55 24070 101 24108
rect -63 24051 -42 24060
rect -132 23999 -113 24051
rect -61 23999 -42 24051
rect -132 23998 -42 23999
rect -132 23990 -97 23998
rect -261 23926 -215 23964
rect -261 23892 -255 23926
rect -221 23892 -215 23926
rect -261 23854 -215 23892
rect -261 23820 -255 23854
rect -221 23820 -215 23854
rect -261 23782 -215 23820
rect -379 23761 -352 23770
rect -442 23709 -423 23761
rect -371 23709 -352 23761
rect -442 23700 -413 23709
rect -577 23661 -531 23676
rect -419 23676 -413 23700
rect -379 23700 -352 23709
rect -261 23748 -255 23782
rect -221 23748 -215 23782
rect -103 23964 -97 23990
rect -63 23990 -42 23998
rect 55 24036 61 24070
rect 95 24036 101 24070
rect 213 24252 219 24286
rect 253 24252 259 24286
rect 348 24324 377 24330
rect 411 24330 417 24358
rect 529 24540 535 24574
rect 569 24540 575 24574
rect 529 24502 575 24540
rect 529 24468 535 24502
rect 569 24468 575 24502
rect 529 24430 575 24468
rect 529 24396 535 24430
rect 569 24396 575 24430
rect 529 24358 575 24396
rect 411 24324 438 24330
rect 348 24321 438 24324
rect 348 24269 367 24321
rect 419 24269 438 24321
rect 348 24260 377 24269
rect 213 24214 259 24252
rect 213 24180 219 24214
rect 253 24180 259 24214
rect 213 24142 259 24180
rect 213 24108 219 24142
rect 253 24108 259 24142
rect 213 24070 259 24108
rect 213 24060 219 24070
rect 55 23998 101 24036
rect -63 23964 -57 23990
rect -103 23926 -57 23964
rect -103 23892 -97 23926
rect -63 23892 -57 23926
rect -103 23854 -57 23892
rect -103 23820 -97 23854
rect -63 23820 -57 23854
rect -103 23782 -57 23820
rect -103 23770 -97 23782
rect -261 23710 -215 23748
rect -379 23676 -373 23700
rect -419 23661 -373 23676
rect -261 23676 -255 23710
rect -221 23676 -215 23710
rect -132 23761 -97 23770
rect -63 23770 -57 23782
rect 55 23964 61 23998
rect 95 23964 101 23998
rect 188 24051 219 24060
rect 253 24060 259 24070
rect 371 24252 377 24260
rect 411 24260 438 24269
rect 529 24324 535 24358
rect 569 24324 575 24358
rect 529 24286 575 24324
rect 411 24252 417 24260
rect 371 24214 417 24252
rect 371 24180 377 24214
rect 411 24180 417 24214
rect 371 24142 417 24180
rect 371 24108 377 24142
rect 411 24108 417 24142
rect 371 24070 417 24108
rect 253 24051 278 24060
rect 188 23999 207 24051
rect 259 23999 278 24051
rect 188 23998 278 23999
rect 188 23990 219 23998
rect 55 23926 101 23964
rect 55 23892 61 23926
rect 95 23892 101 23926
rect 55 23854 101 23892
rect 55 23820 61 23854
rect 95 23820 101 23854
rect 55 23782 101 23820
rect -63 23761 -42 23770
rect -132 23709 -113 23761
rect -61 23709 -42 23761
rect -132 23700 -97 23709
rect -261 23661 -215 23676
rect -103 23676 -97 23700
rect -63 23700 -42 23709
rect 55 23748 61 23782
rect 95 23748 101 23782
rect 213 23964 219 23990
rect 253 23990 278 23998
rect 371 24036 377 24070
rect 411 24036 417 24070
rect 529 24252 535 24286
rect 569 24252 575 24286
rect 529 24214 575 24252
rect 529 24180 535 24214
rect 569 24180 575 24214
rect 529 24142 575 24180
rect 529 24108 535 24142
rect 569 24108 575 24142
rect 529 24070 575 24108
rect 529 24060 535 24070
rect 371 23998 417 24036
rect 253 23964 259 23990
rect 213 23926 259 23964
rect 213 23892 219 23926
rect 253 23892 259 23926
rect 213 23854 259 23892
rect 213 23820 219 23854
rect 253 23820 259 23854
rect 213 23782 259 23820
rect 213 23770 219 23782
rect 55 23710 101 23748
rect -63 23676 -57 23700
rect -103 23661 -57 23676
rect 55 23676 61 23710
rect 95 23676 101 23710
rect 188 23761 219 23770
rect 253 23770 259 23782
rect 371 23964 377 23998
rect 411 23964 417 23998
rect 508 24051 535 24060
rect 569 24060 575 24070
rect 569 24051 598 24060
rect 508 23999 527 24051
rect 579 23999 598 24051
rect 508 23998 598 23999
rect 508 23990 535 23998
rect 371 23926 417 23964
rect 371 23892 377 23926
rect 411 23892 417 23926
rect 371 23854 417 23892
rect 371 23820 377 23854
rect 411 23820 417 23854
rect 371 23782 417 23820
rect 253 23761 278 23770
rect 188 23709 207 23761
rect 259 23709 278 23761
rect 188 23700 219 23709
rect 55 23661 101 23676
rect 213 23676 219 23700
rect 253 23700 278 23709
rect 371 23748 377 23782
rect 411 23748 417 23782
rect 529 23964 535 23990
rect 569 23990 598 23998
rect 569 23964 575 23990
rect 529 23926 575 23964
rect 529 23892 535 23926
rect 569 23892 575 23926
rect 529 23854 575 23892
rect 529 23820 535 23854
rect 569 23820 575 23854
rect 529 23782 575 23820
rect 529 23770 535 23782
rect 371 23710 417 23748
rect 253 23676 259 23700
rect 213 23661 259 23676
rect 371 23676 377 23710
rect 411 23676 417 23710
rect 508 23761 535 23770
rect 569 23770 575 23782
rect 569 23761 598 23770
rect 508 23709 527 23761
rect 579 23709 598 23761
rect 508 23700 535 23709
rect 371 23661 417 23676
rect 529 23676 535 23700
rect 569 23700 598 23709
rect 569 23676 575 23700
rect 529 23661 575 23676
rect 698 23630 778 24690
rect -782 23623 778 23630
rect -782 23589 -492 23623
rect -458 23589 -334 23623
rect -300 23589 -176 23623
rect -142 23589 -18 23623
rect 16 23589 140 23623
rect 174 23589 298 23623
rect 332 23589 456 23623
rect 490 23589 778 23623
rect -782 23580 778 23589
rect -142 23527 138 23530
rect -338 23522 336 23527
rect -338 23521 -124 23522
rect 120 23521 336 23522
rect -338 23487 -306 23521
rect -272 23487 -234 23521
rect -200 23487 -162 23521
rect -128 23487 -124 23521
rect 120 23487 126 23521
rect 160 23487 198 23521
rect 232 23487 270 23521
rect 304 23487 336 23521
rect -338 23481 -124 23487
rect -142 23320 -124 23481
rect -831 23314 -124 23320
rect 120 23481 336 23487
rect 120 23320 138 23481
rect 120 23314 837 23320
rect -831 23280 -806 23314
rect -772 23280 -734 23314
rect -700 23280 -662 23314
rect -628 23280 -590 23314
rect -556 23280 -518 23314
rect -484 23280 -446 23314
rect -412 23280 -374 23314
rect -340 23280 -302 23314
rect -268 23280 -230 23314
rect -196 23280 -158 23314
rect 120 23280 130 23314
rect 164 23280 202 23314
rect 236 23280 274 23314
rect 308 23280 346 23314
rect 380 23280 418 23314
rect 452 23280 490 23314
rect 524 23280 562 23314
rect 596 23280 634 23314
rect 668 23280 706 23314
rect 740 23280 778 23314
rect 812 23280 837 23314
rect -831 23278 -124 23280
rect 120 23278 837 23280
rect -831 23274 837 23278
rect -142 23270 138 23274
rect -2402 23221 -2272 23250
rect -2402 23220 -2363 23221
rect -2412 23170 -2363 23220
rect -2402 23169 -2363 23170
rect -2311 23220 -2272 23221
rect -2152 23221 -2022 23250
rect -2152 23220 -2113 23221
rect -2311 23170 -2113 23220
rect -2311 23169 -2272 23170
rect -2402 23140 -2272 23169
rect -2152 23169 -2113 23170
rect -2061 23220 -2022 23221
rect 1998 23221 2128 23250
rect 1998 23220 2037 23221
rect -2061 23212 2037 23220
rect -2061 23178 -1469 23212
rect -1435 23178 -1397 23212
rect -1363 23178 -1211 23212
rect -1177 23178 -1139 23212
rect -1105 23178 -953 23212
rect -919 23178 -881 23212
rect -847 23178 -695 23212
rect -661 23178 -623 23212
rect -589 23178 -437 23212
rect -403 23178 -365 23212
rect -331 23178 -179 23212
rect -145 23178 -107 23212
rect -73 23178 79 23212
rect 113 23178 151 23212
rect 185 23178 337 23212
rect 371 23178 409 23212
rect 443 23178 595 23212
rect 629 23178 667 23212
rect 701 23178 853 23212
rect 887 23178 925 23212
rect 959 23178 1111 23212
rect 1145 23178 1183 23212
rect 1217 23178 1369 23212
rect 1403 23178 1441 23212
rect 1475 23178 2037 23212
rect -2061 23170 2037 23178
rect -2061 23169 -2022 23170
rect -2152 23140 -2022 23169
rect 1998 23169 2037 23170
rect 2089 23220 2128 23221
rect 2248 23221 2378 23250
rect 2248 23220 2287 23221
rect 2089 23170 2287 23220
rect 2089 23169 2128 23170
rect 1998 23140 2128 23169
rect 2248 23169 2287 23170
rect 2339 23220 2378 23221
rect 2339 23170 2388 23220
rect 2339 23169 2378 23170
rect 2248 23140 2378 23169
rect -1568 23125 -1522 23140
rect -1568 23100 -1562 23125
rect -1592 23091 -1562 23100
rect -1528 23100 -1522 23125
rect -1310 23125 -1264 23140
rect -1528 23091 -1502 23100
rect -1592 23039 -1573 23091
rect -1521 23039 -1502 23091
rect -1592 23030 -1562 23039
rect -1568 23019 -1562 23030
rect -1528 23030 -1502 23039
rect -1310 23091 -1304 23125
rect -1270 23091 -1264 23125
rect -1052 23125 -1006 23140
rect -1052 23100 -1046 23125
rect -1310 23053 -1264 23091
rect -1528 23019 -1522 23030
rect -1568 22981 -1522 23019
rect -1568 22947 -1562 22981
rect -1528 22947 -1522 22981
rect -1568 22920 -1522 22947
rect -1310 23019 -1304 23053
rect -1270 23019 -1264 23053
rect -1072 23091 -1046 23100
rect -1012 23100 -1006 23125
rect -794 23125 -748 23140
rect -1012 23091 -982 23100
rect -1072 23039 -1053 23091
rect -1001 23039 -982 23091
rect -1072 23030 -1046 23039
rect -1310 22981 -1264 23019
rect -1310 22947 -1304 22981
rect -1270 22947 -1264 22981
rect -1592 22911 -1502 22920
rect -1592 22859 -1573 22911
rect -1521 22859 -1502 22911
rect -1592 22850 -1502 22859
rect -1310 22909 -1264 22947
rect -1052 23019 -1046 23030
rect -1012 23030 -982 23039
rect -794 23091 -788 23125
rect -754 23091 -748 23125
rect -536 23125 -490 23140
rect -536 23100 -530 23125
rect -794 23053 -748 23091
rect -1012 23019 -1006 23030
rect -1052 22981 -1006 23019
rect -1052 22947 -1046 22981
rect -1012 22947 -1006 22981
rect -1052 22920 -1006 22947
rect -794 23019 -788 23053
rect -754 23019 -748 23053
rect -562 23091 -530 23100
rect -496 23100 -490 23125
rect -278 23125 -232 23140
rect -496 23091 -472 23100
rect -562 23039 -543 23091
rect -491 23039 -472 23091
rect -562 23030 -530 23039
rect -794 22981 -748 23019
rect -794 22947 -788 22981
rect -754 22947 -748 22981
rect -1310 22875 -1304 22909
rect -1270 22875 -1264 22909
rect -1568 22837 -1522 22850
rect -1568 22803 -1562 22837
rect -1528 22803 -1522 22837
rect -1568 22765 -1522 22803
rect -1568 22731 -1562 22765
rect -1528 22731 -1522 22765
rect -1568 22693 -1522 22731
rect -1568 22659 -1562 22693
rect -1528 22659 -1522 22693
rect -1568 22621 -1522 22659
rect -1568 22587 -1562 22621
rect -1528 22587 -1522 22621
rect -1568 22549 -1522 22587
rect -1568 22515 -1562 22549
rect -1528 22515 -1522 22549
rect -1568 22477 -1522 22515
rect -1568 22443 -1562 22477
rect -1528 22443 -1522 22477
rect -1568 22405 -1522 22443
rect -1310 22837 -1264 22875
rect -1072 22911 -982 22920
rect -1072 22859 -1053 22911
rect -1001 22859 -982 22911
rect -1072 22850 -982 22859
rect -794 22909 -748 22947
rect -536 23019 -530 23030
rect -496 23030 -472 23039
rect -278 23091 -272 23125
rect -238 23091 -232 23125
rect -20 23125 26 23140
rect -20 23100 -14 23125
rect -278 23053 -232 23091
rect -496 23019 -490 23030
rect -536 22981 -490 23019
rect -536 22947 -530 22981
rect -496 22947 -490 22981
rect -536 22920 -490 22947
rect -278 23019 -272 23053
rect -238 23019 -232 23053
rect -42 23091 -14 23100
rect 20 23100 26 23125
rect 238 23125 284 23140
rect 20 23091 48 23100
rect -42 23039 -23 23091
rect 29 23039 48 23091
rect -42 23030 -14 23039
rect -278 22981 -232 23019
rect -278 22947 -272 22981
rect -238 22947 -232 22981
rect -794 22875 -788 22909
rect -754 22875 -748 22909
rect -1310 22803 -1304 22837
rect -1270 22803 -1264 22837
rect -1310 22765 -1264 22803
rect -1310 22731 -1304 22765
rect -1270 22731 -1264 22765
rect -1310 22693 -1264 22731
rect -1310 22659 -1304 22693
rect -1270 22659 -1264 22693
rect -1310 22621 -1264 22659
rect -1310 22587 -1304 22621
rect -1270 22587 -1264 22621
rect -1310 22549 -1264 22587
rect -1310 22515 -1304 22549
rect -1270 22515 -1264 22549
rect -1310 22477 -1264 22515
rect -1310 22443 -1304 22477
rect -1270 22443 -1264 22477
rect -1310 22430 -1264 22443
rect -1052 22837 -1006 22850
rect -1052 22803 -1046 22837
rect -1012 22803 -1006 22837
rect -1052 22765 -1006 22803
rect -1052 22731 -1046 22765
rect -1012 22731 -1006 22765
rect -1052 22693 -1006 22731
rect -1052 22659 -1046 22693
rect -1012 22659 -1006 22693
rect -1052 22621 -1006 22659
rect -1052 22587 -1046 22621
rect -1012 22587 -1006 22621
rect -1052 22549 -1006 22587
rect -1052 22515 -1046 22549
rect -1012 22515 -1006 22549
rect -1052 22477 -1006 22515
rect -1052 22443 -1046 22477
rect -1012 22443 -1006 22477
rect -1568 22371 -1562 22405
rect -1528 22371 -1522 22405
rect -1568 22333 -1522 22371
rect -1332 22421 -1242 22430
rect -1332 22369 -1313 22421
rect -1261 22369 -1242 22421
rect -1332 22360 -1242 22369
rect -1052 22405 -1006 22443
rect -794 22837 -748 22875
rect -562 22911 -472 22920
rect -562 22859 -543 22911
rect -491 22859 -472 22911
rect -562 22850 -472 22859
rect -278 22909 -232 22947
rect -20 23019 -14 23030
rect 20 23030 48 23039
rect 238 23091 244 23125
rect 278 23091 284 23125
rect 496 23125 542 23140
rect 496 23100 502 23125
rect 238 23053 284 23091
rect 20 23019 26 23030
rect -20 22981 26 23019
rect -20 22947 -14 22981
rect 20 22947 26 22981
rect -20 22920 26 22947
rect 238 23019 244 23053
rect 278 23019 284 23053
rect 468 23091 502 23100
rect 536 23100 542 23125
rect 754 23125 800 23140
rect 536 23091 558 23100
rect 468 23039 487 23091
rect 539 23039 558 23091
rect 468 23030 502 23039
rect 238 22981 284 23019
rect 238 22947 244 22981
rect 278 22947 284 22981
rect -278 22875 -272 22909
rect -238 22875 -232 22909
rect -794 22803 -788 22837
rect -754 22803 -748 22837
rect -794 22765 -748 22803
rect -794 22731 -788 22765
rect -754 22731 -748 22765
rect -794 22693 -748 22731
rect -794 22659 -788 22693
rect -754 22659 -748 22693
rect -794 22621 -748 22659
rect -794 22587 -788 22621
rect -754 22587 -748 22621
rect -794 22549 -748 22587
rect -794 22515 -788 22549
rect -754 22515 -748 22549
rect -794 22477 -748 22515
rect -794 22443 -788 22477
rect -754 22443 -748 22477
rect -794 22430 -748 22443
rect -536 22837 -490 22850
rect -536 22803 -530 22837
rect -496 22803 -490 22837
rect -536 22765 -490 22803
rect -536 22731 -530 22765
rect -496 22731 -490 22765
rect -536 22693 -490 22731
rect -536 22659 -530 22693
rect -496 22659 -490 22693
rect -536 22621 -490 22659
rect -536 22587 -530 22621
rect -496 22587 -490 22621
rect -536 22549 -490 22587
rect -536 22515 -530 22549
rect -496 22515 -490 22549
rect -536 22477 -490 22515
rect -536 22443 -530 22477
rect -496 22443 -490 22477
rect -1052 22371 -1046 22405
rect -1012 22371 -1006 22405
rect -1568 22299 -1562 22333
rect -1528 22299 -1522 22333
rect -1568 22261 -1522 22299
rect -1568 22227 -1562 22261
rect -1528 22227 -1522 22261
rect -1310 22333 -1264 22360
rect -1310 22299 -1304 22333
rect -1270 22299 -1264 22333
rect -1310 22261 -1264 22299
rect -1310 22250 -1304 22261
rect -1568 22189 -1522 22227
rect -1568 22155 -1562 22189
rect -1528 22155 -1522 22189
rect -1332 22241 -1304 22250
rect -1270 22250 -1264 22261
rect -1052 22333 -1006 22371
rect -822 22421 -732 22430
rect -822 22369 -803 22421
rect -751 22369 -732 22421
rect -822 22360 -732 22369
rect -536 22405 -490 22443
rect -278 22837 -232 22875
rect -42 22911 48 22920
rect -42 22859 -23 22911
rect 29 22859 48 22911
rect -42 22850 48 22859
rect 238 22909 284 22947
rect 496 23019 502 23030
rect 536 23030 558 23039
rect 754 23091 760 23125
rect 794 23091 800 23125
rect 1012 23125 1058 23140
rect 1012 23100 1018 23125
rect 754 23053 800 23091
rect 536 23019 542 23030
rect 496 22981 542 23019
rect 496 22947 502 22981
rect 536 22947 542 22981
rect 496 22920 542 22947
rect 754 23019 760 23053
rect 794 23019 800 23053
rect 988 23091 1018 23100
rect 1052 23100 1058 23125
rect 1270 23125 1316 23140
rect 1052 23091 1078 23100
rect 988 23039 1007 23091
rect 1059 23039 1078 23091
rect 988 23030 1018 23039
rect 754 22981 800 23019
rect 754 22947 760 22981
rect 794 22947 800 22981
rect 238 22875 244 22909
rect 278 22875 284 22909
rect -278 22803 -272 22837
rect -238 22803 -232 22837
rect -278 22765 -232 22803
rect -278 22731 -272 22765
rect -238 22731 -232 22765
rect -278 22693 -232 22731
rect -278 22659 -272 22693
rect -238 22659 -232 22693
rect -278 22621 -232 22659
rect -278 22587 -272 22621
rect -238 22587 -232 22621
rect -278 22549 -232 22587
rect -278 22515 -272 22549
rect -238 22515 -232 22549
rect -278 22477 -232 22515
rect -278 22443 -272 22477
rect -238 22443 -232 22477
rect -278 22430 -232 22443
rect -20 22837 26 22850
rect -20 22803 -14 22837
rect 20 22803 26 22837
rect -20 22765 26 22803
rect -20 22731 -14 22765
rect 20 22731 26 22765
rect -20 22693 26 22731
rect -20 22659 -14 22693
rect 20 22659 26 22693
rect -20 22621 26 22659
rect -20 22587 -14 22621
rect 20 22587 26 22621
rect -20 22549 26 22587
rect -20 22515 -14 22549
rect 20 22515 26 22549
rect -20 22477 26 22515
rect -20 22443 -14 22477
rect 20 22443 26 22477
rect -536 22371 -530 22405
rect -496 22371 -490 22405
rect -1052 22299 -1046 22333
rect -1012 22299 -1006 22333
rect -1052 22261 -1006 22299
rect -1270 22241 -1242 22250
rect -1332 22189 -1313 22241
rect -1261 22189 -1242 22241
rect -1332 22180 -1304 22189
rect -1568 22140 -1522 22155
rect -1310 22155 -1304 22180
rect -1270 22180 -1242 22189
rect -1052 22227 -1046 22261
rect -1012 22227 -1006 22261
rect -794 22333 -748 22360
rect -794 22299 -788 22333
rect -754 22299 -748 22333
rect -794 22261 -748 22299
rect -794 22250 -788 22261
rect -1052 22189 -1006 22227
rect -1270 22155 -1264 22180
rect -1310 22140 -1264 22155
rect -1052 22155 -1046 22189
rect -1012 22155 -1006 22189
rect -822 22241 -788 22250
rect -754 22250 -748 22261
rect -536 22333 -490 22371
rect -302 22421 -212 22430
rect -302 22369 -283 22421
rect -231 22369 -212 22421
rect -302 22360 -212 22369
rect -20 22405 26 22443
rect 238 22837 284 22875
rect 468 22911 558 22920
rect 468 22859 487 22911
rect 539 22859 558 22911
rect 468 22850 558 22859
rect 754 22909 800 22947
rect 1012 23019 1018 23030
rect 1052 23030 1078 23039
rect 1270 23091 1276 23125
rect 1310 23091 1316 23125
rect 1528 23125 1574 23140
rect 1528 23100 1534 23125
rect 1270 23053 1316 23091
rect 1052 23019 1058 23030
rect 1012 22981 1058 23019
rect 1012 22947 1018 22981
rect 1052 22947 1058 22981
rect 1012 22920 1058 22947
rect 1270 23019 1276 23053
rect 1310 23019 1316 23053
rect 1508 23091 1534 23100
rect 1568 23100 1574 23125
rect 1568 23091 1598 23100
rect 1508 23039 1527 23091
rect 1579 23039 1598 23091
rect 1508 23030 1534 23039
rect 1270 22981 1316 23019
rect 1270 22947 1276 22981
rect 1310 22947 1316 22981
rect 754 22875 760 22909
rect 794 22875 800 22909
rect 238 22803 244 22837
rect 278 22803 284 22837
rect 238 22765 284 22803
rect 238 22731 244 22765
rect 278 22731 284 22765
rect 238 22693 284 22731
rect 238 22659 244 22693
rect 278 22659 284 22693
rect 238 22621 284 22659
rect 238 22587 244 22621
rect 278 22587 284 22621
rect 238 22549 284 22587
rect 238 22515 244 22549
rect 278 22515 284 22549
rect 238 22477 284 22515
rect 238 22443 244 22477
rect 278 22443 284 22477
rect 238 22430 284 22443
rect 496 22837 542 22850
rect 496 22803 502 22837
rect 536 22803 542 22837
rect 496 22765 542 22803
rect 496 22731 502 22765
rect 536 22731 542 22765
rect 496 22693 542 22731
rect 496 22659 502 22693
rect 536 22659 542 22693
rect 496 22621 542 22659
rect 496 22587 502 22621
rect 536 22587 542 22621
rect 496 22549 542 22587
rect 496 22515 502 22549
rect 536 22515 542 22549
rect 496 22477 542 22515
rect 496 22443 502 22477
rect 536 22443 542 22477
rect -20 22371 -14 22405
rect 20 22371 26 22405
rect -536 22299 -530 22333
rect -496 22299 -490 22333
rect -536 22261 -490 22299
rect -754 22241 -732 22250
rect -822 22189 -803 22241
rect -751 22189 -732 22241
rect -822 22180 -788 22189
rect -1052 22140 -1006 22155
rect -794 22155 -788 22180
rect -754 22180 -732 22189
rect -536 22227 -530 22261
rect -496 22227 -490 22261
rect -278 22333 -232 22360
rect -278 22299 -272 22333
rect -238 22299 -232 22333
rect -278 22261 -232 22299
rect -278 22250 -272 22261
rect -536 22189 -490 22227
rect -754 22155 -748 22180
rect -794 22140 -748 22155
rect -536 22155 -530 22189
rect -496 22155 -490 22189
rect -302 22241 -272 22250
rect -238 22250 -232 22261
rect -20 22333 26 22371
rect 218 22421 308 22430
rect 218 22369 237 22421
rect 289 22369 308 22421
rect 218 22360 308 22369
rect 496 22405 542 22443
rect 754 22837 800 22875
rect 988 22911 1078 22920
rect 988 22859 1007 22911
rect 1059 22859 1078 22911
rect 988 22850 1078 22859
rect 1270 22909 1316 22947
rect 1528 23019 1534 23030
rect 1568 23030 1598 23039
rect 1568 23019 1574 23030
rect 1528 22981 1574 23019
rect 1528 22947 1534 22981
rect 1568 22947 1574 22981
rect 1528 22920 1574 22947
rect 1270 22875 1276 22909
rect 1310 22875 1316 22909
rect 754 22803 760 22837
rect 794 22803 800 22837
rect 754 22765 800 22803
rect 754 22731 760 22765
rect 794 22731 800 22765
rect 754 22693 800 22731
rect 754 22659 760 22693
rect 794 22659 800 22693
rect 754 22621 800 22659
rect 754 22587 760 22621
rect 794 22587 800 22621
rect 754 22549 800 22587
rect 754 22515 760 22549
rect 794 22515 800 22549
rect 754 22477 800 22515
rect 754 22443 760 22477
rect 794 22443 800 22477
rect 754 22430 800 22443
rect 1012 22837 1058 22850
rect 1012 22803 1018 22837
rect 1052 22803 1058 22837
rect 1012 22765 1058 22803
rect 1012 22731 1018 22765
rect 1052 22731 1058 22765
rect 1012 22693 1058 22731
rect 1012 22659 1018 22693
rect 1052 22659 1058 22693
rect 1012 22621 1058 22659
rect 1012 22587 1018 22621
rect 1052 22587 1058 22621
rect 1012 22549 1058 22587
rect 1012 22515 1018 22549
rect 1052 22515 1058 22549
rect 1012 22477 1058 22515
rect 1012 22443 1018 22477
rect 1052 22443 1058 22477
rect 496 22371 502 22405
rect 536 22371 542 22405
rect -20 22299 -14 22333
rect 20 22299 26 22333
rect -20 22261 26 22299
rect -238 22241 -212 22250
rect -302 22189 -283 22241
rect -231 22189 -212 22241
rect -302 22180 -272 22189
rect -536 22140 -490 22155
rect -278 22155 -272 22180
rect -238 22180 -212 22189
rect -20 22227 -14 22261
rect 20 22227 26 22261
rect 238 22333 284 22360
rect 238 22299 244 22333
rect 278 22299 284 22333
rect 238 22261 284 22299
rect 238 22250 244 22261
rect -20 22189 26 22227
rect -238 22155 -232 22180
rect -278 22140 -232 22155
rect -20 22155 -14 22189
rect 20 22155 26 22189
rect 218 22241 244 22250
rect 278 22250 284 22261
rect 496 22333 542 22371
rect 728 22421 818 22430
rect 728 22369 747 22421
rect 799 22369 818 22421
rect 728 22360 818 22369
rect 1012 22405 1058 22443
rect 1270 22837 1316 22875
rect 1508 22911 1598 22920
rect 1508 22859 1527 22911
rect 1579 22859 1598 22911
rect 1508 22850 1598 22859
rect 1270 22803 1276 22837
rect 1310 22803 1316 22837
rect 1270 22765 1316 22803
rect 1270 22731 1276 22765
rect 1310 22731 1316 22765
rect 1270 22693 1316 22731
rect 1270 22659 1276 22693
rect 1310 22659 1316 22693
rect 1270 22621 1316 22659
rect 1270 22587 1276 22621
rect 1310 22587 1316 22621
rect 1270 22549 1316 22587
rect 1270 22515 1276 22549
rect 1310 22515 1316 22549
rect 1270 22477 1316 22515
rect 1270 22443 1276 22477
rect 1310 22443 1316 22477
rect 1270 22430 1316 22443
rect 1528 22837 1574 22850
rect 1528 22803 1534 22837
rect 1568 22803 1574 22837
rect 1528 22765 1574 22803
rect 1528 22731 1534 22765
rect 1568 22731 1574 22765
rect 1528 22693 1574 22731
rect 1528 22659 1534 22693
rect 1568 22659 1574 22693
rect 1528 22621 1574 22659
rect 1528 22587 1534 22621
rect 1568 22587 1574 22621
rect 1528 22549 1574 22587
rect 1528 22515 1534 22549
rect 1568 22515 1574 22549
rect 1528 22477 1574 22515
rect 1528 22443 1534 22477
rect 1568 22443 1574 22477
rect 1012 22371 1018 22405
rect 1052 22371 1058 22405
rect 496 22299 502 22333
rect 536 22299 542 22333
rect 496 22261 542 22299
rect 278 22241 308 22250
rect 218 22189 237 22241
rect 289 22189 308 22241
rect 218 22180 244 22189
rect -20 22140 26 22155
rect 238 22155 244 22180
rect 278 22180 308 22189
rect 496 22227 502 22261
rect 536 22227 542 22261
rect 754 22333 800 22360
rect 754 22299 760 22333
rect 794 22299 800 22333
rect 754 22261 800 22299
rect 754 22250 760 22261
rect 496 22189 542 22227
rect 278 22155 284 22180
rect 238 22140 284 22155
rect 496 22155 502 22189
rect 536 22155 542 22189
rect 728 22241 760 22250
rect 794 22250 800 22261
rect 1012 22333 1058 22371
rect 1248 22421 1338 22430
rect 1248 22369 1267 22421
rect 1319 22369 1338 22421
rect 1248 22360 1338 22369
rect 1528 22405 1574 22443
rect 1528 22371 1534 22405
rect 1568 22371 1574 22405
rect 1012 22299 1018 22333
rect 1052 22299 1058 22333
rect 1012 22261 1058 22299
rect 794 22241 818 22250
rect 728 22189 747 22241
rect 799 22189 818 22241
rect 728 22180 760 22189
rect 496 22140 542 22155
rect 754 22155 760 22180
rect 794 22180 818 22189
rect 1012 22227 1018 22261
rect 1052 22227 1058 22261
rect 1270 22333 1316 22360
rect 1270 22299 1276 22333
rect 1310 22299 1316 22333
rect 1270 22261 1316 22299
rect 1270 22250 1276 22261
rect 1012 22189 1058 22227
rect 794 22155 800 22180
rect 754 22140 800 22155
rect 1012 22155 1018 22189
rect 1052 22155 1058 22189
rect 1248 22241 1276 22250
rect 1310 22250 1316 22261
rect 1528 22333 1574 22371
rect 1528 22299 1534 22333
rect 1568 22299 1574 22333
rect 1528 22261 1574 22299
rect 1310 22241 1338 22250
rect 1248 22189 1267 22241
rect 1319 22189 1338 22241
rect 1248 22180 1276 22189
rect 1012 22140 1058 22155
rect 1270 22155 1276 22180
rect 1310 22180 1338 22189
rect 1528 22227 1534 22261
rect 1568 22227 1574 22261
rect 1528 22189 1574 22227
rect 1310 22155 1316 22180
rect 1270 22140 1316 22155
rect 1528 22155 1534 22189
rect 1568 22155 1574 22189
rect 1528 22140 1574 22155
rect -2402 22111 -2272 22140
rect -2402 22110 -2363 22111
rect -2412 22060 -2363 22110
rect -2402 22059 -2363 22060
rect -2311 22110 -2272 22111
rect -2152 22111 -2022 22140
rect -2152 22110 -2113 22111
rect -2311 22060 -2113 22110
rect -2311 22059 -2272 22060
rect -2402 22030 -2272 22059
rect -2152 22059 -2113 22060
rect -2061 22110 -2022 22111
rect 1998 22111 2128 22140
rect 1998 22110 2037 22111
rect -2061 22102 2037 22110
rect -2061 22068 -1469 22102
rect -1435 22068 -1397 22102
rect -1363 22068 -1211 22102
rect -1177 22068 -1139 22102
rect -1105 22068 -953 22102
rect -919 22068 -881 22102
rect -847 22068 -695 22102
rect -661 22068 -623 22102
rect -589 22068 -437 22102
rect -403 22068 -365 22102
rect -331 22068 -179 22102
rect -145 22068 -107 22102
rect -73 22068 79 22102
rect 113 22068 151 22102
rect 185 22068 337 22102
rect 371 22068 409 22102
rect 443 22068 595 22102
rect 629 22068 667 22102
rect 701 22068 853 22102
rect 887 22068 925 22102
rect 959 22068 1111 22102
rect 1145 22068 1183 22102
rect 1217 22068 1369 22102
rect 1403 22068 1441 22102
rect 1475 22068 2037 22102
rect -2061 22060 2037 22068
rect -2061 22059 -2022 22060
rect -2152 22030 -2022 22059
rect 1998 22059 2037 22060
rect 2089 22110 2128 22111
rect 2248 22111 2378 22140
rect 2248 22110 2287 22111
rect 2089 22060 2287 22110
rect 2089 22059 2128 22060
rect 1998 22030 2128 22059
rect 2248 22059 2287 22060
rect 2339 22110 2378 22111
rect 2339 22060 2388 22110
rect 2339 22059 2378 22060
rect 2248 22030 2378 22059
rect -132 22007 138 22010
rect -132 22006 -119 22007
rect -831 22000 -119 22006
rect 125 22006 138 22007
rect 125 22000 837 22006
rect -831 21966 -806 22000
rect -772 21966 -734 22000
rect -700 21966 -662 22000
rect -628 21966 -590 22000
rect -556 21966 -518 22000
rect -484 21966 -446 22000
rect -412 21966 -374 22000
rect -340 21966 -302 22000
rect -268 21966 -230 22000
rect -196 21966 -158 22000
rect -124 21966 -119 22000
rect 125 21966 130 22000
rect 164 21966 202 22000
rect 236 21966 274 22000
rect 308 21966 346 22000
rect 380 21966 418 22000
rect 452 21966 490 22000
rect 524 21966 562 22000
rect 596 21966 634 22000
rect 668 21966 706 22000
rect 740 21966 778 22000
rect 812 21966 837 22000
rect -831 21960 -119 21966
rect -132 21800 -119 21960
rect -962 21794 -119 21800
rect 125 21960 837 21966
rect 125 21800 138 21960
rect 125 21794 964 21800
rect -962 21760 -916 21794
rect -882 21760 -844 21794
rect -810 21760 -772 21794
rect -738 21760 -700 21794
rect -666 21760 -628 21794
rect -594 21760 -556 21794
rect -522 21760 -484 21794
rect -450 21760 -412 21794
rect -378 21760 -340 21794
rect -306 21760 -268 21794
rect -234 21760 -196 21794
rect -162 21760 -124 21794
rect -90 21760 -52 21763
rect -18 21760 20 21763
rect 54 21760 92 21763
rect 126 21760 164 21794
rect 198 21760 236 21794
rect 270 21760 308 21794
rect 342 21760 380 21794
rect 414 21760 452 21794
rect 486 21760 524 21794
rect 558 21760 596 21794
rect 630 21760 668 21794
rect 702 21760 740 21794
rect 774 21760 812 21794
rect 846 21760 884 21794
rect 918 21760 964 21794
rect 5418 21780 6328 29120
rect -6370 21716 -2662 21760
rect -962 21754 964 21760
rect -132 21750 138 21754
rect -6370 21344 -3249 21716
rect -2685 21344 -2662 21716
rect -2402 21701 -2272 21730
rect -2402 21700 -2363 21701
rect -2412 21650 -2363 21700
rect -2402 21649 -2363 21650
rect -2311 21700 -2272 21701
rect -2152 21701 -2022 21730
rect -2152 21700 -2113 21701
rect -2311 21650 -2113 21700
rect -2311 21649 -2272 21650
rect -2402 21620 -2272 21649
rect -2152 21649 -2113 21650
rect -2061 21700 -2022 21701
rect 1998 21701 2128 21730
rect 1998 21700 2037 21701
rect -2061 21692 2037 21700
rect -2061 21658 -1729 21692
rect -1695 21658 -1657 21692
rect -1623 21658 -1471 21692
rect -1437 21658 -1399 21692
rect -1365 21658 -1213 21692
rect -1179 21658 -1141 21692
rect -1107 21658 -955 21692
rect -921 21658 -883 21692
rect -849 21658 -697 21692
rect -663 21658 -625 21692
rect -591 21658 -439 21692
rect -405 21658 -367 21692
rect -333 21658 -181 21692
rect -147 21658 -109 21692
rect -75 21658 77 21692
rect 111 21658 149 21692
rect 183 21658 335 21692
rect 369 21658 407 21692
rect 441 21658 593 21692
rect 627 21658 665 21692
rect 699 21658 851 21692
rect 885 21658 923 21692
rect 957 21658 1109 21692
rect 1143 21658 1181 21692
rect 1215 21658 1367 21692
rect 1401 21658 1439 21692
rect 1473 21658 1625 21692
rect 1659 21658 1697 21692
rect 1731 21658 2037 21692
rect -2061 21650 2037 21658
rect -2061 21649 -2022 21650
rect -2152 21620 -2022 21649
rect 1998 21649 2037 21650
rect 2089 21700 2128 21701
rect 2248 21701 2378 21730
rect 2248 21700 2287 21701
rect 2089 21650 2287 21700
rect 2089 21649 2128 21650
rect 1998 21620 2128 21649
rect 2248 21649 2287 21650
rect 2339 21700 2378 21701
rect 2339 21650 2388 21700
rect 2588 21680 6328 21780
rect 2339 21649 2378 21650
rect 2248 21620 2378 21649
rect -1828 21605 -1782 21620
rect -1828 21580 -1822 21605
rect -1852 21571 -1822 21580
rect -1788 21580 -1782 21605
rect -1570 21605 -1524 21620
rect -1788 21571 -1762 21580
rect -1852 21519 -1833 21571
rect -1781 21519 -1762 21571
rect -1852 21510 -1822 21519
rect -1828 21499 -1822 21510
rect -1788 21510 -1762 21519
rect -1570 21571 -1564 21605
rect -1530 21571 -1524 21605
rect -1312 21605 -1266 21620
rect -1312 21580 -1306 21605
rect -1570 21533 -1524 21571
rect -1788 21499 -1782 21510
rect -1828 21461 -1782 21499
rect -1828 21427 -1822 21461
rect -1788 21427 -1782 21461
rect -1828 21400 -1782 21427
rect -1570 21499 -1564 21533
rect -1530 21499 -1524 21533
rect -1332 21571 -1306 21580
rect -1272 21580 -1266 21605
rect -1054 21605 -1008 21620
rect -1272 21571 -1242 21580
rect -1332 21519 -1313 21571
rect -1261 21519 -1242 21571
rect -1332 21510 -1306 21519
rect -1570 21461 -1524 21499
rect -1570 21427 -1564 21461
rect -1530 21427 -1524 21461
rect -6370 21310 -2662 21344
rect -1852 21391 -1762 21400
rect -1852 21339 -1833 21391
rect -1781 21339 -1762 21391
rect -1852 21330 -1762 21339
rect -1570 21389 -1524 21427
rect -1312 21499 -1306 21510
rect -1272 21510 -1242 21519
rect -1054 21571 -1048 21605
rect -1014 21571 -1008 21605
rect -796 21605 -750 21620
rect -796 21580 -790 21605
rect -1054 21533 -1008 21571
rect -1272 21499 -1266 21510
rect -1312 21461 -1266 21499
rect -1312 21427 -1306 21461
rect -1272 21427 -1266 21461
rect -1312 21400 -1266 21427
rect -1054 21499 -1048 21533
rect -1014 21499 -1008 21533
rect -822 21571 -790 21580
rect -756 21580 -750 21605
rect -538 21605 -492 21620
rect -756 21571 -732 21580
rect -822 21519 -803 21571
rect -751 21519 -732 21571
rect -822 21510 -790 21519
rect -1054 21461 -1008 21499
rect -1054 21427 -1048 21461
rect -1014 21427 -1008 21461
rect -1570 21355 -1564 21389
rect -1530 21355 -1524 21389
rect -1828 21317 -1782 21330
rect -1828 21283 -1822 21317
rect -1788 21283 -1782 21317
rect -1828 21245 -1782 21283
rect -1828 21211 -1822 21245
rect -1788 21211 -1782 21245
rect -1828 21173 -1782 21211
rect -1828 21139 -1822 21173
rect -1788 21139 -1782 21173
rect -1828 21101 -1782 21139
rect -1828 21067 -1822 21101
rect -1788 21067 -1782 21101
rect -1828 21029 -1782 21067
rect -1828 20995 -1822 21029
rect -1788 20995 -1782 21029
rect -1828 20957 -1782 20995
rect -1828 20923 -1822 20957
rect -1788 20923 -1782 20957
rect -1828 20885 -1782 20923
rect -1570 21317 -1524 21355
rect -1332 21391 -1242 21400
rect -1332 21339 -1313 21391
rect -1261 21339 -1242 21391
rect -1332 21330 -1242 21339
rect -1054 21389 -1008 21427
rect -796 21499 -790 21510
rect -756 21510 -732 21519
rect -538 21571 -532 21605
rect -498 21571 -492 21605
rect -280 21605 -234 21620
rect -280 21580 -274 21605
rect -538 21533 -492 21571
rect -756 21499 -750 21510
rect -796 21461 -750 21499
rect -796 21427 -790 21461
rect -756 21427 -750 21461
rect -796 21400 -750 21427
rect -538 21499 -532 21533
rect -498 21499 -492 21533
rect -302 21571 -274 21580
rect -240 21580 -234 21605
rect -22 21605 24 21620
rect -240 21571 -212 21580
rect -302 21519 -283 21571
rect -231 21519 -212 21571
rect -302 21510 -274 21519
rect -538 21461 -492 21499
rect -538 21427 -532 21461
rect -498 21427 -492 21461
rect -1054 21355 -1048 21389
rect -1014 21355 -1008 21389
rect -1570 21283 -1564 21317
rect -1530 21283 -1524 21317
rect -1570 21245 -1524 21283
rect -1570 21211 -1564 21245
rect -1530 21211 -1524 21245
rect -1570 21173 -1524 21211
rect -1570 21139 -1564 21173
rect -1530 21139 -1524 21173
rect -1570 21101 -1524 21139
rect -1570 21067 -1564 21101
rect -1530 21067 -1524 21101
rect -1570 21029 -1524 21067
rect -1570 20995 -1564 21029
rect -1530 20995 -1524 21029
rect -1570 20957 -1524 20995
rect -1570 20923 -1564 20957
rect -1530 20923 -1524 20957
rect -1570 20910 -1524 20923
rect -1312 21317 -1266 21330
rect -1312 21283 -1306 21317
rect -1272 21283 -1266 21317
rect -1312 21245 -1266 21283
rect -1312 21211 -1306 21245
rect -1272 21211 -1266 21245
rect -1312 21173 -1266 21211
rect -1312 21139 -1306 21173
rect -1272 21139 -1266 21173
rect -1312 21101 -1266 21139
rect -1312 21067 -1306 21101
rect -1272 21067 -1266 21101
rect -1312 21029 -1266 21067
rect -1312 20995 -1306 21029
rect -1272 20995 -1266 21029
rect -1312 20957 -1266 20995
rect -1312 20923 -1306 20957
rect -1272 20923 -1266 20957
rect -1828 20851 -1822 20885
rect -1788 20851 -1782 20885
rect -1828 20813 -1782 20851
rect -1592 20901 -1502 20910
rect -1592 20849 -1573 20901
rect -1521 20849 -1502 20901
rect -1592 20840 -1502 20849
rect -1312 20885 -1266 20923
rect -1054 21317 -1008 21355
rect -822 21391 -732 21400
rect -822 21339 -803 21391
rect -751 21339 -732 21391
rect -822 21330 -732 21339
rect -538 21389 -492 21427
rect -280 21499 -274 21510
rect -240 21510 -212 21519
rect -22 21571 -16 21605
rect 18 21571 24 21605
rect 236 21605 282 21620
rect 236 21580 242 21605
rect -22 21533 24 21571
rect -240 21499 -234 21510
rect -280 21461 -234 21499
rect -280 21427 -274 21461
rect -240 21427 -234 21461
rect -280 21400 -234 21427
rect -22 21499 -16 21533
rect 18 21499 24 21533
rect 208 21571 242 21580
rect 276 21580 282 21605
rect 494 21605 540 21620
rect 276 21571 298 21580
rect 208 21519 227 21571
rect 279 21519 298 21571
rect 208 21510 242 21519
rect -22 21461 24 21499
rect -22 21427 -16 21461
rect 18 21427 24 21461
rect -538 21355 -532 21389
rect -498 21355 -492 21389
rect -1054 21283 -1048 21317
rect -1014 21283 -1008 21317
rect -1054 21245 -1008 21283
rect -1054 21211 -1048 21245
rect -1014 21211 -1008 21245
rect -1054 21173 -1008 21211
rect -1054 21139 -1048 21173
rect -1014 21139 -1008 21173
rect -1054 21101 -1008 21139
rect -1054 21067 -1048 21101
rect -1014 21067 -1008 21101
rect -1054 21029 -1008 21067
rect -1054 20995 -1048 21029
rect -1014 20995 -1008 21029
rect -1054 20957 -1008 20995
rect -1054 20923 -1048 20957
rect -1014 20923 -1008 20957
rect -1054 20910 -1008 20923
rect -796 21317 -750 21330
rect -796 21283 -790 21317
rect -756 21283 -750 21317
rect -796 21245 -750 21283
rect -796 21211 -790 21245
rect -756 21211 -750 21245
rect -796 21173 -750 21211
rect -796 21139 -790 21173
rect -756 21139 -750 21173
rect -796 21101 -750 21139
rect -796 21067 -790 21101
rect -756 21067 -750 21101
rect -796 21029 -750 21067
rect -796 20995 -790 21029
rect -756 20995 -750 21029
rect -796 20957 -750 20995
rect -796 20923 -790 20957
rect -756 20923 -750 20957
rect -1312 20851 -1306 20885
rect -1272 20851 -1266 20885
rect -1828 20779 -1822 20813
rect -1788 20779 -1782 20813
rect -1828 20741 -1782 20779
rect -1828 20707 -1822 20741
rect -1788 20707 -1782 20741
rect -1570 20813 -1524 20840
rect -1570 20779 -1564 20813
rect -1530 20779 -1524 20813
rect -1570 20741 -1524 20779
rect -1570 20730 -1564 20741
rect -1828 20669 -1782 20707
rect -1828 20635 -1822 20669
rect -1788 20635 -1782 20669
rect -1592 20721 -1564 20730
rect -1530 20730 -1524 20741
rect -1312 20813 -1266 20851
rect -1082 20901 -992 20910
rect -1082 20849 -1063 20901
rect -1011 20849 -992 20901
rect -1082 20840 -992 20849
rect -796 20885 -750 20923
rect -538 21317 -492 21355
rect -302 21391 -212 21400
rect -302 21339 -283 21391
rect -231 21339 -212 21391
rect -302 21330 -212 21339
rect -22 21389 24 21427
rect 236 21499 242 21510
rect 276 21510 298 21519
rect 494 21571 500 21605
rect 534 21571 540 21605
rect 752 21605 798 21620
rect 752 21580 758 21605
rect 494 21533 540 21571
rect 276 21499 282 21510
rect 236 21461 282 21499
rect 236 21427 242 21461
rect 276 21427 282 21461
rect 236 21400 282 21427
rect 494 21499 500 21533
rect 534 21499 540 21533
rect 728 21571 758 21580
rect 792 21580 798 21605
rect 1010 21605 1056 21620
rect 792 21571 818 21580
rect 728 21519 747 21571
rect 799 21519 818 21571
rect 728 21510 758 21519
rect 494 21461 540 21499
rect 494 21427 500 21461
rect 534 21427 540 21461
rect -22 21355 -16 21389
rect 18 21355 24 21389
rect -538 21283 -532 21317
rect -498 21283 -492 21317
rect -538 21245 -492 21283
rect -538 21211 -532 21245
rect -498 21211 -492 21245
rect -538 21173 -492 21211
rect -538 21139 -532 21173
rect -498 21139 -492 21173
rect -538 21101 -492 21139
rect -538 21067 -532 21101
rect -498 21067 -492 21101
rect -538 21029 -492 21067
rect -538 20995 -532 21029
rect -498 20995 -492 21029
rect -538 20957 -492 20995
rect -538 20923 -532 20957
rect -498 20923 -492 20957
rect -538 20910 -492 20923
rect -280 21317 -234 21330
rect -280 21283 -274 21317
rect -240 21283 -234 21317
rect -280 21245 -234 21283
rect -280 21211 -274 21245
rect -240 21211 -234 21245
rect -280 21173 -234 21211
rect -280 21139 -274 21173
rect -240 21139 -234 21173
rect -280 21101 -234 21139
rect -280 21067 -274 21101
rect -240 21067 -234 21101
rect -280 21029 -234 21067
rect -280 20995 -274 21029
rect -240 20995 -234 21029
rect -280 20957 -234 20995
rect -280 20923 -274 20957
rect -240 20923 -234 20957
rect -796 20851 -790 20885
rect -756 20851 -750 20885
rect -1312 20779 -1306 20813
rect -1272 20779 -1266 20813
rect -1312 20741 -1266 20779
rect -1530 20721 -1502 20730
rect -1592 20669 -1573 20721
rect -1521 20669 -1502 20721
rect -1592 20660 -1564 20669
rect -1828 20620 -1782 20635
rect -1570 20635 -1564 20660
rect -1530 20660 -1502 20669
rect -1312 20707 -1306 20741
rect -1272 20707 -1266 20741
rect -1054 20813 -1008 20840
rect -1054 20779 -1048 20813
rect -1014 20779 -1008 20813
rect -1054 20741 -1008 20779
rect -1054 20730 -1048 20741
rect -1312 20669 -1266 20707
rect -1530 20635 -1524 20660
rect -1570 20620 -1524 20635
rect -1312 20635 -1306 20669
rect -1272 20635 -1266 20669
rect -1082 20721 -1048 20730
rect -1014 20730 -1008 20741
rect -796 20813 -750 20851
rect -562 20901 -472 20910
rect -562 20849 -543 20901
rect -491 20849 -472 20901
rect -562 20840 -472 20849
rect -280 20885 -234 20923
rect -22 21317 24 21355
rect 208 21391 298 21400
rect 208 21339 227 21391
rect 279 21339 298 21391
rect 208 21330 298 21339
rect 494 21389 540 21427
rect 752 21499 758 21510
rect 792 21510 818 21519
rect 1010 21571 1016 21605
rect 1050 21571 1056 21605
rect 1268 21605 1314 21620
rect 1268 21580 1274 21605
rect 1010 21533 1056 21571
rect 792 21499 798 21510
rect 752 21461 798 21499
rect 752 21427 758 21461
rect 792 21427 798 21461
rect 752 21400 798 21427
rect 1010 21499 1016 21533
rect 1050 21499 1056 21533
rect 1248 21571 1274 21580
rect 1308 21580 1314 21605
rect 1526 21605 1572 21620
rect 1308 21571 1338 21580
rect 1248 21519 1267 21571
rect 1319 21519 1338 21571
rect 1248 21510 1274 21519
rect 1010 21461 1056 21499
rect 1010 21427 1016 21461
rect 1050 21427 1056 21461
rect 494 21355 500 21389
rect 534 21355 540 21389
rect -22 21283 -16 21317
rect 18 21283 24 21317
rect -22 21245 24 21283
rect -22 21211 -16 21245
rect 18 21211 24 21245
rect -22 21173 24 21211
rect -22 21139 -16 21173
rect 18 21139 24 21173
rect -22 21101 24 21139
rect -22 21067 -16 21101
rect 18 21067 24 21101
rect -22 21029 24 21067
rect -22 20995 -16 21029
rect 18 20995 24 21029
rect -22 20957 24 20995
rect -22 20923 -16 20957
rect 18 20923 24 20957
rect -22 20910 24 20923
rect 236 21317 282 21330
rect 236 21283 242 21317
rect 276 21283 282 21317
rect 236 21245 282 21283
rect 236 21211 242 21245
rect 276 21211 282 21245
rect 236 21173 282 21211
rect 236 21139 242 21173
rect 276 21139 282 21173
rect 236 21101 282 21139
rect 236 21067 242 21101
rect 276 21067 282 21101
rect 236 21029 282 21067
rect 236 20995 242 21029
rect 276 20995 282 21029
rect 236 20957 282 20995
rect 236 20923 242 20957
rect 276 20923 282 20957
rect -280 20851 -274 20885
rect -240 20851 -234 20885
rect -796 20779 -790 20813
rect -756 20779 -750 20813
rect -796 20741 -750 20779
rect -1014 20721 -992 20730
rect -1082 20669 -1063 20721
rect -1011 20669 -992 20721
rect -1082 20660 -1048 20669
rect -1312 20620 -1266 20635
rect -1054 20635 -1048 20660
rect -1014 20660 -992 20669
rect -796 20707 -790 20741
rect -756 20707 -750 20741
rect -538 20813 -492 20840
rect -538 20779 -532 20813
rect -498 20779 -492 20813
rect -538 20741 -492 20779
rect -538 20730 -532 20741
rect -796 20669 -750 20707
rect -1014 20635 -1008 20660
rect -1054 20620 -1008 20635
rect -796 20635 -790 20669
rect -756 20635 -750 20669
rect -562 20721 -532 20730
rect -498 20730 -492 20741
rect -280 20813 -234 20851
rect -42 20901 48 20910
rect -42 20849 -23 20901
rect 29 20849 48 20901
rect -42 20840 48 20849
rect 236 20885 282 20923
rect 494 21317 540 21355
rect 728 21391 818 21400
rect 728 21339 747 21391
rect 799 21339 818 21391
rect 728 21330 818 21339
rect 1010 21389 1056 21427
rect 1268 21499 1274 21510
rect 1308 21510 1338 21519
rect 1526 21571 1532 21605
rect 1566 21571 1572 21605
rect 1784 21605 1830 21620
rect 1784 21580 1790 21605
rect 1526 21533 1572 21571
rect 1308 21499 1314 21510
rect 1268 21461 1314 21499
rect 1268 21427 1274 21461
rect 1308 21427 1314 21461
rect 1268 21400 1314 21427
rect 1526 21499 1532 21533
rect 1566 21499 1572 21533
rect 1758 21571 1790 21580
rect 1824 21580 1830 21605
rect 1824 21571 1848 21580
rect 1758 21519 1777 21571
rect 1829 21519 1848 21571
rect 1758 21510 1790 21519
rect 1526 21461 1572 21499
rect 1526 21427 1532 21461
rect 1566 21427 1572 21461
rect 1010 21355 1016 21389
rect 1050 21355 1056 21389
rect 494 21283 500 21317
rect 534 21283 540 21317
rect 494 21245 540 21283
rect 494 21211 500 21245
rect 534 21211 540 21245
rect 494 21173 540 21211
rect 494 21139 500 21173
rect 534 21139 540 21173
rect 494 21101 540 21139
rect 494 21067 500 21101
rect 534 21067 540 21101
rect 494 21029 540 21067
rect 494 20995 500 21029
rect 534 20995 540 21029
rect 494 20957 540 20995
rect 494 20923 500 20957
rect 534 20923 540 20957
rect 494 20910 540 20923
rect 752 21317 798 21330
rect 752 21283 758 21317
rect 792 21283 798 21317
rect 752 21245 798 21283
rect 752 21211 758 21245
rect 792 21211 798 21245
rect 752 21173 798 21211
rect 752 21139 758 21173
rect 792 21139 798 21173
rect 752 21101 798 21139
rect 752 21067 758 21101
rect 792 21067 798 21101
rect 752 21029 798 21067
rect 752 20995 758 21029
rect 792 20995 798 21029
rect 752 20957 798 20995
rect 752 20923 758 20957
rect 792 20923 798 20957
rect 236 20851 242 20885
rect 276 20851 282 20885
rect -280 20779 -274 20813
rect -240 20779 -234 20813
rect -280 20741 -234 20779
rect -498 20721 -472 20730
rect -562 20669 -543 20721
rect -491 20669 -472 20721
rect -562 20660 -532 20669
rect -796 20620 -750 20635
rect -538 20635 -532 20660
rect -498 20660 -472 20669
rect -280 20707 -274 20741
rect -240 20707 -234 20741
rect -22 20813 24 20840
rect -22 20779 -16 20813
rect 18 20779 24 20813
rect -22 20741 24 20779
rect -22 20730 -16 20741
rect -280 20669 -234 20707
rect -498 20635 -492 20660
rect -538 20620 -492 20635
rect -280 20635 -274 20669
rect -240 20635 -234 20669
rect -42 20721 -16 20730
rect 18 20730 24 20741
rect 236 20813 282 20851
rect 468 20901 558 20910
rect 468 20849 487 20901
rect 539 20849 558 20901
rect 468 20840 558 20849
rect 752 20885 798 20923
rect 1010 21317 1056 21355
rect 1248 21391 1338 21400
rect 1248 21339 1267 21391
rect 1319 21339 1338 21391
rect 1248 21330 1338 21339
rect 1526 21389 1572 21427
rect 1784 21499 1790 21510
rect 1824 21510 1848 21519
rect 1824 21499 1830 21510
rect 1784 21461 1830 21499
rect 1784 21427 1790 21461
rect 1824 21427 1830 21461
rect 1784 21400 1830 21427
rect 2588 21440 2638 21680
rect 2878 21440 2968 21680
rect 3208 21440 6328 21680
rect 1526 21355 1532 21389
rect 1566 21355 1572 21389
rect 1010 21283 1016 21317
rect 1050 21283 1056 21317
rect 1010 21245 1056 21283
rect 1010 21211 1016 21245
rect 1050 21211 1056 21245
rect 1010 21173 1056 21211
rect 1010 21139 1016 21173
rect 1050 21139 1056 21173
rect 1010 21101 1056 21139
rect 1010 21067 1016 21101
rect 1050 21067 1056 21101
rect 1010 21029 1056 21067
rect 1010 20995 1016 21029
rect 1050 20995 1056 21029
rect 1010 20957 1056 20995
rect 1010 20923 1016 20957
rect 1050 20923 1056 20957
rect 1010 20910 1056 20923
rect 1268 21317 1314 21330
rect 1268 21283 1274 21317
rect 1308 21283 1314 21317
rect 1268 21245 1314 21283
rect 1268 21211 1274 21245
rect 1308 21211 1314 21245
rect 1268 21173 1314 21211
rect 1268 21139 1274 21173
rect 1308 21139 1314 21173
rect 1268 21101 1314 21139
rect 1268 21067 1274 21101
rect 1308 21067 1314 21101
rect 1268 21029 1314 21067
rect 1268 20995 1274 21029
rect 1308 20995 1314 21029
rect 1268 20957 1314 20995
rect 1268 20923 1274 20957
rect 1308 20923 1314 20957
rect 752 20851 758 20885
rect 792 20851 798 20885
rect 236 20779 242 20813
rect 276 20779 282 20813
rect 236 20741 282 20779
rect 18 20721 48 20730
rect -42 20669 -23 20721
rect 29 20669 48 20721
rect -42 20660 -16 20669
rect -280 20620 -234 20635
rect -22 20635 -16 20660
rect 18 20660 48 20669
rect 236 20707 242 20741
rect 276 20707 282 20741
rect 494 20813 540 20840
rect 494 20779 500 20813
rect 534 20779 540 20813
rect 494 20741 540 20779
rect 494 20730 500 20741
rect 236 20669 282 20707
rect 18 20635 24 20660
rect -22 20620 24 20635
rect 236 20635 242 20669
rect 276 20635 282 20669
rect 468 20721 500 20730
rect 534 20730 540 20741
rect 752 20813 798 20851
rect 988 20901 1078 20910
rect 988 20849 1007 20901
rect 1059 20849 1078 20901
rect 988 20840 1078 20849
rect 1268 20885 1314 20923
rect 1526 21317 1572 21355
rect 1758 21391 1848 21400
rect 1758 21339 1777 21391
rect 1829 21339 1848 21391
rect 1758 21330 1848 21339
rect 2588 21330 6328 21440
rect 1526 21283 1532 21317
rect 1566 21283 1572 21317
rect 1526 21245 1572 21283
rect 1526 21211 1532 21245
rect 1566 21211 1572 21245
rect 1526 21173 1572 21211
rect 1526 21139 1532 21173
rect 1566 21139 1572 21173
rect 1526 21101 1572 21139
rect 1526 21067 1532 21101
rect 1566 21067 1572 21101
rect 1526 21029 1572 21067
rect 1526 20995 1532 21029
rect 1566 20995 1572 21029
rect 1526 20957 1572 20995
rect 1526 20923 1532 20957
rect 1566 20923 1572 20957
rect 1526 20910 1572 20923
rect 1784 21317 1830 21330
rect 1784 21283 1790 21317
rect 1824 21283 1830 21317
rect 1784 21245 1830 21283
rect 1784 21211 1790 21245
rect 1824 21211 1830 21245
rect 1784 21173 1830 21211
rect 1784 21139 1790 21173
rect 1824 21139 1830 21173
rect 1784 21101 1830 21139
rect 1784 21067 1790 21101
rect 1824 21067 1830 21101
rect 1784 21029 1830 21067
rect 1784 20995 1790 21029
rect 1824 20995 1830 21029
rect 1784 20957 1830 20995
rect 1784 20923 1790 20957
rect 1824 20923 1830 20957
rect 1268 20851 1274 20885
rect 1308 20851 1314 20885
rect 752 20779 758 20813
rect 792 20779 798 20813
rect 752 20741 798 20779
rect 534 20721 558 20730
rect 468 20669 487 20721
rect 539 20669 558 20721
rect 468 20660 500 20669
rect 236 20620 282 20635
rect 494 20635 500 20660
rect 534 20660 558 20669
rect 752 20707 758 20741
rect 792 20707 798 20741
rect 1010 20813 1056 20840
rect 1010 20779 1016 20813
rect 1050 20779 1056 20813
rect 1010 20741 1056 20779
rect 1010 20730 1016 20741
rect 752 20669 798 20707
rect 534 20635 540 20660
rect 494 20620 540 20635
rect 752 20635 758 20669
rect 792 20635 798 20669
rect 988 20721 1016 20730
rect 1050 20730 1056 20741
rect 1268 20813 1314 20851
rect 1498 20901 1588 20910
rect 1498 20849 1517 20901
rect 1569 20849 1588 20901
rect 1498 20840 1588 20849
rect 1784 20885 1830 20923
rect 1784 20851 1790 20885
rect 1824 20851 1830 20885
rect 1268 20779 1274 20813
rect 1308 20779 1314 20813
rect 1268 20741 1314 20779
rect 1050 20721 1078 20730
rect 988 20669 1007 20721
rect 1059 20669 1078 20721
rect 988 20660 1016 20669
rect 752 20620 798 20635
rect 1010 20635 1016 20660
rect 1050 20660 1078 20669
rect 1268 20707 1274 20741
rect 1308 20707 1314 20741
rect 1526 20813 1572 20840
rect 1526 20779 1532 20813
rect 1566 20779 1572 20813
rect 1526 20741 1572 20779
rect 1526 20730 1532 20741
rect 1268 20669 1314 20707
rect 1050 20635 1056 20660
rect 1010 20620 1056 20635
rect 1268 20635 1274 20669
rect 1308 20635 1314 20669
rect 1498 20721 1532 20730
rect 1566 20730 1572 20741
rect 1784 20813 1830 20851
rect 1784 20779 1790 20813
rect 1824 20779 1830 20813
rect 1784 20741 1830 20779
rect 1566 20721 1588 20730
rect 1498 20669 1517 20721
rect 1569 20669 1588 20721
rect 1498 20660 1532 20669
rect 1268 20620 1314 20635
rect 1526 20635 1532 20660
rect 1566 20660 1588 20669
rect 1784 20707 1790 20741
rect 1824 20707 1830 20741
rect 1784 20669 1830 20707
rect 1566 20635 1572 20660
rect 1526 20620 1572 20635
rect 1784 20635 1790 20669
rect 1824 20635 1830 20669
rect 1784 20620 1830 20635
rect -2402 20591 -2272 20620
rect -2402 20590 -2363 20591
rect -2412 20540 -2363 20590
rect -2402 20539 -2363 20540
rect -2311 20590 -2272 20591
rect -2152 20591 -2022 20620
rect -2152 20590 -2113 20591
rect -2311 20540 -2113 20590
rect -2311 20539 -2272 20540
rect -2402 20510 -2272 20539
rect -2152 20539 -2113 20540
rect -2061 20590 -2022 20591
rect 1998 20591 2128 20620
rect 1998 20590 2037 20591
rect -2061 20582 2037 20590
rect -2061 20548 -1729 20582
rect -1695 20548 -1657 20582
rect -1623 20548 -1471 20582
rect -1437 20548 -1399 20582
rect -1365 20548 -1213 20582
rect -1179 20548 -1141 20582
rect -1107 20548 -955 20582
rect -921 20548 -883 20582
rect -849 20548 -697 20582
rect -663 20548 -625 20582
rect -591 20548 -439 20582
rect -405 20548 -367 20582
rect -333 20548 -181 20582
rect -147 20548 -109 20582
rect -75 20548 77 20582
rect 111 20548 149 20582
rect 183 20548 335 20582
rect 369 20548 407 20582
rect 441 20548 593 20582
rect 627 20548 665 20582
rect 699 20548 851 20582
rect 885 20548 923 20582
rect 957 20548 1109 20582
rect 1143 20548 1181 20582
rect 1215 20548 1367 20582
rect 1401 20548 1439 20582
rect 1473 20548 1625 20582
rect 1659 20548 1697 20582
rect 1731 20548 2037 20582
rect -2061 20540 2037 20548
rect -2061 20539 -2022 20540
rect -2152 20510 -2022 20539
rect 1998 20539 2037 20540
rect 2089 20590 2128 20591
rect 2248 20591 2378 20620
rect 2248 20590 2287 20591
rect 2089 20540 2287 20590
rect 2089 20539 2128 20540
rect 1998 20510 2128 20539
rect 2248 20539 2287 20540
rect 2339 20590 2378 20591
rect 2339 20540 2388 20590
rect 2339 20539 2378 20540
rect 2248 20510 2378 20539
rect -962 20480 964 20486
rect -962 20446 -916 20480
rect -882 20446 -844 20480
rect -810 20446 -772 20480
rect -738 20446 -700 20480
rect -666 20446 -628 20480
rect -594 20446 -556 20480
rect -522 20446 -484 20480
rect -450 20446 -412 20480
rect -378 20446 -340 20480
rect -306 20446 -268 20480
rect -234 20446 -196 20480
rect -162 20446 -124 20480
rect -90 20477 -52 20480
rect -18 20477 20 20480
rect 54 20477 92 20480
rect 126 20446 164 20480
rect 198 20446 236 20480
rect 270 20446 308 20480
rect 342 20446 380 20480
rect 414 20446 452 20480
rect 486 20446 524 20480
rect 558 20446 596 20480
rect 630 20446 668 20480
rect 702 20446 740 20480
rect 774 20446 812 20480
rect 846 20446 884 20480
rect 918 20446 964 20480
rect -962 20440 -119 20446
rect -132 20233 -119 20440
rect 125 20440 964 20446
rect 125 20233 138 20440
rect -132 20230 138 20233
rect -3232 19640 -3048 19646
rect -2172 19640 -1988 19646
rect -712 19640 -528 19646
rect 508 19640 692 19646
rect 1988 19640 2172 19646
rect 2988 19640 3172 19646
rect -3600 19480 -3220 19640
rect -3060 19480 -2160 19640
rect -2000 19480 -700 19640
rect -540 19480 520 19640
rect 680 19480 2000 19640
rect 2160 19480 3000 19640
rect 3160 19480 3600 19640
rect -3600 19432 3600 19480
rect -3600 19398 -3579 19432
rect -2603 19420 -2343 19432
rect -2603 19398 -2580 19420
rect -3678 19370 -3632 19382
rect -3600 19380 -2580 19398
rect -2360 19398 -2343 19420
rect -1367 19420 -1107 19432
rect -1367 19398 -1355 19420
rect -2360 19392 -1355 19398
rect -1120 19398 -1107 19420
rect -131 19420 129 19432
rect -131 19398 -119 19420
rect -1120 19392 -119 19398
rect 117 19398 129 19420
rect 1105 19420 1365 19432
rect 1105 19398 1120 19420
rect 117 19392 1120 19398
rect -3678 19202 -3672 19370
rect -3638 19330 -3632 19370
rect -2550 19370 -2504 19382
rect -2550 19330 -2544 19370
rect -3638 19202 -2544 19330
rect -2510 19330 -2504 19370
rect -2442 19370 -2396 19382
rect -2360 19380 -1360 19392
rect -2442 19330 -2436 19370
rect -2510 19202 -2436 19330
rect -2402 19330 -2396 19370
rect -1314 19370 -1268 19382
rect -1314 19330 -1308 19370
rect -2402 19320 -1308 19330
rect -2402 19250 -1720 19320
rect -1650 19250 -1500 19320
rect -1430 19250 -1308 19320
rect -2402 19202 -1308 19250
rect -1274 19330 -1268 19370
rect -1206 19370 -1160 19382
rect -1120 19380 -120 19392
rect -1206 19330 -1200 19370
rect -1274 19202 -1200 19330
rect -1166 19330 -1160 19370
rect -78 19370 -32 19382
rect -78 19330 -72 19370
rect -1166 19202 -72 19330
rect -38 19330 -32 19370
rect 30 19370 76 19382
rect 120 19380 1120 19392
rect 1340 19398 1365 19420
rect 2341 19420 2601 19432
rect 2341 19398 2360 19420
rect 30 19330 36 19370
rect -38 19202 36 19330
rect 70 19330 76 19370
rect 1158 19370 1204 19382
rect 1158 19330 1164 19370
rect 70 19202 1164 19330
rect 1198 19330 1204 19370
rect 1266 19370 1312 19382
rect 1340 19380 2360 19398
rect 2580 19398 2601 19420
rect 3577 19398 3600 19432
rect 1266 19330 1272 19370
rect 1198 19202 1272 19330
rect 1306 19330 1312 19370
rect 2394 19370 2440 19382
rect 2394 19330 2400 19370
rect 1306 19320 2400 19330
rect 1306 19250 1460 19320
rect 1530 19250 1700 19320
rect 1770 19250 2400 19320
rect 1306 19202 2400 19250
rect 2434 19330 2440 19370
rect 2502 19370 2548 19382
rect 2580 19380 3600 19398
rect 2502 19330 2508 19370
rect 2434 19202 2508 19330
rect 2542 19330 2548 19370
rect 3630 19370 3676 19382
rect 3630 19330 3636 19370
rect 2542 19202 3636 19330
rect 3670 19202 3676 19370
rect -3678 19190 3676 19202
rect -3678 19174 3670 19190
rect -3678 19140 -3579 19174
rect -2603 19140 -2343 19174
rect -1367 19140 -1107 19174
rect -131 19140 129 19174
rect 1105 19140 1365 19174
rect 2341 19140 2601 19174
rect 3577 19140 3670 19174
rect -3678 19118 3670 19140
rect -3232 19060 -3048 19066
rect -2172 19060 -1988 19066
rect -712 19060 -528 19066
rect 508 19060 692 19066
rect 1988 19060 2172 19066
rect 2988 19060 3172 19066
rect -3600 18900 -3220 19060
rect -3060 18900 -2160 19060
rect -2000 18900 -700 19060
rect -540 18900 520 19060
rect 680 18900 2000 19060
rect 2160 18900 3000 19060
rect 3160 18900 3600 19060
rect -3600 18842 3600 18900
rect -3600 18820 -3579 18842
rect -3591 18808 -3579 18820
rect -2603 18830 -2343 18842
rect -2603 18808 -2591 18830
rect -3591 18802 -2591 18808
rect -2355 18808 -2343 18830
rect -1367 18830 -1107 18842
rect -1367 18808 -1355 18830
rect -2355 18802 -1355 18808
rect -1119 18808 -1107 18830
rect -131 18830 129 18842
rect -131 18808 -119 18830
rect -1119 18802 -119 18808
rect 117 18808 129 18830
rect 1105 18830 1365 18842
rect 1105 18808 1117 18830
rect 117 18802 1117 18808
rect 1353 18808 1365 18830
rect 2341 18830 2601 18842
rect 2341 18808 2353 18830
rect 1353 18802 2353 18808
rect 2589 18808 2601 18830
rect 3577 18820 3600 18842
rect 3577 18808 3589 18820
rect 2589 18802 3589 18808
rect -3678 18780 -3632 18792
rect -3678 18740 -3672 18780
rect -3680 18650 -3672 18740
rect -3678 18612 -3672 18650
rect -3638 18740 -3632 18780
rect -2550 18780 -2504 18792
rect -2550 18740 -2544 18780
rect -3638 18650 -2544 18740
rect -3638 18612 -3632 18650
rect -3678 18600 -3632 18612
rect -2550 18612 -2544 18650
rect -2510 18740 -2504 18780
rect -2442 18780 -2396 18792
rect -2442 18740 -2436 18780
rect -2510 18650 -2436 18740
rect -2510 18612 -2504 18650
rect -2550 18600 -2504 18612
rect -2442 18612 -2436 18650
rect -2402 18740 -2396 18780
rect -1314 18780 -1268 18792
rect -1314 18740 -1308 18780
rect -2402 18730 -1308 18740
rect -2402 18660 -1720 18730
rect -1650 18660 -1500 18730
rect -1430 18660 -1308 18730
rect -2402 18650 -1308 18660
rect -2402 18612 -2396 18650
rect -2442 18600 -2396 18612
rect -1314 18612 -1308 18650
rect -1274 18740 -1268 18780
rect -1206 18780 -1160 18792
rect -1206 18740 -1200 18780
rect -1274 18650 -1200 18740
rect -1274 18612 -1268 18650
rect -1314 18600 -1268 18612
rect -1206 18612 -1200 18650
rect -1166 18740 -1160 18780
rect -78 18780 -32 18792
rect -78 18740 -72 18780
rect -1166 18650 -72 18740
rect -1166 18612 -1160 18650
rect -1206 18600 -1160 18612
rect -78 18612 -72 18650
rect -38 18740 -32 18780
rect 30 18780 76 18792
rect 30 18740 36 18780
rect -38 18650 36 18740
rect -38 18612 -32 18650
rect -78 18600 -32 18612
rect 30 18612 36 18650
rect 70 18740 76 18780
rect 1158 18780 1204 18792
rect 1158 18740 1164 18780
rect 70 18650 1164 18740
rect 70 18612 76 18650
rect 30 18600 76 18612
rect 1158 18612 1164 18650
rect 1198 18740 1204 18780
rect 1266 18780 1312 18792
rect 1266 18740 1272 18780
rect 1198 18650 1272 18740
rect 1198 18612 1204 18650
rect 1158 18600 1204 18612
rect 1266 18612 1272 18650
rect 1306 18740 1312 18780
rect 2394 18780 2440 18792
rect 2394 18740 2400 18780
rect 1306 18730 2400 18740
rect 1306 18660 1460 18730
rect 1530 18660 1700 18730
rect 1770 18660 2400 18730
rect 1306 18650 2400 18660
rect 1306 18612 1312 18650
rect 1266 18600 1312 18612
rect 2394 18612 2400 18650
rect 2434 18740 2440 18780
rect 2502 18780 2548 18792
rect 2502 18740 2508 18780
rect 2434 18650 2508 18740
rect 2434 18612 2440 18650
rect 2394 18600 2440 18612
rect 2502 18612 2508 18650
rect 2542 18740 2548 18780
rect 3630 18780 3676 18792
rect 3630 18740 3636 18780
rect 2542 18650 3636 18740
rect 2542 18612 2548 18650
rect 2502 18600 2548 18612
rect 3630 18612 3636 18650
rect 3670 18612 3676 18780
rect 3630 18600 3676 18612
rect -3600 18584 -2591 18590
rect -3600 18550 -3579 18584
rect -2603 18570 -2591 18584
rect -2355 18584 -1355 18590
rect -2355 18570 -2343 18584
rect -2603 18550 -2343 18570
rect -1367 18570 -1355 18584
rect -1119 18584 -119 18590
rect -1119 18570 -1107 18584
rect -131 18570 -119 18584
rect 117 18584 1117 18590
rect 117 18570 129 18584
rect 1105 18570 1117 18584
rect 1353 18584 2353 18590
rect 1353 18570 1365 18584
rect -1367 18550 -1107 18570
rect -131 18550 129 18570
rect 1105 18550 1365 18570
rect 2341 18570 2353 18584
rect 2589 18584 3594 18590
rect 2589 18570 2601 18584
rect 2341 18550 2601 18570
rect 3577 18550 3594 18584
rect -3600 18500 -560 18550
rect -490 18500 -450 18550
rect -380 18500 380 18550
rect 450 18500 490 18550
rect 560 18500 3594 18550
rect -3600 18490 3594 18500
rect -920 18052 900 18080
rect -920 18018 -818 18052
rect -592 18018 -350 18052
rect -124 18018 118 18052
rect 344 18018 586 18052
rect 812 18018 900 18052
rect -920 18010 900 18018
rect -920 18000 380 18010
rect -920 17990 -560 18000
rect -920 17930 -902 17990
rect -908 17822 -902 17930
rect -868 17930 -560 17990
rect -490 17930 -450 18000
rect -380 17990 380 18000
rect -380 17930 -74 17990
rect -868 17850 -542 17930
rect -868 17822 -862 17850
rect -908 17810 -862 17822
rect -550 17822 -542 17850
rect -508 17822 -434 17930
rect -400 17850 -74 17930
rect -400 17822 -390 17850
rect -550 17810 -390 17822
rect -80 17822 -74 17850
rect -40 17822 34 17990
rect 68 17940 380 17990
rect 450 17940 490 18010
rect 560 18002 900 18010
rect 560 17990 902 18002
rect 560 17940 862 17990
rect 68 17850 394 17940
rect 68 17822 75 17850
rect -80 17810 75 17822
rect 388 17822 394 17850
rect 428 17822 502 17940
rect 536 17850 862 17940
rect 536 17822 545 17850
rect 388 17810 545 17822
rect 856 17822 862 17850
rect 896 17822 902 17990
rect 856 17810 902 17822
rect -830 17794 -580 17800
rect -830 17780 -818 17794
rect -840 17760 -818 17780
rect -592 17780 -580 17794
rect -362 17794 -112 17800
rect -362 17780 -350 17794
rect -592 17760 -350 17780
rect -124 17780 -112 17794
rect 106 17794 356 17800
rect 106 17780 118 17794
rect -124 17760 118 17780
rect 344 17780 356 17794
rect 574 17794 824 17800
rect 574 17780 586 17794
rect 344 17760 586 17780
rect 812 17780 824 17794
rect 812 17760 830 17780
rect -840 17740 830 17760
rect -840 17686 870 17740
rect -852 17680 882 17686
rect -852 17530 -840 17680
rect -620 17670 -320 17680
rect -620 17530 -608 17670
rect -852 17524 -608 17530
rect -332 17530 -320 17670
rect -100 17670 100 17680
rect -100 17530 -88 17670
rect -332 17524 -88 17530
rect 88 17530 100 17670
rect 320 17670 650 17680
rect 320 17530 332 17670
rect 88 17524 332 17530
rect 638 17530 650 17670
rect 870 17530 882 17680
rect 638 17524 882 17530
rect 1440 17490 1790 17510
rect -1740 17470 1460 17490
rect -1740 17400 -1720 17470
rect -1650 17400 -1510 17470
rect -1440 17427 1460 17470
rect -1440 17400 -598 17427
rect -1740 17393 -598 17400
rect -122 17393 120 17427
rect 596 17420 1460 17427
rect 1530 17420 1700 17490
rect 1770 17420 1790 17490
rect 596 17400 1790 17420
rect 596 17393 1460 17400
rect -1740 17380 1460 17393
rect -1740 17310 -1720 17380
rect -1650 17310 -1510 17380
rect -1440 17365 1460 17380
rect -1440 17310 -682 17365
rect -1740 17280 -1410 17310
rect -688 17297 -682 17310
rect -648 17310 -72 17365
rect -648 17297 -642 17310
rect -688 17285 -642 17297
rect -78 17297 -72 17310
rect -38 17310 36 17365
rect -38 17297 -32 17310
rect -78 17285 -32 17297
rect 30 17297 36 17310
rect 70 17310 646 17365
rect 70 17297 76 17310
rect 30 17285 76 17297
rect 640 17297 646 17310
rect 680 17330 1460 17365
rect 1530 17330 1700 17400
rect 1770 17330 1790 17400
rect 680 17310 1790 17330
rect 680 17297 686 17310
rect 640 17285 686 17297
rect -610 17269 -110 17275
rect -610 17255 -598 17269
rect -615 17240 -598 17255
rect -122 17255 -110 17269
rect 108 17269 608 17275
rect 108 17255 120 17269
rect -620 17235 -598 17240
rect -122 17235 120 17255
rect 596 17255 608 17269
rect 596 17240 620 17255
rect 596 17235 630 17240
rect -620 17180 -560 17235
rect -490 17180 -450 17235
rect -380 17180 380 17235
rect 450 17180 490 17235
rect 560 17180 630 17235
rect -620 17170 630 17180
rect -1092 17130 -888 17136
rect -3212 17120 -3008 17126
rect -3212 16990 -3200 17120
rect -3020 16990 -3008 17120
rect -3212 16984 -3008 16990
rect -2072 17120 -1868 17126
rect -2072 16990 -2060 17120
rect -1880 16990 -1868 17120
rect -1092 17000 -1080 17130
rect -900 17000 -888 17130
rect -1092 16994 -888 17000
rect -322 17130 -118 17136
rect -322 17000 -310 17130
rect -130 17000 -118 17130
rect -322 16994 -118 17000
rect 118 17130 322 17136
rect 118 17000 130 17130
rect 310 17000 322 17130
rect 1908 17130 2112 17136
rect 118 16994 322 17000
rect 838 17120 1042 17126
rect -2072 16984 -1868 16990
rect 838 16990 850 17120
rect 1030 16990 1042 17120
rect 1908 17000 1920 17130
rect 2100 17000 2112 17130
rect 1908 16994 2112 17000
rect 2908 17130 3112 17136
rect 2908 17000 2920 17130
rect 3100 17000 3112 17130
rect 2908 16994 3112 17000
rect 838 16984 1042 16990
rect -3550 16950 3540 16955
rect -3550 16902 -1720 16950
rect -1650 16902 -1500 16950
rect -1430 16902 1460 16950
rect 1530 16902 1700 16950
rect 1770 16908 3540 16950
rect 1770 16902 3545 16908
rect -3550 16880 -3533 16902
rect -3545 16868 -3533 16880
rect -2557 16880 -2315 16902
rect -1339 16880 -1097 16902
rect -2557 16868 -2545 16880
rect -3545 16862 -2545 16868
rect -2327 16868 -2315 16880
rect -1339 16868 -1327 16880
rect -2327 16862 -1327 16868
rect -1109 16868 -1097 16880
rect -121 16880 121 16902
rect -121 16868 -109 16880
rect -1109 16862 -109 16868
rect 109 16868 121 16880
rect 1097 16880 1339 16902
rect 2315 16880 2557 16902
rect 1097 16868 1109 16880
rect 109 16862 1109 16868
rect 1327 16868 1339 16880
rect 2315 16868 2327 16880
rect 1327 16862 2327 16868
rect 2545 16868 2557 16880
rect 3533 16868 3545 16902
rect 2545 16862 3545 16868
rect -3623 16840 -3577 16852
rect -3623 16672 -3617 16840
rect -3583 16805 -3577 16840
rect -2513 16840 -2467 16852
rect -2513 16805 -2507 16840
rect -3583 16720 -2507 16805
rect -3583 16672 -3577 16720
rect -3623 16660 -3577 16672
rect -2513 16672 -2507 16720
rect -2473 16805 -2467 16840
rect -2405 16840 -2359 16852
rect -2405 16805 -2399 16840
rect -2473 16720 -2399 16805
rect -2473 16672 -2467 16720
rect -2513 16660 -2467 16672
rect -2405 16672 -2399 16720
rect -2365 16805 -2359 16840
rect -1295 16840 -1249 16852
rect -1295 16805 -1289 16840
rect -2365 16720 -1289 16805
rect -2365 16672 -2359 16720
rect -2405 16660 -2359 16672
rect -1295 16672 -1289 16720
rect -1255 16805 -1249 16840
rect -1187 16840 -1141 16852
rect -1187 16805 -1181 16840
rect -1255 16720 -1181 16805
rect -1255 16672 -1249 16720
rect -1295 16660 -1249 16672
rect -1187 16672 -1181 16720
rect -1147 16805 -1141 16840
rect -77 16840 -31 16852
rect -77 16805 -71 16840
rect -1147 16800 -71 16805
rect -1147 16730 -560 16800
rect -490 16730 -450 16800
rect -380 16730 -71 16800
rect -1147 16720 -71 16730
rect -1147 16672 -1141 16720
rect -1187 16660 -1141 16672
rect -77 16672 -71 16720
rect -37 16805 -31 16840
rect 31 16840 77 16852
rect 31 16805 37 16840
rect -37 16720 37 16805
rect -37 16672 -31 16720
rect -77 16660 -31 16672
rect 31 16672 37 16720
rect 71 16805 77 16840
rect 1141 16840 1187 16852
rect 1141 16805 1147 16840
rect 71 16800 1147 16805
rect 71 16730 380 16800
rect 450 16730 490 16800
rect 560 16730 1147 16800
rect 71 16720 1147 16730
rect 71 16672 77 16720
rect 31 16660 77 16672
rect 1141 16672 1147 16720
rect 1181 16805 1187 16840
rect 1249 16840 1295 16852
rect 1249 16805 1255 16840
rect 1181 16720 1255 16805
rect 1181 16672 1187 16720
rect 1141 16660 1187 16672
rect 1249 16672 1255 16720
rect 1289 16805 1295 16840
rect 2359 16840 2405 16852
rect 2359 16805 2365 16840
rect 1289 16720 2365 16805
rect 1289 16672 1295 16720
rect 1249 16660 1295 16672
rect 2359 16672 2365 16720
rect 2399 16805 2405 16840
rect 2467 16840 2513 16852
rect 2467 16805 2473 16840
rect 2399 16720 2473 16805
rect 2399 16672 2405 16720
rect 2359 16660 2405 16672
rect 2467 16672 2473 16720
rect 2507 16805 2513 16840
rect 3577 16840 3623 16852
rect 3577 16805 3583 16840
rect 2507 16720 3583 16805
rect 2507 16672 2513 16720
rect 2467 16660 2513 16672
rect 3577 16672 3583 16720
rect 3617 16672 3623 16840
rect 3577 16660 3623 16672
rect -3545 16644 -2545 16650
rect -3545 16630 -3533 16644
rect -3550 16610 -3533 16630
rect -2557 16630 -2545 16644
rect -2327 16644 -1327 16650
rect -2327 16630 -2315 16644
rect -2557 16610 -2315 16630
rect -1339 16630 -1327 16644
rect -1109 16644 -109 16650
rect -1109 16630 -1097 16644
rect -1339 16610 -1097 16630
rect -121 16630 -109 16644
rect 109 16644 1109 16650
rect 109 16630 121 16644
rect -121 16610 121 16630
rect 1097 16630 1109 16644
rect 1327 16644 2327 16650
rect 1327 16630 1339 16644
rect 1097 16610 1339 16630
rect 2315 16630 2327 16644
rect 2545 16644 3545 16650
rect 2545 16630 2557 16644
rect 2315 16610 2557 16630
rect 3533 16610 3545 16644
rect -3550 16604 3545 16610
rect -3550 16555 3540 16604
rect -2200 16260 -1800 16555
rect -800 16260 -400 16555
rect 500 16260 900 16555
rect 1790 16260 2200 16555
rect -3000 16152 3000 16260
rect -3000 16146 203 16152
rect -3000 15749 -2827 16146
rect -1713 15749 -1307 16146
rect -193 15755 203 16146
rect 1317 15755 1713 16152
rect 2827 15755 3000 16152
rect -193 15749 3000 15755
rect -3000 15660 3000 15749
rect -3252 15220 -3108 15226
rect -3252 15100 -3240 15220
rect -3120 15100 -3108 15220
rect -3252 15094 -3108 15100
rect 3118 15220 3262 15226
rect 3118 15100 3130 15220
rect 3250 15100 3262 15220
rect 3118 15094 3262 15100
rect -3252 12220 -3108 12226
rect -3252 12100 -3240 12220
rect -3120 12100 -3108 12220
rect -3252 12094 -3108 12100
rect 3118 12220 3262 12226
rect 3118 12100 3130 12220
rect 3250 12100 3262 12220
rect 3118 12094 3262 12100
rect -3252 9220 -3108 9226
rect -3252 9100 -3240 9220
rect -3120 9100 -3108 9220
rect -3252 9094 -3108 9100
rect 3118 9220 3262 9226
rect 3118 9100 3130 9220
rect 3250 9100 3262 9220
rect 3118 9094 3262 9100
rect -3252 6220 -3108 6226
rect -3252 6100 -3240 6220
rect -3120 6100 -3108 6220
rect -3252 6094 -3108 6100
rect 3118 6220 3262 6226
rect 3118 6100 3130 6220
rect 3250 6100 3262 6220
rect 3118 6094 3262 6100
rect -3252 3220 -3108 3226
rect -3252 3100 -3240 3220
rect -3120 3100 -3108 3220
rect -3252 3094 -3108 3100
rect 3118 3220 3262 3226
rect 3118 3100 3130 3220
rect 3250 3100 3262 3220
rect 3118 3094 3262 3100
rect -3000 1921 3000 1960
rect -3000 1915 203 1921
rect -3000 1890 -2827 1915
rect -1713 1890 -1307 1915
rect -193 1890 203 1915
rect 1317 1900 1713 1921
rect 2827 1900 3000 1921
rect 1317 1890 1690 1900
rect -3000 1480 -2860 1890
rect -1690 1480 -1350 1890
rect -180 1480 170 1890
rect 1340 1490 1690 1890
rect 2860 1490 3000 1900
rect 1340 1480 3000 1490
rect -3000 1460 3000 1480
<< via1 >>
rect -7912 30560 -7852 30620
rect -7792 30560 -7732 30620
rect -629 31143 -385 31387
rect 421 31143 665 31387
rect -3183 30910 -3172 30911
rect -3172 30910 -3138 30911
rect -3138 30910 -3131 30911
rect -3183 30872 -3131 30910
rect -3183 30859 -3172 30872
rect -3172 30859 -3138 30872
rect -3138 30859 -3131 30872
rect -2863 30910 -2856 30911
rect -2856 30910 -2822 30911
rect -2822 30910 -2811 30911
rect -2863 30872 -2811 30910
rect -2863 30859 -2856 30872
rect -2856 30859 -2822 30872
rect -2822 30859 -2811 30872
rect -3183 30656 -3131 30671
rect -3183 30622 -3172 30656
rect -3172 30622 -3138 30656
rect -3138 30622 -3131 30656
rect -3183 30619 -3131 30622
rect -2553 30910 -2540 30911
rect -2540 30910 -2506 30911
rect -2506 30910 -2501 30911
rect -2553 30872 -2501 30910
rect -2553 30859 -2540 30872
rect -2540 30859 -2506 30872
rect -2506 30859 -2501 30872
rect -2863 30656 -2811 30671
rect -2863 30622 -2856 30656
rect -2856 30622 -2822 30656
rect -2822 30622 -2811 30656
rect -2863 30619 -2811 30622
rect -2233 30910 -2224 30911
rect -2224 30910 -2190 30911
rect -2190 30910 -2181 30911
rect -2233 30872 -2181 30910
rect -2233 30859 -2224 30872
rect -2224 30859 -2190 30872
rect -2190 30859 -2181 30872
rect -3023 30296 -2971 30301
rect -3023 30262 -3014 30296
rect -3014 30262 -2980 30296
rect -2980 30262 -2971 30296
rect -3023 30249 -2971 30262
rect -2553 30656 -2501 30671
rect -2553 30622 -2540 30656
rect -2540 30622 -2506 30656
rect -2506 30622 -2501 30656
rect -2553 30619 -2501 30622
rect -1923 30910 -1908 30911
rect -1908 30910 -1874 30911
rect -1874 30910 -1871 30911
rect -1923 30872 -1871 30910
rect -1923 30859 -1908 30872
rect -1908 30859 -1874 30872
rect -1874 30859 -1871 30872
rect -2713 30296 -2661 30301
rect -2713 30262 -2698 30296
rect -2698 30262 -2664 30296
rect -2664 30262 -2661 30296
rect -2713 30249 -2661 30262
rect -2233 30656 -2181 30671
rect -2233 30622 -2224 30656
rect -2224 30622 -2190 30656
rect -2190 30622 -2181 30656
rect -2233 30619 -2181 30622
rect -1603 30910 -1592 30911
rect -1592 30910 -1558 30911
rect -1558 30910 -1551 30911
rect -1603 30872 -1551 30910
rect -1603 30859 -1592 30872
rect -1592 30859 -1558 30872
rect -1558 30859 -1551 30872
rect -3023 30046 -3014 30061
rect -3014 30046 -2980 30061
rect -2980 30046 -2971 30061
rect -3023 30009 -2971 30046
rect -2393 30296 -2341 30301
rect -2393 30262 -2382 30296
rect -2382 30262 -2348 30296
rect -2348 30262 -2341 30296
rect -2393 30249 -2341 30262
rect -1923 30656 -1871 30671
rect -1923 30622 -1908 30656
rect -1908 30622 -1874 30656
rect -1874 30622 -1871 30656
rect -1923 30619 -1871 30622
rect -1283 30910 -1276 30911
rect -1276 30910 -1242 30911
rect -1242 30910 -1231 30911
rect -1283 30872 -1231 30910
rect -1283 30859 -1276 30872
rect -1276 30859 -1242 30872
rect -1242 30859 -1231 30872
rect -2713 30046 -2698 30061
rect -2698 30046 -2664 30061
rect -2664 30046 -2661 30061
rect -2713 30009 -2661 30046
rect -2073 30296 -2021 30301
rect -2073 30262 -2066 30296
rect -2066 30262 -2032 30296
rect -2032 30262 -2021 30296
rect -2073 30249 -2021 30262
rect -1603 30656 -1551 30671
rect -1603 30622 -1592 30656
rect -1592 30622 -1558 30656
rect -1558 30622 -1551 30656
rect -1603 30619 -1551 30622
rect -973 30910 -960 30911
rect -960 30910 -926 30911
rect -926 30910 -921 30911
rect -973 30872 -921 30910
rect -973 30859 -960 30872
rect -960 30859 -926 30872
rect -926 30859 -921 30872
rect -2393 30046 -2382 30061
rect -2382 30046 -2348 30061
rect -2348 30046 -2341 30061
rect -2393 30009 -2341 30046
rect -1763 30296 -1711 30301
rect -1763 30262 -1750 30296
rect -1750 30262 -1716 30296
rect -1716 30262 -1711 30296
rect -1763 30249 -1711 30262
rect -1283 30656 -1231 30671
rect -1283 30622 -1276 30656
rect -1276 30622 -1242 30656
rect -1242 30622 -1231 30656
rect -1283 30619 -1231 30622
rect -653 30910 -644 30911
rect -644 30910 -610 30911
rect -610 30910 -601 30911
rect -653 30872 -601 30910
rect -653 30859 -644 30872
rect -644 30859 -610 30872
rect -610 30859 -601 30872
rect -2073 30046 -2066 30061
rect -2066 30046 -2032 30061
rect -2032 30046 -2021 30061
rect -2073 30009 -2021 30046
rect -1443 30296 -1391 30301
rect -1443 30262 -1434 30296
rect -1434 30262 -1400 30296
rect -1400 30262 -1391 30296
rect -1443 30249 -1391 30262
rect -973 30656 -921 30671
rect -973 30622 -960 30656
rect -960 30622 -926 30656
rect -926 30622 -921 30656
rect -973 30619 -921 30622
rect -333 30910 -328 30911
rect -328 30910 -294 30911
rect -294 30910 -281 30911
rect -333 30872 -281 30910
rect -333 30859 -328 30872
rect -328 30859 -294 30872
rect -294 30859 -281 30872
rect -1763 30046 -1750 30061
rect -1750 30046 -1716 30061
rect -1716 30046 -1711 30061
rect -1763 30009 -1711 30046
rect -1133 30296 -1081 30301
rect -1133 30262 -1118 30296
rect -1118 30262 -1084 30296
rect -1084 30262 -1081 30296
rect -1133 30249 -1081 30262
rect -653 30656 -601 30671
rect -653 30622 -644 30656
rect -644 30622 -610 30656
rect -610 30622 -601 30656
rect -653 30619 -601 30622
rect -23 30910 -12 30911
rect -12 30910 22 30911
rect 22 30910 29 30911
rect -23 30872 29 30910
rect -23 30859 -12 30872
rect -12 30859 22 30872
rect 22 30859 29 30872
rect -1443 30046 -1434 30061
rect -1434 30046 -1400 30061
rect -1400 30046 -1391 30061
rect -1443 30009 -1391 30046
rect -813 30296 -761 30301
rect -813 30262 -802 30296
rect -802 30262 -768 30296
rect -768 30262 -761 30296
rect -813 30249 -761 30262
rect -333 30656 -281 30671
rect -333 30622 -328 30656
rect -328 30622 -294 30656
rect -294 30622 -281 30656
rect -333 30619 -281 30622
rect 297 30910 304 30911
rect 304 30910 338 30911
rect 338 30910 349 30911
rect 297 30872 349 30910
rect 297 30859 304 30872
rect 304 30859 338 30872
rect 338 30859 349 30872
rect -1133 30046 -1118 30061
rect -1118 30046 -1084 30061
rect -1084 30046 -1081 30061
rect -1133 30009 -1081 30046
rect -493 30296 -441 30301
rect -493 30262 -486 30296
rect -486 30262 -452 30296
rect -452 30262 -441 30296
rect -493 30249 -441 30262
rect -23 30656 29 30671
rect -23 30622 -12 30656
rect -12 30622 22 30656
rect 22 30622 29 30656
rect -23 30619 29 30622
rect 607 30910 620 30911
rect 620 30910 654 30911
rect 654 30910 659 30911
rect 607 30872 659 30910
rect 607 30859 620 30872
rect 620 30859 654 30872
rect 654 30859 659 30872
rect -813 30046 -802 30061
rect -802 30046 -768 30061
rect -768 30046 -761 30061
rect -813 30009 -761 30046
rect -183 30296 -131 30301
rect -183 30262 -170 30296
rect -170 30262 -136 30296
rect -136 30262 -131 30296
rect -183 30249 -131 30262
rect 297 30656 349 30671
rect 297 30622 304 30656
rect 304 30622 338 30656
rect 338 30622 349 30656
rect 297 30619 349 30622
rect 927 30910 936 30911
rect 936 30910 970 30911
rect 970 30910 979 30911
rect 927 30872 979 30910
rect 927 30859 936 30872
rect 936 30859 970 30872
rect 970 30859 979 30872
rect -493 30046 -486 30061
rect -486 30046 -452 30061
rect -452 30046 -441 30061
rect -493 30009 -441 30046
rect 137 30296 189 30301
rect 137 30262 146 30296
rect 146 30262 180 30296
rect 180 30262 189 30296
rect 137 30249 189 30262
rect 607 30656 659 30671
rect 607 30622 620 30656
rect 620 30622 654 30656
rect 654 30622 659 30656
rect 607 30619 659 30622
rect 1247 30910 1252 30911
rect 1252 30910 1286 30911
rect 1286 30910 1299 30911
rect 1247 30872 1299 30910
rect 1247 30859 1252 30872
rect 1252 30859 1286 30872
rect 1286 30859 1299 30872
rect -183 30046 -170 30061
rect -170 30046 -136 30061
rect -136 30046 -131 30061
rect -183 30009 -131 30046
rect 457 30296 509 30301
rect 457 30262 462 30296
rect 462 30262 496 30296
rect 496 30262 509 30296
rect 457 30249 509 30262
rect 927 30656 979 30671
rect 927 30622 936 30656
rect 936 30622 970 30656
rect 970 30622 979 30656
rect 927 30619 979 30622
rect 1557 30910 1568 30911
rect 1568 30910 1602 30911
rect 1602 30910 1609 30911
rect 1557 30872 1609 30910
rect 1557 30859 1568 30872
rect 1568 30859 1602 30872
rect 1602 30859 1609 30872
rect 137 30046 146 30061
rect 146 30046 180 30061
rect 180 30046 189 30061
rect 137 30009 189 30046
rect 767 30296 819 30301
rect 767 30262 778 30296
rect 778 30262 812 30296
rect 812 30262 819 30296
rect 767 30249 819 30262
rect 1247 30656 1299 30671
rect 1247 30622 1252 30656
rect 1252 30622 1286 30656
rect 1286 30622 1299 30656
rect 1247 30619 1299 30622
rect 1877 30910 1884 30911
rect 1884 30910 1918 30911
rect 1918 30910 1929 30911
rect 1877 30872 1929 30910
rect 1877 30859 1884 30872
rect 1884 30859 1918 30872
rect 1918 30859 1929 30872
rect 457 30046 462 30061
rect 462 30046 496 30061
rect 496 30046 509 30061
rect 457 30009 509 30046
rect 1087 30296 1139 30301
rect 1087 30262 1094 30296
rect 1094 30262 1128 30296
rect 1128 30262 1139 30296
rect 1087 30249 1139 30262
rect 1557 30656 1609 30671
rect 1557 30622 1568 30656
rect 1568 30622 1602 30656
rect 1602 30622 1609 30656
rect 1557 30619 1609 30622
rect 2187 30910 2200 30911
rect 2200 30910 2234 30911
rect 2234 30910 2239 30911
rect 2187 30872 2239 30910
rect 2187 30859 2200 30872
rect 2200 30859 2234 30872
rect 2234 30859 2239 30872
rect 767 30046 778 30061
rect 778 30046 812 30061
rect 812 30046 819 30061
rect 767 30009 819 30046
rect 1397 30296 1449 30301
rect 1397 30262 1410 30296
rect 1410 30262 1444 30296
rect 1444 30262 1449 30296
rect 1397 30249 1449 30262
rect 1877 30656 1929 30671
rect 1877 30622 1884 30656
rect 1884 30622 1918 30656
rect 1918 30622 1929 30656
rect 1877 30619 1929 30622
rect 2507 30910 2516 30911
rect 2516 30910 2550 30911
rect 2550 30910 2559 30911
rect 2507 30872 2559 30910
rect 2507 30859 2516 30872
rect 2516 30859 2550 30872
rect 2550 30859 2559 30872
rect 1087 30046 1094 30061
rect 1094 30046 1128 30061
rect 1128 30046 1139 30061
rect 1087 30009 1139 30046
rect 1717 30296 1769 30301
rect 1717 30262 1726 30296
rect 1726 30262 1760 30296
rect 1760 30262 1769 30296
rect 1717 30249 1769 30262
rect 2187 30656 2239 30671
rect 2187 30622 2200 30656
rect 2200 30622 2234 30656
rect 2234 30622 2239 30656
rect 2187 30619 2239 30622
rect 2827 30910 2832 30911
rect 2832 30910 2866 30911
rect 2866 30910 2879 30911
rect 2827 30872 2879 30910
rect 2827 30859 2832 30872
rect 2832 30859 2866 30872
rect 2866 30859 2879 30872
rect 1397 30046 1410 30061
rect 1410 30046 1444 30061
rect 1444 30046 1449 30061
rect 1397 30009 1449 30046
rect 2037 30296 2089 30301
rect 2037 30262 2042 30296
rect 2042 30262 2076 30296
rect 2076 30262 2089 30296
rect 2037 30249 2089 30262
rect 2507 30656 2559 30671
rect 2507 30622 2516 30656
rect 2516 30622 2550 30656
rect 2550 30622 2559 30656
rect 2507 30619 2559 30622
rect 3137 30910 3148 30911
rect 3148 30910 3182 30911
rect 3182 30910 3189 30911
rect 3137 30872 3189 30910
rect 3137 30859 3148 30872
rect 3148 30859 3182 30872
rect 3182 30859 3189 30872
rect 1717 30046 1726 30061
rect 1726 30046 1760 30061
rect 1760 30046 1769 30061
rect 1717 30009 1769 30046
rect 2347 30296 2399 30301
rect 2347 30262 2358 30296
rect 2358 30262 2392 30296
rect 2392 30262 2399 30296
rect 2347 30249 2399 30262
rect 2827 30656 2879 30671
rect 2827 30622 2832 30656
rect 2832 30622 2866 30656
rect 2866 30622 2879 30656
rect 2827 30619 2879 30622
rect 2037 30046 2042 30061
rect 2042 30046 2076 30061
rect 2076 30046 2089 30061
rect 2037 30009 2089 30046
rect 2667 30296 2719 30301
rect 2667 30262 2674 30296
rect 2674 30262 2708 30296
rect 2708 30262 2719 30296
rect 2667 30249 2719 30262
rect 3137 30656 3189 30671
rect 3137 30622 3148 30656
rect 3148 30622 3182 30656
rect 3182 30622 3189 30656
rect 3137 30619 3189 30622
rect 2347 30046 2358 30061
rect 2358 30046 2392 30061
rect 2392 30046 2399 30061
rect 2347 30009 2399 30046
rect 2987 30296 3039 30301
rect 2987 30262 2990 30296
rect 2990 30262 3024 30296
rect 3024 30262 3039 30296
rect 2987 30249 3039 30262
rect 2667 30046 2674 30061
rect 2674 30046 2708 30061
rect 2708 30046 2719 30061
rect 2667 30009 2719 30046
rect 2987 30046 2990 30061
rect 2990 30046 3024 30061
rect 3024 30046 3039 30061
rect 2987 30009 3039 30046
rect -2058 29834 -2006 29886
rect 2002 29834 2054 29886
rect -629 29503 -385 29747
rect 421 29503 665 29747
rect -1683 29240 -1672 29241
rect -1672 29240 -1638 29241
rect -1638 29240 -1631 29241
rect -1683 29202 -1631 29240
rect -1683 29189 -1672 29202
rect -1672 29189 -1638 29202
rect -1638 29189 -1631 29202
rect -1363 29240 -1356 29241
rect -1356 29240 -1322 29241
rect -1322 29240 -1311 29241
rect -1363 29202 -1311 29240
rect -1363 29189 -1356 29202
rect -1356 29189 -1322 29202
rect -1322 29189 -1311 29202
rect -1683 29024 -1672 29031
rect -1672 29024 -1638 29031
rect -1638 29024 -1631 29031
rect -1683 28986 -1631 29024
rect -1683 28979 -1672 28986
rect -1672 28979 -1638 28986
rect -1638 28979 -1631 28986
rect -1053 29240 -1040 29241
rect -1040 29240 -1006 29241
rect -1006 29240 -1001 29241
rect -1053 29202 -1001 29240
rect -1053 29189 -1040 29202
rect -1040 29189 -1006 29202
rect -1006 29189 -1001 29202
rect -1363 29024 -1356 29031
rect -1356 29024 -1322 29031
rect -1322 29024 -1311 29031
rect -1363 28986 -1311 29024
rect -1363 28979 -1356 28986
rect -1356 28979 -1322 28986
rect -1322 28979 -1311 28986
rect -1523 28592 -1514 28601
rect -1514 28592 -1480 28601
rect -1480 28592 -1471 28601
rect -1523 28554 -1471 28592
rect -1523 28549 -1514 28554
rect -1514 28549 -1480 28554
rect -1480 28549 -1471 28554
rect -733 29240 -724 29241
rect -724 29240 -690 29241
rect -690 29240 -681 29241
rect -733 29202 -681 29240
rect -733 29189 -724 29202
rect -724 29189 -690 29202
rect -690 29189 -681 29202
rect -1053 29024 -1040 29031
rect -1040 29024 -1006 29031
rect -1006 29024 -1001 29031
rect -1053 28986 -1001 29024
rect -1053 28979 -1040 28986
rect -1040 28979 -1006 28986
rect -1006 28979 -1001 28986
rect -1203 28592 -1198 28601
rect -1198 28592 -1164 28601
rect -1164 28592 -1151 28601
rect -1203 28554 -1151 28592
rect -1203 28549 -1198 28554
rect -1198 28549 -1164 28554
rect -1164 28549 -1151 28554
rect -1523 28376 -1514 28391
rect -1514 28376 -1480 28391
rect -1480 28376 -1471 28391
rect -1523 28339 -1471 28376
rect -413 29240 -408 29241
rect -408 29240 -374 29241
rect -374 29240 -361 29241
rect -413 29202 -361 29240
rect -413 29189 -408 29202
rect -408 29189 -374 29202
rect -374 29189 -361 29202
rect -733 29024 -724 29031
rect -724 29024 -690 29031
rect -690 29024 -681 29031
rect -733 28986 -681 29024
rect -733 28979 -724 28986
rect -724 28979 -690 28986
rect -690 28979 -681 28986
rect -893 28592 -882 28601
rect -882 28592 -848 28601
rect -848 28592 -841 28601
rect -893 28554 -841 28592
rect -893 28549 -882 28554
rect -882 28549 -848 28554
rect -848 28549 -841 28554
rect -1203 28376 -1198 28391
rect -1198 28376 -1164 28391
rect -1164 28376 -1151 28391
rect -1203 28339 -1151 28376
rect -103 29240 -92 29241
rect -92 29240 -58 29241
rect -58 29240 -51 29241
rect -103 29202 -51 29240
rect -103 29189 -92 29202
rect -92 29189 -58 29202
rect -58 29189 -51 29202
rect -413 29024 -408 29031
rect -408 29024 -374 29031
rect -374 29024 -361 29031
rect -413 28986 -361 29024
rect -413 28979 -408 28986
rect -408 28979 -374 28986
rect -374 28979 -361 28986
rect -573 28592 -566 28601
rect -566 28592 -532 28601
rect -532 28592 -521 28601
rect -573 28554 -521 28592
rect -573 28549 -566 28554
rect -566 28549 -532 28554
rect -532 28549 -521 28554
rect -893 28376 -882 28391
rect -882 28376 -848 28391
rect -848 28376 -841 28391
rect -893 28339 -841 28376
rect 217 29240 224 29241
rect 224 29240 258 29241
rect 258 29240 269 29241
rect 217 29202 269 29240
rect 217 29189 224 29202
rect 224 29189 258 29202
rect 258 29189 269 29202
rect -103 29024 -92 29031
rect -92 29024 -58 29031
rect -58 29024 -51 29031
rect -103 28986 -51 29024
rect -103 28979 -92 28986
rect -92 28979 -58 28986
rect -58 28979 -51 28986
rect -253 28592 -250 28601
rect -250 28592 -216 28601
rect -216 28592 -201 28601
rect -253 28554 -201 28592
rect -253 28549 -250 28554
rect -250 28549 -216 28554
rect -216 28549 -201 28554
rect -573 28376 -566 28391
rect -566 28376 -532 28391
rect -532 28376 -521 28391
rect -573 28339 -521 28376
rect 537 29240 540 29241
rect 540 29240 574 29241
rect 574 29240 589 29241
rect 537 29202 589 29240
rect 537 29189 540 29202
rect 540 29189 574 29202
rect 574 29189 589 29202
rect 217 29024 224 29031
rect 224 29024 258 29031
rect 258 29024 269 29031
rect 217 28986 269 29024
rect 217 28979 224 28986
rect 224 28979 258 28986
rect 258 28979 269 28986
rect 57 28592 66 28601
rect 66 28592 100 28601
rect 100 28592 109 28601
rect 57 28554 109 28592
rect 57 28549 66 28554
rect 66 28549 100 28554
rect 100 28549 109 28554
rect -253 28376 -250 28391
rect -250 28376 -216 28391
rect -216 28376 -201 28391
rect -253 28339 -201 28376
rect 847 29240 856 29241
rect 856 29240 890 29241
rect 890 29240 899 29241
rect 847 29202 899 29240
rect 847 29189 856 29202
rect 856 29189 890 29202
rect 890 29189 899 29202
rect 537 29024 540 29031
rect 540 29024 574 29031
rect 574 29024 589 29031
rect 537 28986 589 29024
rect 537 28979 540 28986
rect 540 28979 574 28986
rect 574 28979 589 28986
rect 377 28592 382 28601
rect 382 28592 416 28601
rect 416 28592 429 28601
rect 377 28554 429 28592
rect 377 28549 382 28554
rect 382 28549 416 28554
rect 416 28549 429 28554
rect 57 28376 66 28391
rect 66 28376 100 28391
rect 100 28376 109 28391
rect 57 28339 109 28376
rect 1167 29240 1172 29241
rect 1172 29240 1206 29241
rect 1206 29240 1219 29241
rect 1167 29202 1219 29240
rect 1167 29189 1172 29202
rect 1172 29189 1206 29202
rect 1206 29189 1219 29202
rect 847 29024 856 29031
rect 856 29024 890 29031
rect 890 29024 899 29031
rect 847 28986 899 29024
rect 847 28979 856 28986
rect 856 28979 890 28986
rect 890 28979 899 28986
rect 687 28592 698 28601
rect 698 28592 732 28601
rect 732 28592 739 28601
rect 687 28554 739 28592
rect 687 28549 698 28554
rect 698 28549 732 28554
rect 732 28549 739 28554
rect 377 28376 382 28391
rect 382 28376 416 28391
rect 416 28376 429 28391
rect 377 28339 429 28376
rect 1477 29240 1488 29241
rect 1488 29240 1522 29241
rect 1522 29240 1529 29241
rect 1477 29202 1529 29240
rect 1477 29189 1488 29202
rect 1488 29189 1522 29202
rect 1522 29189 1529 29202
rect 1167 29024 1172 29031
rect 1172 29024 1206 29031
rect 1206 29024 1219 29031
rect 1167 28986 1219 29024
rect 1167 28979 1172 28986
rect 1172 28979 1206 28986
rect 1206 28979 1219 28986
rect 1007 28592 1014 28601
rect 1014 28592 1048 28601
rect 1048 28592 1059 28601
rect 1007 28554 1059 28592
rect 1007 28549 1014 28554
rect 1014 28549 1048 28554
rect 1048 28549 1059 28554
rect 687 28376 698 28391
rect 698 28376 732 28391
rect 732 28376 739 28391
rect 687 28339 739 28376
rect 1477 29024 1488 29031
rect 1488 29024 1522 29031
rect 1522 29024 1529 29031
rect 1477 28986 1529 29024
rect 1477 28979 1488 28986
rect 1488 28979 1522 28986
rect 1522 28979 1529 28986
rect 1327 28592 1330 28601
rect 1330 28592 1364 28601
rect 1364 28592 1379 28601
rect 1327 28554 1379 28592
rect 1327 28549 1330 28554
rect 1330 28549 1364 28554
rect 1364 28549 1379 28554
rect 1007 28376 1014 28391
rect 1014 28376 1048 28391
rect 1048 28376 1059 28391
rect 1007 28339 1059 28376
rect 1637 28592 1646 28601
rect 1646 28592 1680 28601
rect 1680 28592 1689 28601
rect 1637 28554 1689 28592
rect 1637 28549 1646 28554
rect 1646 28549 1680 28554
rect 1680 28549 1689 28554
rect 1327 28376 1330 28391
rect 1330 28376 1364 28391
rect 1364 28376 1379 28391
rect 1327 28339 1379 28376
rect 1637 28376 1646 28391
rect 1646 28376 1680 28391
rect 1680 28376 1689 28391
rect 1637 28339 1689 28376
rect 8002 30564 8054 30616
rect 8112 30564 8164 30616
rect -864 28109 -620 28142
rect -864 27931 -620 28109
rect -864 27898 -620 27931
rect 636 28109 880 28142
rect 636 27931 880 28109
rect 636 27898 880 27931
rect -1683 27662 -1631 27691
rect -1683 27639 -1672 27662
rect -1672 27639 -1638 27662
rect -1638 27639 -1631 27662
rect -1363 27662 -1311 27691
rect -1363 27639 -1356 27662
rect -1356 27639 -1322 27662
rect -1322 27639 -1311 27662
rect -1683 27446 -1631 27481
rect -1683 27429 -1672 27446
rect -1672 27429 -1638 27446
rect -1638 27429 -1631 27446
rect -1053 27662 -1001 27691
rect -1053 27639 -1040 27662
rect -1040 27639 -1006 27662
rect -1006 27639 -1001 27662
rect -1363 27446 -1311 27481
rect -1363 27429 -1356 27446
rect -1356 27429 -1322 27446
rect -1322 27429 -1311 27446
rect -1523 27052 -1514 27061
rect -1514 27052 -1480 27061
rect -1480 27052 -1471 27061
rect -1523 27014 -1471 27052
rect -1523 27009 -1514 27014
rect -1514 27009 -1480 27014
rect -1480 27009 -1471 27014
rect -733 27662 -681 27691
rect -733 27639 -724 27662
rect -724 27639 -690 27662
rect -690 27639 -681 27662
rect -1053 27446 -1001 27481
rect -1053 27429 -1040 27446
rect -1040 27429 -1006 27446
rect -1006 27429 -1001 27446
rect -1203 27052 -1198 27061
rect -1198 27052 -1164 27061
rect -1164 27052 -1151 27061
rect -1203 27014 -1151 27052
rect -1203 27009 -1198 27014
rect -1198 27009 -1164 27014
rect -1164 27009 -1151 27014
rect -1523 26836 -1514 26851
rect -1514 26836 -1480 26851
rect -1480 26836 -1471 26851
rect -1523 26799 -1471 26836
rect -413 27662 -361 27691
rect -413 27639 -408 27662
rect -408 27639 -374 27662
rect -374 27639 -361 27662
rect -733 27446 -681 27481
rect -733 27429 -724 27446
rect -724 27429 -690 27446
rect -690 27429 -681 27446
rect -893 27052 -882 27061
rect -882 27052 -848 27061
rect -848 27052 -841 27061
rect -893 27014 -841 27052
rect -893 27009 -882 27014
rect -882 27009 -848 27014
rect -848 27009 -841 27014
rect -1203 26836 -1198 26851
rect -1198 26836 -1164 26851
rect -1164 26836 -1151 26851
rect -1203 26799 -1151 26836
rect -103 27662 -51 27691
rect -103 27639 -92 27662
rect -92 27639 -58 27662
rect -58 27639 -51 27662
rect -413 27446 -361 27481
rect -413 27429 -408 27446
rect -408 27429 -374 27446
rect -374 27429 -361 27446
rect -573 27052 -566 27061
rect -566 27052 -532 27061
rect -532 27052 -521 27061
rect -573 27014 -521 27052
rect -573 27009 -566 27014
rect -566 27009 -532 27014
rect -532 27009 -521 27014
rect -893 26836 -882 26851
rect -882 26836 -848 26851
rect -848 26836 -841 26851
rect -893 26799 -841 26836
rect 217 27662 269 27691
rect 217 27639 224 27662
rect 224 27639 258 27662
rect 258 27639 269 27662
rect -103 27446 -51 27481
rect -103 27429 -92 27446
rect -92 27429 -58 27446
rect -58 27429 -51 27446
rect -263 27052 -250 27061
rect -250 27052 -216 27061
rect -216 27052 -211 27061
rect -263 27014 -211 27052
rect -263 27009 -250 27014
rect -250 27009 -216 27014
rect -216 27009 -211 27014
rect -573 26836 -566 26851
rect -566 26836 -532 26851
rect -532 26836 -521 26851
rect -573 26799 -521 26836
rect 527 27662 579 27691
rect 527 27639 540 27662
rect 540 27639 574 27662
rect 574 27639 579 27662
rect 217 27446 269 27481
rect 217 27429 224 27446
rect 224 27429 258 27446
rect 258 27429 269 27446
rect 57 27052 66 27061
rect 66 27052 100 27061
rect 100 27052 109 27061
rect 57 27014 109 27052
rect 57 27009 66 27014
rect 66 27009 100 27014
rect 100 27009 109 27014
rect -263 26836 -250 26851
rect -250 26836 -216 26851
rect -216 26836 -211 26851
rect -263 26799 -211 26836
rect 847 27662 899 27691
rect 847 27639 856 27662
rect 856 27639 890 27662
rect 890 27639 899 27662
rect 527 27446 579 27481
rect 527 27429 540 27446
rect 540 27429 574 27446
rect 574 27429 579 27446
rect 377 27052 382 27061
rect 382 27052 416 27061
rect 416 27052 429 27061
rect 377 27014 429 27052
rect 377 27009 382 27014
rect 382 27009 416 27014
rect 416 27009 429 27014
rect 57 26836 66 26851
rect 66 26836 100 26851
rect 100 26836 109 26851
rect 57 26799 109 26836
rect 1167 27662 1219 27691
rect 1167 27639 1172 27662
rect 1172 27639 1206 27662
rect 1206 27639 1219 27662
rect 847 27446 899 27481
rect 847 27429 856 27446
rect 856 27429 890 27446
rect 890 27429 899 27446
rect 687 27052 698 27061
rect 698 27052 732 27061
rect 732 27052 739 27061
rect 687 27014 739 27052
rect 687 27009 698 27014
rect 698 27009 732 27014
rect 732 27009 739 27014
rect 377 26836 382 26851
rect 382 26836 416 26851
rect 416 26836 429 26851
rect 377 26799 429 26836
rect 1477 27662 1529 27691
rect 1477 27639 1488 27662
rect 1488 27639 1522 27662
rect 1522 27639 1529 27662
rect 1167 27446 1219 27481
rect 1167 27429 1172 27446
rect 1172 27429 1206 27446
rect 1206 27429 1219 27446
rect 1007 27052 1014 27061
rect 1014 27052 1048 27061
rect 1048 27052 1059 27061
rect 1007 27014 1059 27052
rect 1007 27009 1014 27014
rect 1014 27009 1048 27014
rect 1048 27009 1059 27014
rect 687 26836 698 26851
rect 698 26836 732 26851
rect 732 26836 739 26851
rect 687 26799 739 26836
rect 1477 27446 1529 27481
rect 1477 27429 1488 27446
rect 1488 27429 1522 27446
rect 1522 27429 1529 27446
rect 1317 27052 1330 27061
rect 1330 27052 1364 27061
rect 1364 27052 1369 27061
rect 1317 27014 1369 27052
rect 1317 27009 1330 27014
rect 1330 27009 1364 27014
rect 1364 27009 1369 27014
rect 1007 26836 1014 26851
rect 1014 26836 1048 26851
rect 1048 26836 1059 26851
rect 1007 26799 1059 26836
rect 1637 27052 1646 27061
rect 1646 27052 1680 27061
rect 1680 27052 1689 27061
rect 1637 27014 1689 27052
rect 1637 27009 1646 27014
rect 1646 27009 1680 27014
rect 1680 27009 1689 27014
rect 1317 26836 1330 26851
rect 1330 26836 1364 26851
rect 1364 26836 1369 26851
rect 1317 26799 1369 26836
rect 1637 26836 1646 26851
rect 1646 26836 1680 26851
rect 1680 26836 1689 26851
rect 1637 26799 1689 26836
rect -583 26094 -531 26131
rect -583 26079 -571 26094
rect -571 26079 -537 26094
rect -537 26079 -531 26094
rect -263 26094 -211 26131
rect -263 26079 -255 26094
rect -255 26079 -221 26094
rect -221 26079 -211 26094
rect -583 25806 -531 25841
rect -583 25789 -571 25806
rect -571 25789 -537 25806
rect -537 25789 -531 25806
rect 47 26094 99 26131
rect 47 26079 61 26094
rect 61 26079 95 26094
rect 95 26079 99 26094
rect -263 25806 -211 25841
rect -263 25789 -255 25806
rect -255 25789 -221 25806
rect -221 25789 -211 25806
rect -423 25556 -413 25571
rect -413 25556 -379 25571
rect -379 25556 -371 25571
rect -423 25519 -371 25556
rect 367 26094 419 26131
rect 367 26079 377 26094
rect 377 26079 411 26094
rect 411 26079 419 26094
rect 47 25806 99 25841
rect 47 25789 61 25806
rect 61 25789 95 25806
rect 95 25789 99 25806
rect -113 25556 -97 25571
rect -97 25556 -63 25571
rect -63 25556 -61 25571
rect -113 25519 -61 25556
rect -423 25268 -413 25281
rect -413 25268 -379 25281
rect -379 25268 -371 25281
rect -423 25230 -371 25268
rect -423 25229 -413 25230
rect -413 25229 -379 25230
rect -379 25229 -371 25230
rect 367 25806 419 25841
rect 367 25789 377 25806
rect 377 25789 411 25806
rect 411 25789 419 25806
rect 207 25556 219 25571
rect 219 25556 253 25571
rect 253 25556 259 25571
rect 207 25519 259 25556
rect -113 25268 -97 25281
rect -97 25268 -63 25281
rect -63 25268 -61 25281
rect -113 25230 -61 25268
rect -113 25229 -97 25230
rect -97 25229 -63 25230
rect -63 25229 -61 25230
rect 527 25556 535 25571
rect 535 25556 569 25571
rect 569 25556 579 25571
rect 527 25519 579 25556
rect 207 25268 219 25281
rect 219 25268 253 25281
rect 253 25268 259 25281
rect 207 25230 259 25268
rect 207 25229 219 25230
rect 219 25229 253 25230
rect 253 25229 259 25230
rect 527 25268 535 25281
rect 535 25268 569 25281
rect 569 25268 579 25281
rect 527 25230 579 25268
rect 527 25229 535 25230
rect 535 25229 569 25230
rect 569 25229 579 25230
rect -124 25041 120 25042
rect -124 25007 -90 25041
rect -90 25007 -56 25041
rect -56 25007 -18 25041
rect -18 25007 16 25041
rect 16 25007 54 25041
rect 54 25007 88 25041
rect 88 25007 120 25041
rect -124 24835 120 25007
rect -124 24801 -90 24835
rect -90 24801 -56 24835
rect -56 24801 -18 24835
rect -18 24801 16 24835
rect 16 24801 54 24835
rect 54 24801 88 24835
rect 88 24801 120 24835
rect -124 24798 120 24801
rect -583 24574 -531 24611
rect -583 24559 -571 24574
rect -571 24559 -537 24574
rect -537 24559 -531 24574
rect -263 24574 -211 24611
rect -263 24559 -255 24574
rect -255 24559 -221 24574
rect -221 24559 -211 24574
rect -583 24286 -531 24321
rect -583 24269 -571 24286
rect -571 24269 -537 24286
rect -537 24269 -531 24286
rect 47 24574 99 24611
rect 47 24559 61 24574
rect 61 24559 95 24574
rect 95 24559 99 24574
rect -263 24286 -211 24321
rect -263 24269 -255 24286
rect -255 24269 -221 24286
rect -221 24269 -211 24286
rect -423 24036 -413 24051
rect -413 24036 -379 24051
rect -379 24036 -371 24051
rect -423 23999 -371 24036
rect 367 24574 419 24611
rect 367 24559 377 24574
rect 377 24559 411 24574
rect 411 24559 419 24574
rect 47 24286 99 24321
rect 47 24269 61 24286
rect 61 24269 95 24286
rect 95 24269 99 24286
rect -113 24036 -97 24051
rect -97 24036 -63 24051
rect -63 24036 -61 24051
rect -113 23999 -61 24036
rect -423 23748 -413 23761
rect -413 23748 -379 23761
rect -379 23748 -371 23761
rect -423 23710 -371 23748
rect -423 23709 -413 23710
rect -413 23709 -379 23710
rect -379 23709 -371 23710
rect 367 24286 419 24321
rect 367 24269 377 24286
rect 377 24269 411 24286
rect 411 24269 419 24286
rect 207 24036 219 24051
rect 219 24036 253 24051
rect 253 24036 259 24051
rect 207 23999 259 24036
rect -113 23748 -97 23761
rect -97 23748 -63 23761
rect -63 23748 -61 23761
rect -113 23710 -61 23748
rect -113 23709 -97 23710
rect -97 23709 -63 23710
rect -63 23709 -61 23710
rect 527 24036 535 24051
rect 535 24036 569 24051
rect 569 24036 579 24051
rect 527 23999 579 24036
rect 207 23748 219 23761
rect 219 23748 253 23761
rect 253 23748 259 23761
rect 207 23710 259 23748
rect 207 23709 219 23710
rect 219 23709 253 23710
rect 253 23709 259 23710
rect 527 23748 535 23761
rect 535 23748 569 23761
rect 569 23748 579 23761
rect 527 23710 579 23748
rect 527 23709 535 23710
rect 535 23709 569 23710
rect 569 23709 579 23710
rect -124 23521 120 23522
rect -124 23487 -90 23521
rect -90 23487 -56 23521
rect -56 23487 -18 23521
rect -18 23487 16 23521
rect 16 23487 54 23521
rect 54 23487 88 23521
rect 88 23487 120 23521
rect -124 23314 120 23487
rect -124 23280 -86 23314
rect -86 23280 -52 23314
rect -52 23280 -14 23314
rect -14 23280 20 23314
rect 20 23280 58 23314
rect 58 23280 92 23314
rect 92 23280 120 23314
rect -124 23278 120 23280
rect -2363 23169 -2311 23221
rect -2113 23169 -2061 23221
rect 2037 23169 2089 23221
rect 2287 23169 2339 23221
rect -1573 23053 -1521 23091
rect -1573 23039 -1562 23053
rect -1562 23039 -1528 23053
rect -1528 23039 -1521 23053
rect -1053 23053 -1001 23091
rect -1053 23039 -1046 23053
rect -1046 23039 -1012 23053
rect -1012 23039 -1001 23053
rect -1573 22909 -1521 22911
rect -1573 22875 -1562 22909
rect -1562 22875 -1528 22909
rect -1528 22875 -1521 22909
rect -1573 22859 -1521 22875
rect -543 23053 -491 23091
rect -543 23039 -530 23053
rect -530 23039 -496 23053
rect -496 23039 -491 23053
rect -1053 22909 -1001 22911
rect -1053 22875 -1046 22909
rect -1046 22875 -1012 22909
rect -1012 22875 -1001 22909
rect -1053 22859 -1001 22875
rect -23 23053 29 23091
rect -23 23039 -14 23053
rect -14 23039 20 23053
rect 20 23039 29 23053
rect -1313 22405 -1261 22421
rect -1313 22371 -1304 22405
rect -1304 22371 -1270 22405
rect -1270 22371 -1261 22405
rect -1313 22369 -1261 22371
rect -543 22909 -491 22911
rect -543 22875 -530 22909
rect -530 22875 -496 22909
rect -496 22875 -491 22909
rect -543 22859 -491 22875
rect 487 23053 539 23091
rect 487 23039 502 23053
rect 502 23039 536 23053
rect 536 23039 539 23053
rect -803 22405 -751 22421
rect -803 22371 -788 22405
rect -788 22371 -754 22405
rect -754 22371 -751 22405
rect -803 22369 -751 22371
rect -23 22909 29 22911
rect -23 22875 -14 22909
rect -14 22875 20 22909
rect 20 22875 29 22909
rect -23 22859 29 22875
rect 1007 23053 1059 23091
rect 1007 23039 1018 23053
rect 1018 23039 1052 23053
rect 1052 23039 1059 23053
rect -1313 22227 -1304 22241
rect -1304 22227 -1270 22241
rect -1270 22227 -1261 22241
rect -1313 22189 -1261 22227
rect -283 22405 -231 22421
rect -283 22371 -272 22405
rect -272 22371 -238 22405
rect -238 22371 -231 22405
rect -283 22369 -231 22371
rect 487 22909 539 22911
rect 487 22875 502 22909
rect 502 22875 536 22909
rect 536 22875 539 22909
rect 487 22859 539 22875
rect 1527 23053 1579 23091
rect 1527 23039 1534 23053
rect 1534 23039 1568 23053
rect 1568 23039 1579 23053
rect -803 22227 -788 22241
rect -788 22227 -754 22241
rect -754 22227 -751 22241
rect -803 22189 -751 22227
rect 237 22405 289 22421
rect 237 22371 244 22405
rect 244 22371 278 22405
rect 278 22371 289 22405
rect 237 22369 289 22371
rect 1007 22909 1059 22911
rect 1007 22875 1018 22909
rect 1018 22875 1052 22909
rect 1052 22875 1059 22909
rect 1007 22859 1059 22875
rect -283 22227 -272 22241
rect -272 22227 -238 22241
rect -238 22227 -231 22241
rect -283 22189 -231 22227
rect 747 22405 799 22421
rect 747 22371 760 22405
rect 760 22371 794 22405
rect 794 22371 799 22405
rect 747 22369 799 22371
rect 1527 22909 1579 22911
rect 1527 22875 1534 22909
rect 1534 22875 1568 22909
rect 1568 22875 1579 22909
rect 1527 22859 1579 22875
rect 237 22227 244 22241
rect 244 22227 278 22241
rect 278 22227 289 22241
rect 237 22189 289 22227
rect 1267 22405 1319 22421
rect 1267 22371 1276 22405
rect 1276 22371 1310 22405
rect 1310 22371 1319 22405
rect 1267 22369 1319 22371
rect 747 22227 760 22241
rect 760 22227 794 22241
rect 794 22227 799 22241
rect 747 22189 799 22227
rect 1267 22227 1276 22241
rect 1276 22227 1310 22241
rect 1310 22227 1319 22241
rect 1267 22189 1319 22227
rect -2363 22059 -2311 22111
rect -2113 22059 -2061 22111
rect 2037 22059 2089 22111
rect 2287 22059 2339 22111
rect -119 22000 125 22007
rect -119 21966 -86 22000
rect -86 21966 -52 22000
rect -52 21966 -14 22000
rect -14 21966 20 22000
rect 20 21966 58 22000
rect 58 21966 92 22000
rect 92 21966 125 22000
rect -119 21794 125 21966
rect -119 21763 -90 21794
rect -90 21763 -52 21794
rect -52 21763 -18 21794
rect -18 21763 20 21794
rect 20 21763 54 21794
rect 54 21763 92 21794
rect 92 21763 125 21794
rect -3249 21344 -2685 21716
rect -2363 21649 -2311 21701
rect -2113 21649 -2061 21701
rect 2037 21649 2089 21701
rect 2287 21649 2339 21701
rect -1833 21533 -1781 21571
rect -1833 21519 -1822 21533
rect -1822 21519 -1788 21533
rect -1788 21519 -1781 21533
rect -1313 21533 -1261 21571
rect -1313 21519 -1306 21533
rect -1306 21519 -1272 21533
rect -1272 21519 -1261 21533
rect -1833 21389 -1781 21391
rect -1833 21355 -1822 21389
rect -1822 21355 -1788 21389
rect -1788 21355 -1781 21389
rect -1833 21339 -1781 21355
rect -803 21533 -751 21571
rect -803 21519 -790 21533
rect -790 21519 -756 21533
rect -756 21519 -751 21533
rect -1313 21389 -1261 21391
rect -1313 21355 -1306 21389
rect -1306 21355 -1272 21389
rect -1272 21355 -1261 21389
rect -1313 21339 -1261 21355
rect -283 21533 -231 21571
rect -283 21519 -274 21533
rect -274 21519 -240 21533
rect -240 21519 -231 21533
rect -1573 20885 -1521 20901
rect -1573 20851 -1564 20885
rect -1564 20851 -1530 20885
rect -1530 20851 -1521 20885
rect -1573 20849 -1521 20851
rect -803 21389 -751 21391
rect -803 21355 -790 21389
rect -790 21355 -756 21389
rect -756 21355 -751 21389
rect -803 21339 -751 21355
rect 227 21533 279 21571
rect 227 21519 242 21533
rect 242 21519 276 21533
rect 276 21519 279 21533
rect -1063 20885 -1011 20901
rect -1063 20851 -1048 20885
rect -1048 20851 -1014 20885
rect -1014 20851 -1011 20885
rect -1063 20849 -1011 20851
rect -283 21389 -231 21391
rect -283 21355 -274 21389
rect -274 21355 -240 21389
rect -240 21355 -231 21389
rect -283 21339 -231 21355
rect 747 21533 799 21571
rect 747 21519 758 21533
rect 758 21519 792 21533
rect 792 21519 799 21533
rect -1573 20707 -1564 20721
rect -1564 20707 -1530 20721
rect -1530 20707 -1521 20721
rect -1573 20669 -1521 20707
rect -543 20885 -491 20901
rect -543 20851 -532 20885
rect -532 20851 -498 20885
rect -498 20851 -491 20885
rect -543 20849 -491 20851
rect 227 21389 279 21391
rect 227 21355 242 21389
rect 242 21355 276 21389
rect 276 21355 279 21389
rect 227 21339 279 21355
rect 1267 21533 1319 21571
rect 1267 21519 1274 21533
rect 1274 21519 1308 21533
rect 1308 21519 1319 21533
rect -1063 20707 -1048 20721
rect -1048 20707 -1014 20721
rect -1014 20707 -1011 20721
rect -1063 20669 -1011 20707
rect -23 20885 29 20901
rect -23 20851 -16 20885
rect -16 20851 18 20885
rect 18 20851 29 20885
rect -23 20849 29 20851
rect 747 21389 799 21391
rect 747 21355 758 21389
rect 758 21355 792 21389
rect 792 21355 799 21389
rect 747 21339 799 21355
rect 1777 21533 1829 21571
rect 1777 21519 1790 21533
rect 1790 21519 1824 21533
rect 1824 21519 1829 21533
rect -543 20707 -532 20721
rect -532 20707 -498 20721
rect -498 20707 -491 20721
rect -543 20669 -491 20707
rect 487 20885 539 20901
rect 487 20851 500 20885
rect 500 20851 534 20885
rect 534 20851 539 20885
rect 487 20849 539 20851
rect 1267 21389 1319 21391
rect 1267 21355 1274 21389
rect 1274 21355 1308 21389
rect 1308 21355 1319 21389
rect 1267 21339 1319 21355
rect 2638 21440 2878 21680
rect 2968 21440 3208 21680
rect -23 20707 -16 20721
rect -16 20707 18 20721
rect 18 20707 29 20721
rect -23 20669 29 20707
rect 1007 20885 1059 20901
rect 1007 20851 1016 20885
rect 1016 20851 1050 20885
rect 1050 20851 1059 20885
rect 1007 20849 1059 20851
rect 1777 21389 1829 21391
rect 1777 21355 1790 21389
rect 1790 21355 1824 21389
rect 1824 21355 1829 21389
rect 1777 21339 1829 21355
rect 487 20707 500 20721
rect 500 20707 534 20721
rect 534 20707 539 20721
rect 487 20669 539 20707
rect 1517 20885 1569 20901
rect 1517 20851 1532 20885
rect 1532 20851 1566 20885
rect 1566 20851 1569 20885
rect 1517 20849 1569 20851
rect 1007 20707 1016 20721
rect 1016 20707 1050 20721
rect 1050 20707 1059 20721
rect 1007 20669 1059 20707
rect 1517 20707 1532 20721
rect 1532 20707 1566 20721
rect 1566 20707 1569 20721
rect 1517 20669 1569 20707
rect -2363 20539 -2311 20591
rect -2113 20539 -2061 20591
rect 2037 20539 2089 20591
rect 2287 20539 2339 20591
rect -119 20446 -90 20477
rect -90 20446 -52 20477
rect -52 20446 -18 20477
rect -18 20446 20 20477
rect 20 20446 54 20477
rect 54 20446 92 20477
rect 92 20446 125 20477
rect -119 20233 125 20446
rect -3220 19480 -3060 19640
rect -2160 19480 -2000 19640
rect -700 19480 -540 19640
rect 520 19480 680 19640
rect 2000 19480 2160 19640
rect 3000 19480 3160 19640
rect -1720 19250 -1650 19320
rect -1500 19250 -1430 19320
rect 1460 19250 1530 19320
rect 1700 19250 1770 19320
rect -3220 18900 -3060 19060
rect -2160 18900 -2000 19060
rect -700 18900 -540 19060
rect 520 18900 680 19060
rect 2000 18900 2160 19060
rect 3000 18900 3160 19060
rect -1720 18660 -1650 18730
rect -1500 18660 -1430 18730
rect 1460 18660 1530 18730
rect 1700 18660 1770 18730
rect -560 18550 -490 18570
rect -450 18550 -380 18570
rect 380 18550 450 18570
rect 490 18550 560 18570
rect -560 18500 -490 18550
rect -450 18500 -380 18550
rect 380 18500 450 18550
rect 490 18500 560 18550
rect -560 17990 -490 18000
rect -560 17930 -542 17990
rect -542 17930 -508 17990
rect -508 17930 -490 17990
rect -450 17990 -380 18000
rect 380 17990 450 18010
rect -450 17930 -434 17990
rect -434 17930 -400 17990
rect -400 17930 -380 17990
rect 380 17940 394 17990
rect 394 17940 428 17990
rect 428 17940 450 17990
rect 490 17990 560 18010
rect 490 17940 502 17990
rect 502 17940 536 17990
rect 536 17940 560 17990
rect -840 17530 -620 17680
rect -320 17530 -100 17680
rect 100 17530 320 17680
rect 650 17530 870 17680
rect -1720 17400 -1650 17470
rect -1510 17400 -1440 17470
rect 1460 17420 1530 17490
rect 1700 17420 1770 17490
rect -1720 17310 -1650 17380
rect -1510 17310 -1440 17380
rect 1460 17330 1530 17400
rect 1700 17330 1770 17400
rect -560 17235 -490 17250
rect -450 17235 -380 17250
rect 380 17235 450 17250
rect 490 17235 560 17250
rect -560 17180 -490 17235
rect -450 17180 -380 17235
rect 380 17180 450 17235
rect 490 17180 560 17235
rect -3200 16990 -3020 17120
rect -2060 16990 -1880 17120
rect -1080 17000 -900 17130
rect -310 17000 -130 17130
rect 130 17000 310 17130
rect 850 16990 1030 17120
rect 1920 17000 2100 17130
rect 2920 17000 3100 17130
rect -1720 16902 -1650 16950
rect -1500 16902 -1430 16950
rect 1460 16902 1530 16950
rect 1700 16902 1770 16950
rect -1720 16880 -1650 16902
rect -1500 16880 -1430 16902
rect 1460 16880 1530 16902
rect 1700 16880 1770 16902
rect -560 16730 -490 16800
rect -450 16730 -380 16800
rect 380 16730 450 16800
rect 490 16730 560 16800
rect -3240 15100 -3120 15220
rect 3130 15100 3250 15220
rect -3240 12100 -3120 12220
rect 3130 12100 3250 12220
rect -3240 9100 -3120 9220
rect 3130 9100 3250 9220
rect -3240 6100 -3120 6220
rect 3130 6100 3250 6220
rect -3240 3100 -3120 3220
rect 3130 3100 3250 3220
rect -2860 1518 -2827 1890
rect -2827 1518 -1713 1890
rect -1713 1518 -1690 1890
rect -2860 1480 -1690 1518
rect -1350 1518 -1307 1890
rect -1307 1518 -193 1890
rect -193 1518 -180 1890
rect -1350 1480 -180 1518
rect 170 1524 203 1890
rect 203 1524 1317 1890
rect 1317 1524 1340 1890
rect 170 1480 1340 1524
rect 1690 1524 1713 1900
rect 1713 1524 2827 1900
rect 2827 1524 2860 1900
rect 1690 1490 2860 1524
<< metal2 >>
rect -642 31387 -372 31410
rect -642 31143 -629 31387
rect -385 31143 -372 31387
rect -642 31120 -372 31143
rect 408 31387 678 31410
rect 408 31143 421 31387
rect 665 31143 678 31387
rect 408 31120 678 31143
rect -3192 30913 -3122 30930
rect -3192 30857 -3185 30913
rect -3129 30857 -3122 30913
rect -3192 30840 -3122 30857
rect -2872 30913 -2802 30930
rect -2872 30857 -2865 30913
rect -2809 30857 -2802 30913
rect -2872 30840 -2802 30857
rect -2562 30913 -2492 30930
rect -2562 30857 -2555 30913
rect -2499 30857 -2492 30913
rect -2562 30840 -2492 30857
rect -2242 30913 -2172 30930
rect -2242 30857 -2235 30913
rect -2179 30857 -2172 30913
rect -2242 30840 -2172 30857
rect -1932 30913 -1862 30930
rect -1932 30857 -1925 30913
rect -1869 30857 -1862 30913
rect -1932 30840 -1862 30857
rect -1612 30913 -1542 30930
rect -1612 30857 -1605 30913
rect -1549 30857 -1542 30913
rect -1612 30840 -1542 30857
rect -1292 30913 -1222 30930
rect -1292 30857 -1285 30913
rect -1229 30857 -1222 30913
rect -1292 30840 -1222 30857
rect -982 30913 -912 30930
rect -982 30857 -975 30913
rect -919 30857 -912 30913
rect -982 30840 -912 30857
rect -662 30913 -592 30930
rect -662 30857 -655 30913
rect -599 30857 -592 30913
rect -662 30840 -592 30857
rect -342 30913 -272 30930
rect -342 30857 -335 30913
rect -279 30857 -272 30913
rect -342 30840 -272 30857
rect -32 30913 38 30930
rect -32 30857 -25 30913
rect 31 30857 38 30913
rect -32 30840 38 30857
rect 288 30913 358 30930
rect 288 30857 295 30913
rect 351 30857 358 30913
rect 288 30840 358 30857
rect 598 30913 668 30930
rect 598 30857 605 30913
rect 661 30857 668 30913
rect 598 30840 668 30857
rect 918 30913 988 30930
rect 918 30857 925 30913
rect 981 30857 988 30913
rect 918 30840 988 30857
rect 1238 30913 1308 30930
rect 1238 30857 1245 30913
rect 1301 30857 1308 30913
rect 1238 30840 1308 30857
rect 1548 30913 1618 30930
rect 1548 30857 1555 30913
rect 1611 30857 1618 30913
rect 1548 30840 1618 30857
rect 1868 30913 1938 30930
rect 1868 30857 1875 30913
rect 1931 30857 1938 30913
rect 1868 30840 1938 30857
rect 2178 30913 2248 30930
rect 2178 30857 2185 30913
rect 2241 30857 2248 30913
rect 2178 30840 2248 30857
rect 2498 30913 2568 30930
rect 2498 30857 2505 30913
rect 2561 30857 2568 30913
rect 2498 30840 2568 30857
rect 2818 30913 2888 30930
rect 2818 30857 2825 30913
rect 2881 30857 2888 30913
rect 2818 30840 2888 30857
rect 3128 30913 3198 30930
rect 3128 30857 3135 30913
rect 3191 30857 3198 30913
rect 3128 30840 3198 30857
rect -3192 30673 -3122 30690
rect -7912 30620 -7852 30630
rect -7912 30550 -7852 30560
rect -7792 30620 -7732 30630
rect -3192 30617 -3185 30673
rect -3129 30617 -3122 30673
rect -3192 30600 -3122 30617
rect -2872 30673 -2802 30690
rect -2872 30617 -2865 30673
rect -2809 30617 -2802 30673
rect -2872 30600 -2802 30617
rect -2562 30673 -2492 30690
rect -2562 30617 -2555 30673
rect -2499 30617 -2492 30673
rect -2562 30600 -2492 30617
rect -2242 30673 -2172 30690
rect -2242 30617 -2235 30673
rect -2179 30617 -2172 30673
rect -2242 30600 -2172 30617
rect -1932 30673 -1862 30690
rect -1932 30617 -1925 30673
rect -1869 30617 -1862 30673
rect -1932 30600 -1862 30617
rect -1612 30673 -1542 30690
rect -1612 30617 -1605 30673
rect -1549 30617 -1542 30673
rect -1612 30600 -1542 30617
rect -1292 30673 -1222 30690
rect -1292 30617 -1285 30673
rect -1229 30617 -1222 30673
rect -1292 30600 -1222 30617
rect -982 30673 -912 30690
rect -982 30617 -975 30673
rect -919 30617 -912 30673
rect -982 30600 -912 30617
rect -662 30673 -592 30690
rect -662 30617 -655 30673
rect -599 30617 -592 30673
rect -662 30600 -592 30617
rect -342 30673 -272 30690
rect -342 30617 -335 30673
rect -279 30617 -272 30673
rect -342 30600 -272 30617
rect -32 30673 38 30690
rect -32 30617 -25 30673
rect 31 30617 38 30673
rect -32 30600 38 30617
rect 288 30673 358 30690
rect 288 30617 295 30673
rect 351 30617 358 30673
rect 288 30600 358 30617
rect 598 30673 668 30690
rect 598 30617 605 30673
rect 661 30617 668 30673
rect 598 30600 668 30617
rect 918 30673 988 30690
rect 918 30617 925 30673
rect 981 30617 988 30673
rect 918 30600 988 30617
rect 1238 30673 1308 30690
rect 1238 30617 1245 30673
rect 1301 30617 1308 30673
rect 1238 30600 1308 30617
rect 1548 30673 1618 30690
rect 1548 30617 1555 30673
rect 1611 30617 1618 30673
rect 1548 30600 1618 30617
rect 1868 30673 1938 30690
rect 1868 30617 1875 30673
rect 1931 30617 1938 30673
rect 1868 30600 1938 30617
rect 2178 30673 2248 30690
rect 2178 30617 2185 30673
rect 2241 30617 2248 30673
rect 2178 30600 2248 30617
rect 2498 30673 2568 30690
rect 2498 30617 2505 30673
rect 2561 30617 2568 30673
rect 2498 30600 2568 30617
rect 2818 30673 2888 30690
rect 2818 30617 2825 30673
rect 2881 30617 2888 30673
rect 2818 30600 2888 30617
rect 3128 30673 3198 30690
rect 3128 30617 3135 30673
rect 3191 30617 3198 30673
rect 3128 30600 3198 30617
rect 7988 30618 8068 30640
rect -7792 30550 -7732 30560
rect 7988 30562 8000 30618
rect 8056 30562 8068 30618
rect 7988 30540 8068 30562
rect 8098 30618 8178 30640
rect 8098 30562 8110 30618
rect 8166 30562 8178 30618
rect 8098 30540 8178 30562
rect -3062 30303 -2932 30320
rect -3062 30247 -3025 30303
rect -2969 30247 -2932 30303
rect -3062 30063 -2932 30247
rect -2722 30303 -2652 30320
rect -2722 30247 -2715 30303
rect -2659 30247 -2652 30303
rect -2722 30230 -2652 30247
rect -2402 30303 -2332 30320
rect -2402 30247 -2395 30303
rect -2339 30247 -2332 30303
rect -2402 30230 -2332 30247
rect -2082 30303 -2012 30320
rect -2082 30247 -2075 30303
rect -2019 30247 -2012 30303
rect -2082 30230 -2012 30247
rect -1772 30303 -1702 30320
rect -1772 30247 -1765 30303
rect -1709 30247 -1702 30303
rect -1772 30230 -1702 30247
rect -1452 30303 -1382 30320
rect -1452 30247 -1445 30303
rect -1389 30247 -1382 30303
rect -1452 30230 -1382 30247
rect -1142 30303 -1072 30320
rect -1142 30247 -1135 30303
rect -1079 30247 -1072 30303
rect -1142 30230 -1072 30247
rect -822 30303 -752 30320
rect -822 30247 -815 30303
rect -759 30247 -752 30303
rect -822 30230 -752 30247
rect -502 30303 -432 30320
rect -502 30247 -495 30303
rect -439 30247 -432 30303
rect -502 30230 -432 30247
rect -192 30303 -122 30320
rect -192 30247 -185 30303
rect -129 30247 -122 30303
rect -192 30230 -122 30247
rect 128 30303 198 30320
rect 128 30247 135 30303
rect 191 30247 198 30303
rect 128 30230 198 30247
rect 448 30303 518 30320
rect 448 30247 455 30303
rect 511 30247 518 30303
rect 448 30230 518 30247
rect 758 30303 828 30320
rect 758 30247 765 30303
rect 821 30247 828 30303
rect 758 30230 828 30247
rect 1078 30303 1148 30320
rect 1078 30247 1085 30303
rect 1141 30247 1148 30303
rect 1078 30230 1148 30247
rect 1388 30303 1458 30320
rect 1388 30247 1395 30303
rect 1451 30247 1458 30303
rect 1388 30230 1458 30247
rect 1708 30303 1778 30320
rect 1708 30247 1715 30303
rect 1771 30247 1778 30303
rect 1708 30230 1778 30247
rect 2028 30303 2098 30320
rect 2028 30247 2035 30303
rect 2091 30247 2098 30303
rect 2028 30230 2098 30247
rect 2338 30303 2408 30320
rect 2338 30247 2345 30303
rect 2401 30247 2408 30303
rect 2338 30230 2408 30247
rect 2658 30303 2728 30320
rect 2658 30247 2665 30303
rect 2721 30247 2728 30303
rect 2658 30230 2728 30247
rect 2948 30303 3078 30320
rect 2948 30247 2985 30303
rect 3041 30247 3078 30303
rect -3062 30007 -3025 30063
rect -2969 30007 -2932 30063
rect -3062 29693 -2932 30007
rect -2722 30063 -2652 30080
rect -2722 30007 -2715 30063
rect -2659 30007 -2652 30063
rect -2722 29990 -2652 30007
rect -2402 30063 -2332 30080
rect -2402 30007 -2395 30063
rect -2339 30007 -2332 30063
rect -2402 29990 -2332 30007
rect -2082 30063 -2012 30080
rect -2082 30007 -2075 30063
rect -2019 30007 -2012 30063
rect -2082 29990 -2012 30007
rect -1772 30063 -1702 30080
rect -1772 30007 -1765 30063
rect -1709 30007 -1702 30063
rect -1772 29990 -1702 30007
rect -1452 30063 -1382 30080
rect -1452 30007 -1445 30063
rect -1389 30007 -1382 30063
rect -1452 29990 -1382 30007
rect -1142 30063 -1072 30080
rect -1142 30007 -1135 30063
rect -1079 30007 -1072 30063
rect -1142 29990 -1072 30007
rect -822 30063 -752 30080
rect -822 30007 -815 30063
rect -759 30007 -752 30063
rect -822 29990 -752 30007
rect -502 30063 -432 30080
rect -502 30007 -495 30063
rect -439 30007 -432 30063
rect -502 29990 -432 30007
rect -192 30063 -122 30080
rect -192 30007 -185 30063
rect -129 30007 -122 30063
rect -192 29990 -122 30007
rect 128 30063 198 30080
rect 128 30007 135 30063
rect 191 30007 198 30063
rect 128 29990 198 30007
rect 448 30063 518 30080
rect 448 30007 455 30063
rect 511 30007 518 30063
rect 448 29990 518 30007
rect 758 30063 828 30080
rect 758 30007 765 30063
rect 821 30007 828 30063
rect 758 29990 828 30007
rect 1078 30063 1148 30080
rect 1078 30007 1085 30063
rect 1141 30007 1148 30063
rect 1078 29990 1148 30007
rect 1388 30063 1458 30080
rect 1388 30007 1395 30063
rect 1451 30007 1458 30063
rect 1388 29990 1458 30007
rect 1708 30063 1778 30080
rect 1708 30007 1715 30063
rect 1771 30007 1778 30063
rect 1708 29990 1778 30007
rect 2028 30063 2098 30080
rect 2028 30007 2035 30063
rect 2091 30007 2098 30063
rect 2028 29990 2098 30007
rect 2338 30063 2408 30080
rect 2338 30007 2345 30063
rect 2401 30007 2408 30063
rect 2338 29990 2408 30007
rect 2658 30063 2728 30080
rect 2658 30007 2665 30063
rect 2721 30007 2728 30063
rect 2658 29990 2728 30007
rect 2948 30063 3078 30247
rect 2948 30007 2985 30063
rect 3041 30007 3078 30063
rect -3062 29637 -3025 29693
rect -2969 29637 -2932 29693
rect -3062 23083 -2932 29637
rect -2112 29886 -1952 29920
rect -2112 29834 -2058 29886
rect -2006 29834 -1952 29886
rect -2112 28588 -1952 29834
rect 1948 29886 2108 29920
rect 1948 29834 2002 29886
rect 2054 29834 2108 29886
rect -642 29747 -372 29770
rect -642 29503 -629 29747
rect -385 29503 -372 29747
rect -642 29480 -372 29503
rect 408 29747 678 29770
rect 408 29503 421 29747
rect 665 29503 678 29747
rect 408 29480 678 29503
rect -1692 29243 -1622 29260
rect -1692 29187 -1685 29243
rect -1629 29187 -1622 29243
rect -1692 29170 -1622 29187
rect -1372 29243 -1302 29260
rect -1372 29187 -1365 29243
rect -1309 29187 -1302 29243
rect -1372 29170 -1302 29187
rect -1062 29243 -992 29260
rect -1062 29187 -1055 29243
rect -999 29187 -992 29243
rect -1062 29170 -992 29187
rect -742 29243 -672 29260
rect -742 29187 -735 29243
rect -679 29187 -672 29243
rect -742 29170 -672 29187
rect -422 29243 -352 29260
rect -422 29187 -415 29243
rect -359 29187 -352 29243
rect -422 29170 -352 29187
rect -112 29243 -42 29260
rect -112 29187 -105 29243
rect -49 29187 -42 29243
rect -112 29170 -42 29187
rect 208 29243 278 29260
rect 208 29187 215 29243
rect 271 29187 278 29243
rect 208 29170 278 29187
rect 528 29243 598 29260
rect 528 29187 535 29243
rect 591 29187 598 29243
rect 528 29170 598 29187
rect 838 29243 908 29260
rect 838 29187 845 29243
rect 901 29187 908 29243
rect 838 29170 908 29187
rect 1158 29243 1228 29260
rect 1158 29187 1165 29243
rect 1221 29187 1228 29243
rect 1158 29170 1228 29187
rect 1468 29243 1538 29260
rect 1468 29187 1475 29243
rect 1531 29187 1538 29243
rect 1468 29170 1538 29187
rect -1692 29033 -1622 29050
rect -1692 28977 -1685 29033
rect -1629 28977 -1622 29033
rect -1692 28960 -1622 28977
rect -1372 29033 -1302 29050
rect -1372 28977 -1365 29033
rect -1309 28977 -1302 29033
rect -1372 28960 -1302 28977
rect -1062 29033 -992 29050
rect -1062 28977 -1055 29033
rect -999 28977 -992 29033
rect -1062 28960 -992 28977
rect -742 29033 -672 29050
rect -742 28977 -735 29033
rect -679 28977 -672 29033
rect -742 28960 -672 28977
rect -422 29033 -352 29050
rect -422 28977 -415 29033
rect -359 28977 -352 29033
rect -422 28960 -352 28977
rect -112 29033 -42 29050
rect -112 28977 -105 29033
rect -49 28977 -42 29033
rect -112 28960 -42 28977
rect 208 29033 278 29050
rect 208 28977 215 29033
rect 271 28977 278 29033
rect 208 28960 278 28977
rect 528 29033 598 29050
rect 528 28977 535 29033
rect 591 28977 598 29033
rect 528 28960 598 28977
rect 838 29033 908 29050
rect 838 28977 845 29033
rect 901 28977 908 29033
rect 838 28960 908 28977
rect 1158 29033 1228 29050
rect 1158 28977 1165 29033
rect 1221 28977 1228 29033
rect 1158 28960 1228 28977
rect 1468 29033 1538 29050
rect 1468 28977 1475 29033
rect 1531 28977 1538 29033
rect 1468 28960 1538 28977
rect -2112 28532 -2060 28588
rect -2004 28532 -1952 28588
rect -2112 28408 -1952 28532
rect -1532 28603 -1462 28620
rect -1532 28547 -1525 28603
rect -1469 28547 -1462 28603
rect -1532 28530 -1462 28547
rect -1212 28603 -1142 28620
rect -1212 28547 -1205 28603
rect -1149 28547 -1142 28603
rect -1212 28530 -1142 28547
rect -902 28603 -832 28620
rect -902 28547 -895 28603
rect -839 28547 -832 28603
rect -902 28530 -832 28547
rect -582 28603 -512 28620
rect -582 28547 -575 28603
rect -519 28547 -512 28603
rect -582 28530 -512 28547
rect -262 28603 -192 28620
rect -262 28547 -255 28603
rect -199 28547 -192 28603
rect -262 28530 -192 28547
rect 48 28603 118 28620
rect 48 28547 55 28603
rect 111 28547 118 28603
rect 48 28530 118 28547
rect 368 28603 438 28620
rect 368 28547 375 28603
rect 431 28547 438 28603
rect 368 28530 438 28547
rect 678 28603 748 28620
rect 678 28547 685 28603
rect 741 28547 748 28603
rect 678 28530 748 28547
rect 998 28603 1068 28620
rect 998 28547 1005 28603
rect 1061 28547 1068 28603
rect 998 28530 1068 28547
rect 1318 28603 1388 28620
rect 1318 28547 1325 28603
rect 1381 28547 1388 28603
rect 1318 28530 1388 28547
rect 1628 28603 1698 28620
rect 1628 28547 1635 28603
rect 1691 28547 1698 28603
rect 1628 28530 1698 28547
rect 1948 28588 2108 29834
rect 1948 28532 2000 28588
rect 2056 28532 2108 28588
rect -2112 28352 -2060 28408
rect -2004 28352 -1952 28408
rect -2112 26098 -1952 28352
rect -1532 28393 -1462 28410
rect -1532 28337 -1525 28393
rect -1469 28337 -1462 28393
rect -1532 28320 -1462 28337
rect -1212 28393 -1142 28410
rect -1212 28337 -1205 28393
rect -1149 28337 -1142 28393
rect -1212 28320 -1142 28337
rect -902 28393 -832 28410
rect -902 28337 -895 28393
rect -839 28337 -832 28393
rect -902 28320 -832 28337
rect -582 28393 -512 28410
rect -582 28337 -575 28393
rect -519 28337 -512 28393
rect -582 28320 -512 28337
rect -262 28393 -192 28410
rect -262 28337 -255 28393
rect -199 28337 -192 28393
rect -262 28320 -192 28337
rect 48 28393 118 28410
rect 48 28337 55 28393
rect 111 28337 118 28393
rect 48 28320 118 28337
rect 368 28393 438 28410
rect 368 28337 375 28393
rect 431 28337 438 28393
rect 368 28320 438 28337
rect 678 28393 748 28410
rect 678 28337 685 28393
rect 741 28337 748 28393
rect 678 28320 748 28337
rect 998 28393 1068 28410
rect 998 28337 1005 28393
rect 1061 28337 1068 28393
rect 998 28320 1068 28337
rect 1318 28393 1388 28410
rect 1318 28337 1325 28393
rect 1381 28337 1388 28393
rect 1318 28320 1388 28337
rect 1628 28393 1698 28410
rect 1628 28337 1635 28393
rect 1691 28337 1698 28393
rect 1628 28320 1698 28337
rect 1948 28408 2108 28532
rect 1948 28352 2000 28408
rect 2056 28352 2108 28408
rect -872 28142 -612 28160
rect -872 27898 -864 28142
rect -620 27898 -612 28142
rect -872 27880 -612 27898
rect 628 28142 888 28160
rect 628 27898 636 28142
rect 880 27898 888 28142
rect 628 27880 888 27898
rect -1692 27693 -1622 27710
rect -1692 27637 -1685 27693
rect -1629 27637 -1622 27693
rect -1692 27620 -1622 27637
rect -1372 27693 -1302 27710
rect -1372 27637 -1365 27693
rect -1309 27637 -1302 27693
rect -1372 27620 -1302 27637
rect -1062 27693 -992 27710
rect -1062 27637 -1055 27693
rect -999 27637 -992 27693
rect -1062 27620 -992 27637
rect -742 27693 -672 27710
rect -742 27637 -735 27693
rect -679 27637 -672 27693
rect -742 27620 -672 27637
rect -422 27693 -352 27710
rect -422 27637 -415 27693
rect -359 27637 -352 27693
rect -422 27620 -352 27637
rect -112 27693 -42 27710
rect -112 27637 -105 27693
rect -49 27637 -42 27693
rect -112 27620 -42 27637
rect 208 27693 278 27710
rect 208 27637 215 27693
rect 271 27637 278 27693
rect 208 27620 278 27637
rect 518 27693 588 27710
rect 518 27637 525 27693
rect 581 27637 588 27693
rect 518 27620 588 27637
rect 838 27693 908 27710
rect 838 27637 845 27693
rect 901 27637 908 27693
rect 838 27620 908 27637
rect 1158 27693 1228 27710
rect 1158 27637 1165 27693
rect 1221 27637 1228 27693
rect 1158 27620 1228 27637
rect 1468 27693 1538 27710
rect 1468 27637 1475 27693
rect 1531 27637 1538 27693
rect 1468 27620 1538 27637
rect -1692 27483 -1622 27500
rect -1692 27427 -1685 27483
rect -1629 27427 -1622 27483
rect -1692 27410 -1622 27427
rect -1372 27483 -1302 27500
rect -1372 27427 -1365 27483
rect -1309 27427 -1302 27483
rect -1372 27410 -1302 27427
rect -1062 27483 -992 27500
rect -1062 27427 -1055 27483
rect -999 27427 -992 27483
rect -1062 27410 -992 27427
rect -742 27483 -672 27500
rect -742 27427 -735 27483
rect -679 27427 -672 27483
rect -742 27410 -672 27427
rect -422 27483 -352 27500
rect -422 27427 -415 27483
rect -359 27427 -352 27483
rect -422 27410 -352 27427
rect -112 27483 -42 27500
rect -112 27427 -105 27483
rect -49 27427 -42 27483
rect -112 27410 -42 27427
rect 208 27483 278 27500
rect 208 27427 215 27483
rect 271 27427 278 27483
rect 208 27410 278 27427
rect 518 27483 588 27500
rect 518 27427 525 27483
rect 581 27427 588 27483
rect 518 27410 588 27427
rect 838 27483 908 27500
rect 838 27427 845 27483
rect 901 27427 908 27483
rect 838 27410 908 27427
rect 1158 27483 1228 27500
rect 1158 27427 1165 27483
rect 1221 27427 1228 27483
rect 1158 27410 1228 27427
rect 1468 27483 1538 27500
rect 1468 27427 1475 27483
rect 1531 27427 1538 27483
rect 1468 27410 1538 27427
rect -1532 27063 -1462 27080
rect -1532 27007 -1525 27063
rect -1469 27007 -1462 27063
rect -1532 26990 -1462 27007
rect -1242 27063 -1112 27080
rect -1242 27007 -1205 27063
rect -1149 27007 -1112 27063
rect -1532 26853 -1462 26870
rect -1532 26797 -1525 26853
rect -1469 26797 -1462 26853
rect -1532 26780 -1462 26797
rect -1242 26853 -1112 27007
rect -902 27063 -832 27080
rect -902 27007 -895 27063
rect -839 27007 -832 27063
rect -902 26990 -832 27007
rect -582 27063 -512 27080
rect -582 27007 -575 27063
rect -519 27007 -512 27063
rect -582 26990 -512 27007
rect -272 27063 -202 27080
rect -272 27007 -265 27063
rect -209 27007 -202 27063
rect -272 26990 -202 27007
rect 48 27063 118 27080
rect 48 27007 55 27063
rect 111 27007 118 27063
rect 48 26990 118 27007
rect 368 27063 438 27080
rect 368 27007 375 27063
rect 431 27007 438 27063
rect 368 26990 438 27007
rect 678 27063 748 27080
rect 678 27007 685 27063
rect 741 27007 748 27063
rect 678 26990 748 27007
rect 998 27063 1068 27080
rect 998 27007 1005 27063
rect 1061 27007 1068 27063
rect 998 26990 1068 27007
rect 1278 27063 1408 27080
rect 1278 27007 1315 27063
rect 1371 27007 1408 27063
rect -1242 26797 -1205 26853
rect -1149 26797 -1112 26853
rect -2112 26042 -2060 26098
rect -2004 26042 -1952 26098
rect -2112 25878 -1952 26042
rect -2112 25822 -2060 25878
rect -2004 25822 -1952 25878
rect -2112 25770 -1952 25822
rect -1872 25538 -1712 25590
rect -1872 25482 -1820 25538
rect -1764 25482 -1712 25538
rect -1872 25318 -1712 25482
rect -1872 25262 -1820 25318
rect -1764 25262 -1712 25318
rect -1872 24578 -1712 25262
rect -1872 24522 -1820 24578
rect -1764 24522 -1712 24578
rect -1872 24358 -1712 24522
rect -1872 24302 -1820 24358
rect -1764 24302 -1712 24358
rect -3062 23027 -3025 23083
rect -2969 23027 -2932 23083
rect -3062 22923 -2932 23027
rect -3062 22867 -3025 22923
rect -2969 22867 -2932 22923
rect -3062 22840 -2932 22867
rect -2412 23221 -2012 23370
rect -2412 23169 -2363 23221
rect -2311 23169 -2113 23221
rect -2061 23169 -2012 23221
rect -2412 22111 -2012 23169
rect -2412 22059 -2363 22111
rect -2311 22059 -2113 22111
rect -2061 22059 -2012 22111
rect -3262 21718 -2672 21750
rect -3262 21716 -3235 21718
rect -2699 21716 -2672 21718
rect -3262 21344 -3249 21716
rect -2685 21344 -2672 21716
rect -3262 21342 -3235 21344
rect -2699 21342 -2672 21344
rect -3262 21310 -2672 21342
rect -2412 21701 -2012 22059
rect -2412 21649 -2363 21701
rect -2311 21649 -2113 21701
rect -2061 21649 -2012 21701
rect -2412 20591 -2012 21649
rect -1872 21573 -1712 24302
rect -1242 24033 -1112 26797
rect -902 26853 -832 26870
rect -902 26797 -895 26853
rect -839 26797 -832 26853
rect -902 26780 -832 26797
rect -582 26853 -512 26870
rect -582 26797 -575 26853
rect -519 26797 -512 26853
rect -582 26780 -512 26797
rect -272 26853 -202 26870
rect -272 26797 -265 26853
rect -209 26797 -202 26853
rect -272 26780 -202 26797
rect 48 26853 118 26870
rect 48 26797 55 26853
rect 111 26797 118 26853
rect 48 26780 118 26797
rect 368 26853 438 26870
rect 368 26797 375 26853
rect 431 26797 438 26853
rect 368 26780 438 26797
rect 678 26853 748 26870
rect 678 26797 685 26853
rect 741 26797 748 26853
rect 678 26780 748 26797
rect 998 26853 1068 26870
rect 998 26797 1005 26853
rect 1061 26797 1068 26853
rect 998 26780 1068 26797
rect 1278 26853 1408 27007
rect 1628 27063 1698 27080
rect 1628 27007 1635 27063
rect 1691 27007 1698 27063
rect 1628 26990 1698 27007
rect 1278 26797 1315 26853
rect 1371 26797 1408 26853
rect -592 26133 -522 26150
rect -592 26077 -585 26133
rect -529 26077 -522 26133
rect -592 26060 -522 26077
rect -272 26133 -202 26150
rect -272 26077 -265 26133
rect -209 26077 -202 26133
rect -272 26060 -202 26077
rect 38 26133 108 26150
rect 38 26077 45 26133
rect 101 26077 108 26133
rect 38 26060 108 26077
rect 358 26133 428 26150
rect 358 26077 365 26133
rect 421 26077 428 26133
rect 358 26060 428 26077
rect -592 25843 -522 25860
rect -592 25787 -585 25843
rect -529 25787 -522 25843
rect -592 25770 -522 25787
rect -272 25843 -202 25860
rect -272 25787 -265 25843
rect -209 25787 -202 25843
rect -272 25770 -202 25787
rect 38 25843 108 25860
rect 38 25787 45 25843
rect 101 25787 108 25843
rect 38 25770 108 25787
rect 358 25843 428 25860
rect 358 25787 365 25843
rect 421 25787 428 25843
rect 358 25770 428 25787
rect -432 25573 -362 25590
rect -432 25517 -425 25573
rect -369 25517 -362 25573
rect -432 25500 -362 25517
rect -122 25573 -52 25590
rect -122 25517 -115 25573
rect -59 25517 -52 25573
rect -122 25500 -52 25517
rect 198 25573 268 25590
rect 198 25517 205 25573
rect 261 25517 268 25573
rect 198 25500 268 25517
rect 518 25573 588 25590
rect 518 25517 525 25573
rect 581 25517 588 25573
rect 518 25500 588 25517
rect -432 25283 -362 25300
rect -432 25227 -425 25283
rect -369 25227 -362 25283
rect -432 25210 -362 25227
rect -122 25283 -52 25300
rect -122 25227 -115 25283
rect -59 25227 -52 25283
rect -122 25210 -52 25227
rect 198 25283 268 25300
rect 198 25227 205 25283
rect 261 25227 268 25283
rect 198 25210 268 25227
rect 518 25283 588 25300
rect 518 25227 525 25283
rect 581 25227 588 25283
rect 518 25210 588 25227
rect -132 25042 128 25060
rect -132 24798 -124 25042
rect 120 24798 128 25042
rect -132 24780 128 24798
rect -592 24613 -522 24630
rect -592 24557 -585 24613
rect -529 24557 -522 24613
rect -592 24540 -522 24557
rect -272 24613 -202 24630
rect -272 24557 -265 24613
rect -209 24557 -202 24613
rect -272 24540 -202 24557
rect 38 24613 108 24630
rect 38 24557 45 24613
rect 101 24557 108 24613
rect 38 24540 108 24557
rect 358 24613 428 24630
rect 358 24557 365 24613
rect 421 24557 428 24613
rect 358 24540 428 24557
rect -592 24323 -522 24340
rect -592 24267 -585 24323
rect -529 24267 -522 24323
rect -592 24250 -522 24267
rect -272 24323 -202 24340
rect -272 24267 -265 24323
rect -209 24267 -202 24323
rect -272 24250 -202 24267
rect 38 24323 108 24340
rect 38 24267 45 24323
rect 101 24267 108 24323
rect 38 24250 108 24267
rect 358 24323 428 24340
rect 358 24267 365 24323
rect 421 24267 428 24323
rect 358 24250 428 24267
rect -1242 23977 -1205 24033
rect -1149 23977 -1112 24033
rect -432 24053 -362 24070
rect -432 23997 -425 24053
rect -369 23997 -362 24053
rect -432 23980 -362 23997
rect -122 24053 -52 24070
rect -122 23997 -115 24053
rect -59 23997 -52 24053
rect -122 23980 -52 23997
rect 198 24053 268 24070
rect 198 23997 205 24053
rect 261 23997 268 24053
rect 198 23980 268 23997
rect 518 24053 588 24070
rect 518 23997 525 24053
rect 581 23997 588 24053
rect 518 23980 588 23997
rect 1278 24033 1408 26797
rect 1628 26853 1698 26870
rect 1628 26797 1635 26853
rect 1691 26797 1698 26853
rect 1628 26780 1698 26797
rect 1948 26098 2108 28352
rect 1948 26042 2000 26098
rect 2056 26042 2108 26098
rect 1948 25878 2108 26042
rect 1948 25822 2000 25878
rect 2056 25822 2108 25878
rect 1948 25770 2108 25822
rect 2948 29693 3078 30007
rect 2948 29637 2985 29693
rect 3041 29637 3078 29693
rect -1242 23783 -1112 23977
rect -1242 23727 -1205 23783
rect -1149 23727 -1112 23783
rect 1278 23977 1315 24033
rect 1371 23977 1408 24033
rect 1278 23783 1408 23977
rect -1242 23690 -1112 23727
rect -432 23763 -362 23780
rect -432 23707 -425 23763
rect -369 23707 -362 23763
rect -432 23690 -362 23707
rect -122 23763 -52 23780
rect -122 23707 -115 23763
rect -59 23707 -52 23763
rect -122 23690 -52 23707
rect 198 23763 268 23780
rect 198 23707 205 23763
rect 261 23707 268 23763
rect 198 23690 268 23707
rect 518 23763 588 23780
rect 518 23707 525 23763
rect 581 23707 588 23763
rect 518 23690 588 23707
rect 1278 23727 1315 23783
rect 1371 23727 1408 23783
rect 1278 23690 1408 23727
rect 1708 25538 1868 25590
rect 1708 25482 1760 25538
rect 1816 25482 1868 25538
rect 1708 25318 1868 25482
rect 1708 25262 1760 25318
rect 1816 25262 1868 25318
rect 1708 24578 1868 25262
rect 1708 24522 1760 24578
rect 1816 24522 1868 24578
rect 1708 24358 1868 24522
rect 1708 24302 1760 24358
rect 1816 24302 1868 24358
rect -132 23522 128 23540
rect -132 23278 -124 23522
rect 120 23278 128 23522
rect -132 23260 128 23278
rect -1582 23093 -1512 23110
rect -1582 23037 -1575 23093
rect -1519 23037 -1512 23093
rect -1582 23020 -1512 23037
rect -1062 23093 -992 23110
rect -1062 23037 -1055 23093
rect -999 23037 -992 23093
rect -1062 23020 -992 23037
rect -552 23093 -482 23110
rect -552 23037 -545 23093
rect -489 23037 -482 23093
rect -552 23020 -482 23037
rect -32 23093 38 23110
rect -32 23037 -25 23093
rect 31 23037 38 23093
rect -32 23020 38 23037
rect 478 23093 548 23110
rect 478 23037 485 23093
rect 541 23037 548 23093
rect 478 23020 548 23037
rect 998 23093 1068 23110
rect 998 23037 1005 23093
rect 1061 23037 1068 23093
rect 998 23020 1068 23037
rect 1518 23093 1588 23110
rect 1518 23037 1525 23093
rect 1581 23037 1588 23093
rect 1518 23020 1588 23037
rect -1582 22913 -1512 22930
rect -1582 22857 -1575 22913
rect -1519 22857 -1512 22913
rect -1582 22840 -1512 22857
rect -1062 22913 -992 22930
rect -1062 22857 -1055 22913
rect -999 22857 -992 22913
rect -1062 22840 -992 22857
rect -552 22913 -482 22930
rect -552 22857 -545 22913
rect -489 22857 -482 22913
rect -552 22840 -482 22857
rect -32 22913 38 22930
rect -32 22857 -25 22913
rect 31 22857 38 22913
rect -32 22840 38 22857
rect 478 22913 548 22930
rect 478 22857 485 22913
rect 541 22857 548 22913
rect 478 22840 548 22857
rect 998 22913 1068 22930
rect 998 22857 1005 22913
rect 1061 22857 1068 22913
rect 998 22840 1068 22857
rect 1518 22913 1588 22930
rect 1518 22857 1525 22913
rect 1581 22857 1588 22913
rect 1518 22840 1588 22857
rect -1322 22423 -1252 22440
rect -1322 22367 -1315 22423
rect -1259 22367 -1252 22423
rect -1322 22350 -1252 22367
rect -812 22423 -742 22440
rect -812 22367 -805 22423
rect -749 22367 -742 22423
rect -812 22350 -742 22367
rect -292 22423 -222 22440
rect -292 22367 -285 22423
rect -229 22367 -222 22423
rect -292 22350 -222 22367
rect 228 22423 298 22440
rect 228 22367 235 22423
rect 291 22367 298 22423
rect 228 22350 298 22367
rect 738 22423 808 22440
rect 738 22367 745 22423
rect 801 22367 808 22423
rect 738 22350 808 22367
rect 1258 22423 1328 22440
rect 1258 22367 1265 22423
rect 1321 22367 1328 22423
rect 1258 22350 1328 22367
rect -1322 22243 -1252 22260
rect -1322 22187 -1315 22243
rect -1259 22187 -1252 22243
rect -1322 22170 -1252 22187
rect -812 22243 -742 22260
rect -812 22187 -805 22243
rect -749 22187 -742 22243
rect -812 22170 -742 22187
rect -292 22243 -222 22260
rect -292 22187 -285 22243
rect -229 22187 -222 22243
rect -292 22170 -222 22187
rect 228 22243 298 22260
rect 228 22187 235 22243
rect 291 22187 298 22243
rect 228 22170 298 22187
rect 738 22243 808 22260
rect 738 22187 745 22243
rect 801 22187 808 22243
rect 738 22170 808 22187
rect 1258 22243 1328 22260
rect 1258 22187 1265 22243
rect 1321 22187 1328 22243
rect 1258 22170 1328 22187
rect -122 22007 128 22020
rect -122 21763 -119 22007
rect 125 21763 128 22007
rect -122 21750 128 21763
rect -1872 21517 -1835 21573
rect -1779 21517 -1712 21573
rect -1872 21393 -1712 21517
rect -1322 21573 -1252 21590
rect -1322 21517 -1315 21573
rect -1259 21517 -1252 21573
rect -1322 21500 -1252 21517
rect -812 21573 -742 21590
rect -812 21517 -805 21573
rect -749 21517 -742 21573
rect -812 21500 -742 21517
rect -292 21573 -222 21590
rect -292 21517 -285 21573
rect -229 21517 -222 21573
rect -292 21500 -222 21517
rect 218 21573 288 21590
rect 218 21517 225 21573
rect 281 21517 288 21573
rect 218 21500 288 21517
rect 738 21573 808 21590
rect 738 21517 745 21573
rect 801 21517 808 21573
rect 738 21500 808 21517
rect 1258 21573 1328 21590
rect 1258 21517 1265 21573
rect 1321 21517 1328 21573
rect 1258 21500 1328 21517
rect 1708 21573 1868 24302
rect 1708 21517 1775 21573
rect 1831 21517 1868 21573
rect -1872 21337 -1835 21393
rect -1779 21337 -1712 21393
rect -1872 21320 -1712 21337
rect -1322 21393 -1252 21410
rect -1322 21337 -1315 21393
rect -1259 21337 -1252 21393
rect -1322 21320 -1252 21337
rect -812 21393 -742 21410
rect -812 21337 -805 21393
rect -749 21337 -742 21393
rect -812 21320 -742 21337
rect -292 21393 -222 21410
rect -292 21337 -285 21393
rect -229 21337 -222 21393
rect -292 21320 -222 21337
rect 218 21393 288 21410
rect 218 21337 225 21393
rect 281 21337 288 21393
rect 218 21320 288 21337
rect 738 21393 808 21410
rect 738 21337 745 21393
rect 801 21337 808 21393
rect 738 21320 808 21337
rect 1258 21393 1328 21410
rect 1258 21337 1265 21393
rect 1321 21337 1328 21393
rect 1258 21320 1328 21337
rect 1708 21393 1868 21517
rect 1708 21337 1775 21393
rect 1831 21337 1868 21393
rect 1708 21320 1868 21337
rect 1988 23221 2388 23370
rect 1988 23169 2037 23221
rect 2089 23169 2287 23221
rect 2339 23169 2388 23221
rect 1988 22111 2388 23169
rect 2948 23083 3078 29637
rect 2948 23027 2985 23083
rect 3041 23027 3078 23083
rect 2948 22923 3078 23027
rect 2948 22867 2985 22923
rect 3041 22867 3078 22923
rect 2948 22840 3078 22867
rect 1988 22059 2037 22111
rect 2089 22059 2287 22111
rect 2339 22059 2388 22111
rect 1988 21701 2388 22059
rect 1988 21649 2037 21701
rect 2089 21649 2287 21701
rect 2339 21649 2388 21701
rect -1582 20903 -1512 20920
rect -1582 20847 -1575 20903
rect -1519 20847 -1512 20903
rect -1582 20830 -1512 20847
rect -1072 20903 -1002 20920
rect -1072 20847 -1065 20903
rect -1009 20847 -1002 20903
rect -1072 20830 -1002 20847
rect -552 20903 -482 20920
rect -552 20847 -545 20903
rect -489 20847 -482 20903
rect -552 20830 -482 20847
rect -32 20903 38 20920
rect -32 20847 -25 20903
rect 31 20847 38 20903
rect -32 20830 38 20847
rect 478 20903 548 20920
rect 478 20847 485 20903
rect 541 20847 548 20903
rect 478 20830 548 20847
rect 998 20903 1068 20920
rect 998 20847 1005 20903
rect 1061 20847 1068 20903
rect 998 20830 1068 20847
rect 1508 20903 1578 20920
rect 1508 20847 1515 20903
rect 1571 20847 1578 20903
rect 1508 20830 1578 20847
rect -1582 20723 -1512 20740
rect -1582 20667 -1575 20723
rect -1519 20667 -1512 20723
rect -1582 20650 -1512 20667
rect -1072 20723 -1002 20740
rect -1072 20667 -1065 20723
rect -1009 20667 -1002 20723
rect -1072 20650 -1002 20667
rect -552 20723 -482 20740
rect -552 20667 -545 20723
rect -489 20667 -482 20723
rect -552 20650 -482 20667
rect -32 20723 38 20740
rect -32 20667 -25 20723
rect 31 20667 38 20723
rect -32 20650 38 20667
rect 478 20723 548 20740
rect 478 20667 485 20723
rect 541 20667 548 20723
rect 478 20650 548 20667
rect 998 20723 1068 20740
rect 998 20667 1005 20723
rect 1061 20667 1068 20723
rect 998 20650 1068 20667
rect 1508 20723 1578 20740
rect 1508 20667 1515 20723
rect 1571 20667 1578 20723
rect 1508 20650 1578 20667
rect -2412 20539 -2363 20591
rect -2311 20539 -2113 20591
rect -2061 20539 -2012 20591
rect -2412 20370 -2012 20539
rect 1988 20591 2388 21649
rect 2638 21680 2878 21690
rect 2638 21430 2878 21440
rect 2968 21680 3208 21690
rect 2968 21430 3208 21440
rect 1988 20539 2037 20591
rect 2089 20539 2287 20591
rect 2339 20539 2388 20591
rect -122 20477 128 20490
rect -2410 20170 -330 20370
rect -122 20233 -119 20477
rect 125 20233 128 20477
rect 1988 20370 2388 20539
rect -122 20220 128 20233
rect -3220 19640 -3060 19650
rect -3220 19470 -3060 19480
rect -2160 19640 -2000 19650
rect -2160 19470 -2000 19480
rect -700 19640 -540 19650
rect -700 19470 -540 19480
rect -1740 19250 -1720 19320
rect -1650 19250 -1500 19320
rect -1430 19250 -1410 19320
rect -3220 19060 -3060 19070
rect -3220 18890 -3060 18900
rect -2160 19060 -2000 19070
rect -2160 18890 -2000 18900
rect -1740 18730 -1410 19250
rect -700 19060 -540 19070
rect -700 18890 -540 18900
rect -480 18830 -330 20170
rect 330 20170 2390 20370
rect 330 18830 480 20170
rect 520 19640 680 19650
rect 520 19470 680 19480
rect 2000 19640 2160 19650
rect 2000 19470 2160 19480
rect 3000 19640 3160 19650
rect 3000 19470 3160 19480
rect 1440 19320 1790 19330
rect 1440 19250 1460 19320
rect 1530 19250 1700 19320
rect 1770 19250 1790 19320
rect 520 19060 680 19070
rect 520 18890 680 18900
rect -1740 18660 -1720 18730
rect -1650 18660 -1500 18730
rect -1430 18660 -1410 18730
rect -1740 17470 -1410 18660
rect -580 18570 -360 18830
rect -580 18500 -560 18570
rect -490 18500 -450 18570
rect -380 18500 -360 18570
rect -580 18000 -360 18500
rect -580 17930 -560 18000
rect -490 17930 -450 18000
rect -380 17930 -360 18000
rect -840 17680 -620 17690
rect -840 17520 -620 17530
rect -1740 17400 -1720 17470
rect -1650 17400 -1510 17470
rect -1440 17400 -1410 17470
rect -1740 17380 -1410 17400
rect -1740 17310 -1720 17380
rect -1650 17310 -1510 17380
rect -1440 17310 -1410 17380
rect -3200 17120 -3020 17130
rect -3200 16980 -3020 16990
rect -2060 17120 -1880 17130
rect -2060 16980 -1880 16990
rect -1740 16950 -1410 17310
rect -580 17250 -360 17930
rect 360 18570 580 18830
rect 360 18500 380 18570
rect 450 18500 490 18570
rect 560 18500 580 18570
rect 360 18010 580 18500
rect 360 17940 380 18010
rect 450 17940 490 18010
rect 560 17940 580 18010
rect -320 17680 -100 17690
rect -320 17520 -100 17530
rect 100 17680 320 17690
rect 100 17520 320 17530
rect -580 17180 -560 17250
rect -490 17180 -450 17250
rect -380 17180 -360 17250
rect -1080 17130 -900 17140
rect -1080 16990 -900 17000
rect -1740 16880 -1720 16950
rect -1650 16880 -1500 16950
rect -1430 16880 -1410 16950
rect -1740 16870 -1410 16880
rect -580 16800 -360 17180
rect 360 17250 580 17940
rect 1440 18730 1790 19250
rect 2000 19060 2160 19070
rect 2000 18890 2160 18900
rect 3000 19060 3160 19070
rect 3000 18890 3160 18900
rect 1440 18660 1460 18730
rect 1530 18660 1700 18730
rect 1770 18660 1790 18730
rect 650 17680 870 17690
rect 650 17520 870 17530
rect 360 17180 380 17250
rect 450 17180 490 17250
rect 560 17180 580 17250
rect -310 17130 -130 17140
rect -310 16990 -130 17000
rect 130 17130 310 17140
rect 130 16990 310 17000
rect -580 16730 -560 16800
rect -490 16730 -450 16800
rect -380 16730 -360 16800
rect -580 16660 -360 16730
rect 360 16800 580 17180
rect 1440 17490 1790 18660
rect 1440 17420 1460 17490
rect 1530 17420 1700 17490
rect 1770 17420 1790 17490
rect 1440 17400 1790 17420
rect 1440 17330 1460 17400
rect 1530 17330 1700 17400
rect 1770 17330 1790 17400
rect 850 17120 1030 17130
rect 850 16980 1030 16990
rect 1440 16950 1790 17330
rect 1920 17130 2100 17140
rect 1920 16990 2100 17000
rect 2920 17130 3100 17140
rect 2920 16990 3100 17000
rect 1440 16880 1460 16950
rect 1530 16880 1700 16950
rect 1770 16880 1790 16950
rect 1440 16850 1790 16880
rect 360 16730 380 16800
rect 450 16730 490 16800
rect 560 16730 580 16800
rect 360 16670 580 16730
rect -3240 15220 -3120 15230
rect -3240 15090 -3120 15100
rect 3130 15220 3250 15230
rect 3130 15090 3250 15100
rect -3240 12220 -3120 12230
rect -3240 12090 -3120 12100
rect 3130 12220 3250 12230
rect 3130 12090 3250 12100
rect -3240 9220 -3120 9230
rect -3240 9090 -3120 9100
rect 3130 9220 3250 9230
rect 3130 9090 3250 9100
rect -3240 6220 -3120 6230
rect -3240 6090 -3120 6100
rect 3130 6220 3250 6230
rect 3130 6090 3250 6100
rect -3240 3220 -3120 3230
rect -3240 3090 -3120 3100
rect 3130 3220 3250 3230
rect 3130 3090 3250 3100
rect 1690 1900 2860 1910
rect -2860 1890 -1690 1900
rect -2860 1470 -1690 1480
rect -1350 1890 -180 1900
rect -1350 1470 -180 1480
rect 170 1890 1340 1900
rect 1690 1480 2860 1490
rect 170 1470 1340 1480
<< via2 >>
rect -615 31157 -399 31373
rect 435 31157 651 31373
rect -3185 30911 -3129 30913
rect -3185 30859 -3183 30911
rect -3183 30859 -3131 30911
rect -3131 30859 -3129 30911
rect -3185 30857 -3129 30859
rect -2865 30911 -2809 30913
rect -2865 30859 -2863 30911
rect -2863 30859 -2811 30911
rect -2811 30859 -2809 30911
rect -2865 30857 -2809 30859
rect -2555 30911 -2499 30913
rect -2555 30859 -2553 30911
rect -2553 30859 -2501 30911
rect -2501 30859 -2499 30911
rect -2555 30857 -2499 30859
rect -2235 30911 -2179 30913
rect -2235 30859 -2233 30911
rect -2233 30859 -2181 30911
rect -2181 30859 -2179 30911
rect -2235 30857 -2179 30859
rect -1925 30911 -1869 30913
rect -1925 30859 -1923 30911
rect -1923 30859 -1871 30911
rect -1871 30859 -1869 30911
rect -1925 30857 -1869 30859
rect -1605 30911 -1549 30913
rect -1605 30859 -1603 30911
rect -1603 30859 -1551 30911
rect -1551 30859 -1549 30911
rect -1605 30857 -1549 30859
rect -1285 30911 -1229 30913
rect -1285 30859 -1283 30911
rect -1283 30859 -1231 30911
rect -1231 30859 -1229 30911
rect -1285 30857 -1229 30859
rect -975 30911 -919 30913
rect -975 30859 -973 30911
rect -973 30859 -921 30911
rect -921 30859 -919 30911
rect -975 30857 -919 30859
rect -655 30911 -599 30913
rect -655 30859 -653 30911
rect -653 30859 -601 30911
rect -601 30859 -599 30911
rect -655 30857 -599 30859
rect -335 30911 -279 30913
rect -335 30859 -333 30911
rect -333 30859 -281 30911
rect -281 30859 -279 30911
rect -335 30857 -279 30859
rect -25 30911 31 30913
rect -25 30859 -23 30911
rect -23 30859 29 30911
rect 29 30859 31 30911
rect -25 30857 31 30859
rect 295 30911 351 30913
rect 295 30859 297 30911
rect 297 30859 349 30911
rect 349 30859 351 30911
rect 295 30857 351 30859
rect 605 30911 661 30913
rect 605 30859 607 30911
rect 607 30859 659 30911
rect 659 30859 661 30911
rect 605 30857 661 30859
rect 925 30911 981 30913
rect 925 30859 927 30911
rect 927 30859 979 30911
rect 979 30859 981 30911
rect 925 30857 981 30859
rect 1245 30911 1301 30913
rect 1245 30859 1247 30911
rect 1247 30859 1299 30911
rect 1299 30859 1301 30911
rect 1245 30857 1301 30859
rect 1555 30911 1611 30913
rect 1555 30859 1557 30911
rect 1557 30859 1609 30911
rect 1609 30859 1611 30911
rect 1555 30857 1611 30859
rect 1875 30911 1931 30913
rect 1875 30859 1877 30911
rect 1877 30859 1929 30911
rect 1929 30859 1931 30911
rect 1875 30857 1931 30859
rect 2185 30911 2241 30913
rect 2185 30859 2187 30911
rect 2187 30859 2239 30911
rect 2239 30859 2241 30911
rect 2185 30857 2241 30859
rect 2505 30911 2561 30913
rect 2505 30859 2507 30911
rect 2507 30859 2559 30911
rect 2559 30859 2561 30911
rect 2505 30857 2561 30859
rect 2825 30911 2881 30913
rect 2825 30859 2827 30911
rect 2827 30859 2879 30911
rect 2879 30859 2881 30911
rect 2825 30857 2881 30859
rect 3135 30911 3191 30913
rect 3135 30859 3137 30911
rect 3137 30859 3189 30911
rect 3189 30859 3191 30911
rect 3135 30857 3191 30859
rect -7912 30560 -7852 30620
rect -7792 30560 -7732 30620
rect -3185 30671 -3129 30673
rect -3185 30619 -3183 30671
rect -3183 30619 -3131 30671
rect -3131 30619 -3129 30671
rect -3185 30617 -3129 30619
rect -2865 30671 -2809 30673
rect -2865 30619 -2863 30671
rect -2863 30619 -2811 30671
rect -2811 30619 -2809 30671
rect -2865 30617 -2809 30619
rect -2555 30671 -2499 30673
rect -2555 30619 -2553 30671
rect -2553 30619 -2501 30671
rect -2501 30619 -2499 30671
rect -2555 30617 -2499 30619
rect -2235 30671 -2179 30673
rect -2235 30619 -2233 30671
rect -2233 30619 -2181 30671
rect -2181 30619 -2179 30671
rect -2235 30617 -2179 30619
rect -1925 30671 -1869 30673
rect -1925 30619 -1923 30671
rect -1923 30619 -1871 30671
rect -1871 30619 -1869 30671
rect -1925 30617 -1869 30619
rect -1605 30671 -1549 30673
rect -1605 30619 -1603 30671
rect -1603 30619 -1551 30671
rect -1551 30619 -1549 30671
rect -1605 30617 -1549 30619
rect -1285 30671 -1229 30673
rect -1285 30619 -1283 30671
rect -1283 30619 -1231 30671
rect -1231 30619 -1229 30671
rect -1285 30617 -1229 30619
rect -975 30671 -919 30673
rect -975 30619 -973 30671
rect -973 30619 -921 30671
rect -921 30619 -919 30671
rect -975 30617 -919 30619
rect -655 30671 -599 30673
rect -655 30619 -653 30671
rect -653 30619 -601 30671
rect -601 30619 -599 30671
rect -655 30617 -599 30619
rect -335 30671 -279 30673
rect -335 30619 -333 30671
rect -333 30619 -281 30671
rect -281 30619 -279 30671
rect -335 30617 -279 30619
rect -25 30671 31 30673
rect -25 30619 -23 30671
rect -23 30619 29 30671
rect 29 30619 31 30671
rect -25 30617 31 30619
rect 295 30671 351 30673
rect 295 30619 297 30671
rect 297 30619 349 30671
rect 349 30619 351 30671
rect 295 30617 351 30619
rect 605 30671 661 30673
rect 605 30619 607 30671
rect 607 30619 659 30671
rect 659 30619 661 30671
rect 605 30617 661 30619
rect 925 30671 981 30673
rect 925 30619 927 30671
rect 927 30619 979 30671
rect 979 30619 981 30671
rect 925 30617 981 30619
rect 1245 30671 1301 30673
rect 1245 30619 1247 30671
rect 1247 30619 1299 30671
rect 1299 30619 1301 30671
rect 1245 30617 1301 30619
rect 1555 30671 1611 30673
rect 1555 30619 1557 30671
rect 1557 30619 1609 30671
rect 1609 30619 1611 30671
rect 1555 30617 1611 30619
rect 1875 30671 1931 30673
rect 1875 30619 1877 30671
rect 1877 30619 1929 30671
rect 1929 30619 1931 30671
rect 1875 30617 1931 30619
rect 2185 30671 2241 30673
rect 2185 30619 2187 30671
rect 2187 30619 2239 30671
rect 2239 30619 2241 30671
rect 2185 30617 2241 30619
rect 2505 30671 2561 30673
rect 2505 30619 2507 30671
rect 2507 30619 2559 30671
rect 2559 30619 2561 30671
rect 2505 30617 2561 30619
rect 2825 30671 2881 30673
rect 2825 30619 2827 30671
rect 2827 30619 2879 30671
rect 2879 30619 2881 30671
rect 2825 30617 2881 30619
rect 3135 30671 3191 30673
rect 3135 30619 3137 30671
rect 3137 30619 3189 30671
rect 3189 30619 3191 30671
rect 3135 30617 3191 30619
rect 8000 30616 8056 30618
rect 8000 30564 8002 30616
rect 8002 30564 8054 30616
rect 8054 30564 8056 30616
rect 8000 30562 8056 30564
rect 8110 30616 8166 30618
rect 8110 30564 8112 30616
rect 8112 30564 8164 30616
rect 8164 30564 8166 30616
rect 8110 30562 8166 30564
rect -3025 30301 -2969 30303
rect -3025 30249 -3023 30301
rect -3023 30249 -2971 30301
rect -2971 30249 -2969 30301
rect -3025 30247 -2969 30249
rect -2715 30301 -2659 30303
rect -2715 30249 -2713 30301
rect -2713 30249 -2661 30301
rect -2661 30249 -2659 30301
rect -2715 30247 -2659 30249
rect -2395 30301 -2339 30303
rect -2395 30249 -2393 30301
rect -2393 30249 -2341 30301
rect -2341 30249 -2339 30301
rect -2395 30247 -2339 30249
rect -2075 30301 -2019 30303
rect -2075 30249 -2073 30301
rect -2073 30249 -2021 30301
rect -2021 30249 -2019 30301
rect -2075 30247 -2019 30249
rect -1765 30301 -1709 30303
rect -1765 30249 -1763 30301
rect -1763 30249 -1711 30301
rect -1711 30249 -1709 30301
rect -1765 30247 -1709 30249
rect -1445 30301 -1389 30303
rect -1445 30249 -1443 30301
rect -1443 30249 -1391 30301
rect -1391 30249 -1389 30301
rect -1445 30247 -1389 30249
rect -1135 30301 -1079 30303
rect -1135 30249 -1133 30301
rect -1133 30249 -1081 30301
rect -1081 30249 -1079 30301
rect -1135 30247 -1079 30249
rect -815 30301 -759 30303
rect -815 30249 -813 30301
rect -813 30249 -761 30301
rect -761 30249 -759 30301
rect -815 30247 -759 30249
rect -495 30301 -439 30303
rect -495 30249 -493 30301
rect -493 30249 -441 30301
rect -441 30249 -439 30301
rect -495 30247 -439 30249
rect -185 30301 -129 30303
rect -185 30249 -183 30301
rect -183 30249 -131 30301
rect -131 30249 -129 30301
rect -185 30247 -129 30249
rect 135 30301 191 30303
rect 135 30249 137 30301
rect 137 30249 189 30301
rect 189 30249 191 30301
rect 135 30247 191 30249
rect 455 30301 511 30303
rect 455 30249 457 30301
rect 457 30249 509 30301
rect 509 30249 511 30301
rect 455 30247 511 30249
rect 765 30301 821 30303
rect 765 30249 767 30301
rect 767 30249 819 30301
rect 819 30249 821 30301
rect 765 30247 821 30249
rect 1085 30301 1141 30303
rect 1085 30249 1087 30301
rect 1087 30249 1139 30301
rect 1139 30249 1141 30301
rect 1085 30247 1141 30249
rect 1395 30301 1451 30303
rect 1395 30249 1397 30301
rect 1397 30249 1449 30301
rect 1449 30249 1451 30301
rect 1395 30247 1451 30249
rect 1715 30301 1771 30303
rect 1715 30249 1717 30301
rect 1717 30249 1769 30301
rect 1769 30249 1771 30301
rect 1715 30247 1771 30249
rect 2035 30301 2091 30303
rect 2035 30249 2037 30301
rect 2037 30249 2089 30301
rect 2089 30249 2091 30301
rect 2035 30247 2091 30249
rect 2345 30301 2401 30303
rect 2345 30249 2347 30301
rect 2347 30249 2399 30301
rect 2399 30249 2401 30301
rect 2345 30247 2401 30249
rect 2665 30301 2721 30303
rect 2665 30249 2667 30301
rect 2667 30249 2719 30301
rect 2719 30249 2721 30301
rect 2665 30247 2721 30249
rect 2985 30301 3041 30303
rect 2985 30249 2987 30301
rect 2987 30249 3039 30301
rect 3039 30249 3041 30301
rect 2985 30247 3041 30249
rect -3025 30061 -2969 30063
rect -3025 30009 -3023 30061
rect -3023 30009 -2971 30061
rect -2971 30009 -2969 30061
rect -3025 30007 -2969 30009
rect -2715 30061 -2659 30063
rect -2715 30009 -2713 30061
rect -2713 30009 -2661 30061
rect -2661 30009 -2659 30061
rect -2715 30007 -2659 30009
rect -2395 30061 -2339 30063
rect -2395 30009 -2393 30061
rect -2393 30009 -2341 30061
rect -2341 30009 -2339 30061
rect -2395 30007 -2339 30009
rect -2075 30061 -2019 30063
rect -2075 30009 -2073 30061
rect -2073 30009 -2021 30061
rect -2021 30009 -2019 30061
rect -2075 30007 -2019 30009
rect -1765 30061 -1709 30063
rect -1765 30009 -1763 30061
rect -1763 30009 -1711 30061
rect -1711 30009 -1709 30061
rect -1765 30007 -1709 30009
rect -1445 30061 -1389 30063
rect -1445 30009 -1443 30061
rect -1443 30009 -1391 30061
rect -1391 30009 -1389 30061
rect -1445 30007 -1389 30009
rect -1135 30061 -1079 30063
rect -1135 30009 -1133 30061
rect -1133 30009 -1081 30061
rect -1081 30009 -1079 30061
rect -1135 30007 -1079 30009
rect -815 30061 -759 30063
rect -815 30009 -813 30061
rect -813 30009 -761 30061
rect -761 30009 -759 30061
rect -815 30007 -759 30009
rect -495 30061 -439 30063
rect -495 30009 -493 30061
rect -493 30009 -441 30061
rect -441 30009 -439 30061
rect -495 30007 -439 30009
rect -185 30061 -129 30063
rect -185 30009 -183 30061
rect -183 30009 -131 30061
rect -131 30009 -129 30061
rect -185 30007 -129 30009
rect 135 30061 191 30063
rect 135 30009 137 30061
rect 137 30009 189 30061
rect 189 30009 191 30061
rect 135 30007 191 30009
rect 455 30061 511 30063
rect 455 30009 457 30061
rect 457 30009 509 30061
rect 509 30009 511 30061
rect 455 30007 511 30009
rect 765 30061 821 30063
rect 765 30009 767 30061
rect 767 30009 819 30061
rect 819 30009 821 30061
rect 765 30007 821 30009
rect 1085 30061 1141 30063
rect 1085 30009 1087 30061
rect 1087 30009 1139 30061
rect 1139 30009 1141 30061
rect 1085 30007 1141 30009
rect 1395 30061 1451 30063
rect 1395 30009 1397 30061
rect 1397 30009 1449 30061
rect 1449 30009 1451 30061
rect 1395 30007 1451 30009
rect 1715 30061 1771 30063
rect 1715 30009 1717 30061
rect 1717 30009 1769 30061
rect 1769 30009 1771 30061
rect 1715 30007 1771 30009
rect 2035 30061 2091 30063
rect 2035 30009 2037 30061
rect 2037 30009 2089 30061
rect 2089 30009 2091 30061
rect 2035 30007 2091 30009
rect 2345 30061 2401 30063
rect 2345 30009 2347 30061
rect 2347 30009 2399 30061
rect 2399 30009 2401 30061
rect 2345 30007 2401 30009
rect 2665 30061 2721 30063
rect 2665 30009 2667 30061
rect 2667 30009 2719 30061
rect 2719 30009 2721 30061
rect 2665 30007 2721 30009
rect 2985 30061 3041 30063
rect 2985 30009 2987 30061
rect 2987 30009 3039 30061
rect 3039 30009 3041 30061
rect 2985 30007 3041 30009
rect -3025 29637 -2969 29693
rect -615 29517 -399 29733
rect 435 29517 651 29733
rect -1685 29241 -1629 29243
rect -1685 29189 -1683 29241
rect -1683 29189 -1631 29241
rect -1631 29189 -1629 29241
rect -1685 29187 -1629 29189
rect -1365 29241 -1309 29243
rect -1365 29189 -1363 29241
rect -1363 29189 -1311 29241
rect -1311 29189 -1309 29241
rect -1365 29187 -1309 29189
rect -1055 29241 -999 29243
rect -1055 29189 -1053 29241
rect -1053 29189 -1001 29241
rect -1001 29189 -999 29241
rect -1055 29187 -999 29189
rect -735 29241 -679 29243
rect -735 29189 -733 29241
rect -733 29189 -681 29241
rect -681 29189 -679 29241
rect -735 29187 -679 29189
rect -415 29241 -359 29243
rect -415 29189 -413 29241
rect -413 29189 -361 29241
rect -361 29189 -359 29241
rect -415 29187 -359 29189
rect -105 29241 -49 29243
rect -105 29189 -103 29241
rect -103 29189 -51 29241
rect -51 29189 -49 29241
rect -105 29187 -49 29189
rect 215 29241 271 29243
rect 215 29189 217 29241
rect 217 29189 269 29241
rect 269 29189 271 29241
rect 215 29187 271 29189
rect 535 29241 591 29243
rect 535 29189 537 29241
rect 537 29189 589 29241
rect 589 29189 591 29241
rect 535 29187 591 29189
rect 845 29241 901 29243
rect 845 29189 847 29241
rect 847 29189 899 29241
rect 899 29189 901 29241
rect 845 29187 901 29189
rect 1165 29241 1221 29243
rect 1165 29189 1167 29241
rect 1167 29189 1219 29241
rect 1219 29189 1221 29241
rect 1165 29187 1221 29189
rect 1475 29241 1531 29243
rect 1475 29189 1477 29241
rect 1477 29189 1529 29241
rect 1529 29189 1531 29241
rect 1475 29187 1531 29189
rect -1685 29031 -1629 29033
rect -1685 28979 -1683 29031
rect -1683 28979 -1631 29031
rect -1631 28979 -1629 29031
rect -1685 28977 -1629 28979
rect -1365 29031 -1309 29033
rect -1365 28979 -1363 29031
rect -1363 28979 -1311 29031
rect -1311 28979 -1309 29031
rect -1365 28977 -1309 28979
rect -1055 29031 -999 29033
rect -1055 28979 -1053 29031
rect -1053 28979 -1001 29031
rect -1001 28979 -999 29031
rect -1055 28977 -999 28979
rect -735 29031 -679 29033
rect -735 28979 -733 29031
rect -733 28979 -681 29031
rect -681 28979 -679 29031
rect -735 28977 -679 28979
rect -415 29031 -359 29033
rect -415 28979 -413 29031
rect -413 28979 -361 29031
rect -361 28979 -359 29031
rect -415 28977 -359 28979
rect -105 29031 -49 29033
rect -105 28979 -103 29031
rect -103 28979 -51 29031
rect -51 28979 -49 29031
rect -105 28977 -49 28979
rect 215 29031 271 29033
rect 215 28979 217 29031
rect 217 28979 269 29031
rect 269 28979 271 29031
rect 215 28977 271 28979
rect 535 29031 591 29033
rect 535 28979 537 29031
rect 537 28979 589 29031
rect 589 28979 591 29031
rect 535 28977 591 28979
rect 845 29031 901 29033
rect 845 28979 847 29031
rect 847 28979 899 29031
rect 899 28979 901 29031
rect 845 28977 901 28979
rect 1165 29031 1221 29033
rect 1165 28979 1167 29031
rect 1167 28979 1219 29031
rect 1219 28979 1221 29031
rect 1165 28977 1221 28979
rect 1475 29031 1531 29033
rect 1475 28979 1477 29031
rect 1477 28979 1529 29031
rect 1529 28979 1531 29031
rect 1475 28977 1531 28979
rect -2060 28532 -2004 28588
rect -1525 28601 -1469 28603
rect -1525 28549 -1523 28601
rect -1523 28549 -1471 28601
rect -1471 28549 -1469 28601
rect -1525 28547 -1469 28549
rect -1205 28601 -1149 28603
rect -1205 28549 -1203 28601
rect -1203 28549 -1151 28601
rect -1151 28549 -1149 28601
rect -1205 28547 -1149 28549
rect -895 28601 -839 28603
rect -895 28549 -893 28601
rect -893 28549 -841 28601
rect -841 28549 -839 28601
rect -895 28547 -839 28549
rect -575 28601 -519 28603
rect -575 28549 -573 28601
rect -573 28549 -521 28601
rect -521 28549 -519 28601
rect -575 28547 -519 28549
rect -255 28601 -199 28603
rect -255 28549 -253 28601
rect -253 28549 -201 28601
rect -201 28549 -199 28601
rect -255 28547 -199 28549
rect 55 28601 111 28603
rect 55 28549 57 28601
rect 57 28549 109 28601
rect 109 28549 111 28601
rect 55 28547 111 28549
rect 375 28601 431 28603
rect 375 28549 377 28601
rect 377 28549 429 28601
rect 429 28549 431 28601
rect 375 28547 431 28549
rect 685 28601 741 28603
rect 685 28549 687 28601
rect 687 28549 739 28601
rect 739 28549 741 28601
rect 685 28547 741 28549
rect 1005 28601 1061 28603
rect 1005 28549 1007 28601
rect 1007 28549 1059 28601
rect 1059 28549 1061 28601
rect 1005 28547 1061 28549
rect 1325 28601 1381 28603
rect 1325 28549 1327 28601
rect 1327 28549 1379 28601
rect 1379 28549 1381 28601
rect 1325 28547 1381 28549
rect 1635 28601 1691 28603
rect 1635 28549 1637 28601
rect 1637 28549 1689 28601
rect 1689 28549 1691 28601
rect 1635 28547 1691 28549
rect 2000 28532 2056 28588
rect -2060 28352 -2004 28408
rect -1525 28391 -1469 28393
rect -1525 28339 -1523 28391
rect -1523 28339 -1471 28391
rect -1471 28339 -1469 28391
rect -1525 28337 -1469 28339
rect -1205 28391 -1149 28393
rect -1205 28339 -1203 28391
rect -1203 28339 -1151 28391
rect -1151 28339 -1149 28391
rect -1205 28337 -1149 28339
rect -895 28391 -839 28393
rect -895 28339 -893 28391
rect -893 28339 -841 28391
rect -841 28339 -839 28391
rect -895 28337 -839 28339
rect -575 28391 -519 28393
rect -575 28339 -573 28391
rect -573 28339 -521 28391
rect -521 28339 -519 28391
rect -575 28337 -519 28339
rect -255 28391 -199 28393
rect -255 28339 -253 28391
rect -253 28339 -201 28391
rect -201 28339 -199 28391
rect -255 28337 -199 28339
rect 55 28391 111 28393
rect 55 28339 57 28391
rect 57 28339 109 28391
rect 109 28339 111 28391
rect 55 28337 111 28339
rect 375 28391 431 28393
rect 375 28339 377 28391
rect 377 28339 429 28391
rect 429 28339 431 28391
rect 375 28337 431 28339
rect 685 28391 741 28393
rect 685 28339 687 28391
rect 687 28339 739 28391
rect 739 28339 741 28391
rect 685 28337 741 28339
rect 1005 28391 1061 28393
rect 1005 28339 1007 28391
rect 1007 28339 1059 28391
rect 1059 28339 1061 28391
rect 1005 28337 1061 28339
rect 1325 28391 1381 28393
rect 1325 28339 1327 28391
rect 1327 28339 1379 28391
rect 1379 28339 1381 28391
rect 1325 28337 1381 28339
rect 1635 28391 1691 28393
rect 1635 28339 1637 28391
rect 1637 28339 1689 28391
rect 1689 28339 1691 28391
rect 1635 28337 1691 28339
rect 2000 28352 2056 28408
rect -850 27912 -634 28128
rect 650 27912 866 28128
rect -1685 27691 -1629 27693
rect -1685 27639 -1683 27691
rect -1683 27639 -1631 27691
rect -1631 27639 -1629 27691
rect -1685 27637 -1629 27639
rect -1365 27691 -1309 27693
rect -1365 27639 -1363 27691
rect -1363 27639 -1311 27691
rect -1311 27639 -1309 27691
rect -1365 27637 -1309 27639
rect -1055 27691 -999 27693
rect -1055 27639 -1053 27691
rect -1053 27639 -1001 27691
rect -1001 27639 -999 27691
rect -1055 27637 -999 27639
rect -735 27691 -679 27693
rect -735 27639 -733 27691
rect -733 27639 -681 27691
rect -681 27639 -679 27691
rect -735 27637 -679 27639
rect -415 27691 -359 27693
rect -415 27639 -413 27691
rect -413 27639 -361 27691
rect -361 27639 -359 27691
rect -415 27637 -359 27639
rect -105 27691 -49 27693
rect -105 27639 -103 27691
rect -103 27639 -51 27691
rect -51 27639 -49 27691
rect -105 27637 -49 27639
rect 215 27691 271 27693
rect 215 27639 217 27691
rect 217 27639 269 27691
rect 269 27639 271 27691
rect 215 27637 271 27639
rect 525 27691 581 27693
rect 525 27639 527 27691
rect 527 27639 579 27691
rect 579 27639 581 27691
rect 525 27637 581 27639
rect 845 27691 901 27693
rect 845 27639 847 27691
rect 847 27639 899 27691
rect 899 27639 901 27691
rect 845 27637 901 27639
rect 1165 27691 1221 27693
rect 1165 27639 1167 27691
rect 1167 27639 1219 27691
rect 1219 27639 1221 27691
rect 1165 27637 1221 27639
rect 1475 27691 1531 27693
rect 1475 27639 1477 27691
rect 1477 27639 1529 27691
rect 1529 27639 1531 27691
rect 1475 27637 1531 27639
rect -1685 27481 -1629 27483
rect -1685 27429 -1683 27481
rect -1683 27429 -1631 27481
rect -1631 27429 -1629 27481
rect -1685 27427 -1629 27429
rect -1365 27481 -1309 27483
rect -1365 27429 -1363 27481
rect -1363 27429 -1311 27481
rect -1311 27429 -1309 27481
rect -1365 27427 -1309 27429
rect -1055 27481 -999 27483
rect -1055 27429 -1053 27481
rect -1053 27429 -1001 27481
rect -1001 27429 -999 27481
rect -1055 27427 -999 27429
rect -735 27481 -679 27483
rect -735 27429 -733 27481
rect -733 27429 -681 27481
rect -681 27429 -679 27481
rect -735 27427 -679 27429
rect -415 27481 -359 27483
rect -415 27429 -413 27481
rect -413 27429 -361 27481
rect -361 27429 -359 27481
rect -415 27427 -359 27429
rect -105 27481 -49 27483
rect -105 27429 -103 27481
rect -103 27429 -51 27481
rect -51 27429 -49 27481
rect -105 27427 -49 27429
rect 215 27481 271 27483
rect 215 27429 217 27481
rect 217 27429 269 27481
rect 269 27429 271 27481
rect 215 27427 271 27429
rect 525 27481 581 27483
rect 525 27429 527 27481
rect 527 27429 579 27481
rect 579 27429 581 27481
rect 525 27427 581 27429
rect 845 27481 901 27483
rect 845 27429 847 27481
rect 847 27429 899 27481
rect 899 27429 901 27481
rect 845 27427 901 27429
rect 1165 27481 1221 27483
rect 1165 27429 1167 27481
rect 1167 27429 1219 27481
rect 1219 27429 1221 27481
rect 1165 27427 1221 27429
rect 1475 27481 1531 27483
rect 1475 27429 1477 27481
rect 1477 27429 1529 27481
rect 1529 27429 1531 27481
rect 1475 27427 1531 27429
rect -1525 27061 -1469 27063
rect -1525 27009 -1523 27061
rect -1523 27009 -1471 27061
rect -1471 27009 -1469 27061
rect -1525 27007 -1469 27009
rect -1205 27061 -1149 27063
rect -1205 27009 -1203 27061
rect -1203 27009 -1151 27061
rect -1151 27009 -1149 27061
rect -1205 27007 -1149 27009
rect -1525 26851 -1469 26853
rect -1525 26799 -1523 26851
rect -1523 26799 -1471 26851
rect -1471 26799 -1469 26851
rect -1525 26797 -1469 26799
rect -895 27061 -839 27063
rect -895 27009 -893 27061
rect -893 27009 -841 27061
rect -841 27009 -839 27061
rect -895 27007 -839 27009
rect -575 27061 -519 27063
rect -575 27009 -573 27061
rect -573 27009 -521 27061
rect -521 27009 -519 27061
rect -575 27007 -519 27009
rect -265 27061 -209 27063
rect -265 27009 -263 27061
rect -263 27009 -211 27061
rect -211 27009 -209 27061
rect -265 27007 -209 27009
rect 55 27061 111 27063
rect 55 27009 57 27061
rect 57 27009 109 27061
rect 109 27009 111 27061
rect 55 27007 111 27009
rect 375 27061 431 27063
rect 375 27009 377 27061
rect 377 27009 429 27061
rect 429 27009 431 27061
rect 375 27007 431 27009
rect 685 27061 741 27063
rect 685 27009 687 27061
rect 687 27009 739 27061
rect 739 27009 741 27061
rect 685 27007 741 27009
rect 1005 27061 1061 27063
rect 1005 27009 1007 27061
rect 1007 27009 1059 27061
rect 1059 27009 1061 27061
rect 1005 27007 1061 27009
rect 1315 27061 1371 27063
rect 1315 27009 1317 27061
rect 1317 27009 1369 27061
rect 1369 27009 1371 27061
rect 1315 27007 1371 27009
rect -1205 26851 -1149 26853
rect -1205 26799 -1203 26851
rect -1203 26799 -1151 26851
rect -1151 26799 -1149 26851
rect -1205 26797 -1149 26799
rect -2060 26042 -2004 26098
rect -2060 25822 -2004 25878
rect -1820 25482 -1764 25538
rect -1820 25262 -1764 25318
rect -1820 24522 -1764 24578
rect -1820 24302 -1764 24358
rect -3025 23027 -2969 23083
rect -3025 22867 -2969 22923
rect -3235 21716 -2699 21718
rect -3235 21344 -2699 21716
rect -3235 21342 -2699 21344
rect -895 26851 -839 26853
rect -895 26799 -893 26851
rect -893 26799 -841 26851
rect -841 26799 -839 26851
rect -895 26797 -839 26799
rect -575 26851 -519 26853
rect -575 26799 -573 26851
rect -573 26799 -521 26851
rect -521 26799 -519 26851
rect -575 26797 -519 26799
rect -265 26851 -209 26853
rect -265 26799 -263 26851
rect -263 26799 -211 26851
rect -211 26799 -209 26851
rect -265 26797 -209 26799
rect 55 26851 111 26853
rect 55 26799 57 26851
rect 57 26799 109 26851
rect 109 26799 111 26851
rect 55 26797 111 26799
rect 375 26851 431 26853
rect 375 26799 377 26851
rect 377 26799 429 26851
rect 429 26799 431 26851
rect 375 26797 431 26799
rect 685 26851 741 26853
rect 685 26799 687 26851
rect 687 26799 739 26851
rect 739 26799 741 26851
rect 685 26797 741 26799
rect 1005 26851 1061 26853
rect 1005 26799 1007 26851
rect 1007 26799 1059 26851
rect 1059 26799 1061 26851
rect 1005 26797 1061 26799
rect 1635 27061 1691 27063
rect 1635 27009 1637 27061
rect 1637 27009 1689 27061
rect 1689 27009 1691 27061
rect 1635 27007 1691 27009
rect 1315 26851 1371 26853
rect 1315 26799 1317 26851
rect 1317 26799 1369 26851
rect 1369 26799 1371 26851
rect 1315 26797 1371 26799
rect -585 26131 -529 26133
rect -585 26079 -583 26131
rect -583 26079 -531 26131
rect -531 26079 -529 26131
rect -585 26077 -529 26079
rect -265 26131 -209 26133
rect -265 26079 -263 26131
rect -263 26079 -211 26131
rect -211 26079 -209 26131
rect -265 26077 -209 26079
rect 45 26131 101 26133
rect 45 26079 47 26131
rect 47 26079 99 26131
rect 99 26079 101 26131
rect 45 26077 101 26079
rect 365 26131 421 26133
rect 365 26079 367 26131
rect 367 26079 419 26131
rect 419 26079 421 26131
rect 365 26077 421 26079
rect -585 25841 -529 25843
rect -585 25789 -583 25841
rect -583 25789 -531 25841
rect -531 25789 -529 25841
rect -585 25787 -529 25789
rect -265 25841 -209 25843
rect -265 25789 -263 25841
rect -263 25789 -211 25841
rect -211 25789 -209 25841
rect -265 25787 -209 25789
rect 45 25841 101 25843
rect 45 25789 47 25841
rect 47 25789 99 25841
rect 99 25789 101 25841
rect 45 25787 101 25789
rect 365 25841 421 25843
rect 365 25789 367 25841
rect 367 25789 419 25841
rect 419 25789 421 25841
rect 365 25787 421 25789
rect -425 25571 -369 25573
rect -425 25519 -423 25571
rect -423 25519 -371 25571
rect -371 25519 -369 25571
rect -425 25517 -369 25519
rect -115 25571 -59 25573
rect -115 25519 -113 25571
rect -113 25519 -61 25571
rect -61 25519 -59 25571
rect -115 25517 -59 25519
rect 205 25571 261 25573
rect 205 25519 207 25571
rect 207 25519 259 25571
rect 259 25519 261 25571
rect 205 25517 261 25519
rect 525 25571 581 25573
rect 525 25519 527 25571
rect 527 25519 579 25571
rect 579 25519 581 25571
rect 525 25517 581 25519
rect -425 25281 -369 25283
rect -425 25229 -423 25281
rect -423 25229 -371 25281
rect -371 25229 -369 25281
rect -425 25227 -369 25229
rect -115 25281 -59 25283
rect -115 25229 -113 25281
rect -113 25229 -61 25281
rect -61 25229 -59 25281
rect -115 25227 -59 25229
rect 205 25281 261 25283
rect 205 25229 207 25281
rect 207 25229 259 25281
rect 259 25229 261 25281
rect 205 25227 261 25229
rect 525 25281 581 25283
rect 525 25229 527 25281
rect 527 25229 579 25281
rect 579 25229 581 25281
rect 525 25227 581 25229
rect -110 24812 106 25028
rect -585 24611 -529 24613
rect -585 24559 -583 24611
rect -583 24559 -531 24611
rect -531 24559 -529 24611
rect -585 24557 -529 24559
rect -265 24611 -209 24613
rect -265 24559 -263 24611
rect -263 24559 -211 24611
rect -211 24559 -209 24611
rect -265 24557 -209 24559
rect 45 24611 101 24613
rect 45 24559 47 24611
rect 47 24559 99 24611
rect 99 24559 101 24611
rect 45 24557 101 24559
rect 365 24611 421 24613
rect 365 24559 367 24611
rect 367 24559 419 24611
rect 419 24559 421 24611
rect 365 24557 421 24559
rect -585 24321 -529 24323
rect -585 24269 -583 24321
rect -583 24269 -531 24321
rect -531 24269 -529 24321
rect -585 24267 -529 24269
rect -265 24321 -209 24323
rect -265 24269 -263 24321
rect -263 24269 -211 24321
rect -211 24269 -209 24321
rect -265 24267 -209 24269
rect 45 24321 101 24323
rect 45 24269 47 24321
rect 47 24269 99 24321
rect 99 24269 101 24321
rect 45 24267 101 24269
rect 365 24321 421 24323
rect 365 24269 367 24321
rect 367 24269 419 24321
rect 419 24269 421 24321
rect 365 24267 421 24269
rect -1205 23977 -1149 24033
rect -425 24051 -369 24053
rect -425 23999 -423 24051
rect -423 23999 -371 24051
rect -371 23999 -369 24051
rect -425 23997 -369 23999
rect -115 24051 -59 24053
rect -115 23999 -113 24051
rect -113 23999 -61 24051
rect -61 23999 -59 24051
rect -115 23997 -59 23999
rect 205 24051 261 24053
rect 205 23999 207 24051
rect 207 23999 259 24051
rect 259 23999 261 24051
rect 205 23997 261 23999
rect 525 24051 581 24053
rect 525 23999 527 24051
rect 527 23999 579 24051
rect 579 23999 581 24051
rect 525 23997 581 23999
rect 1635 26851 1691 26853
rect 1635 26799 1637 26851
rect 1637 26799 1689 26851
rect 1689 26799 1691 26851
rect 1635 26797 1691 26799
rect 2000 26042 2056 26098
rect 2000 25822 2056 25878
rect 2985 29637 3041 29693
rect -1205 23727 -1149 23783
rect 1315 23977 1371 24033
rect -425 23761 -369 23763
rect -425 23709 -423 23761
rect -423 23709 -371 23761
rect -371 23709 -369 23761
rect -425 23707 -369 23709
rect -115 23761 -59 23763
rect -115 23709 -113 23761
rect -113 23709 -61 23761
rect -61 23709 -59 23761
rect -115 23707 -59 23709
rect 205 23761 261 23763
rect 205 23709 207 23761
rect 207 23709 259 23761
rect 259 23709 261 23761
rect 205 23707 261 23709
rect 525 23761 581 23763
rect 525 23709 527 23761
rect 527 23709 579 23761
rect 579 23709 581 23761
rect 525 23707 581 23709
rect 1315 23727 1371 23783
rect 1760 25482 1816 25538
rect 1760 25262 1816 25318
rect 1760 24522 1816 24578
rect 1760 24302 1816 24358
rect -110 23292 106 23508
rect -1575 23091 -1519 23093
rect -1575 23039 -1573 23091
rect -1573 23039 -1521 23091
rect -1521 23039 -1519 23091
rect -1575 23037 -1519 23039
rect -1055 23091 -999 23093
rect -1055 23039 -1053 23091
rect -1053 23039 -1001 23091
rect -1001 23039 -999 23091
rect -1055 23037 -999 23039
rect -545 23091 -489 23093
rect -545 23039 -543 23091
rect -543 23039 -491 23091
rect -491 23039 -489 23091
rect -545 23037 -489 23039
rect -25 23091 31 23093
rect -25 23039 -23 23091
rect -23 23039 29 23091
rect 29 23039 31 23091
rect -25 23037 31 23039
rect 485 23091 541 23093
rect 485 23039 487 23091
rect 487 23039 539 23091
rect 539 23039 541 23091
rect 485 23037 541 23039
rect 1005 23091 1061 23093
rect 1005 23039 1007 23091
rect 1007 23039 1059 23091
rect 1059 23039 1061 23091
rect 1005 23037 1061 23039
rect 1525 23091 1581 23093
rect 1525 23039 1527 23091
rect 1527 23039 1579 23091
rect 1579 23039 1581 23091
rect 1525 23037 1581 23039
rect -1575 22911 -1519 22913
rect -1575 22859 -1573 22911
rect -1573 22859 -1521 22911
rect -1521 22859 -1519 22911
rect -1575 22857 -1519 22859
rect -1055 22911 -999 22913
rect -1055 22859 -1053 22911
rect -1053 22859 -1001 22911
rect -1001 22859 -999 22911
rect -1055 22857 -999 22859
rect -545 22911 -489 22913
rect -545 22859 -543 22911
rect -543 22859 -491 22911
rect -491 22859 -489 22911
rect -545 22857 -489 22859
rect -25 22911 31 22913
rect -25 22859 -23 22911
rect -23 22859 29 22911
rect 29 22859 31 22911
rect -25 22857 31 22859
rect 485 22911 541 22913
rect 485 22859 487 22911
rect 487 22859 539 22911
rect 539 22859 541 22911
rect 485 22857 541 22859
rect 1005 22911 1061 22913
rect 1005 22859 1007 22911
rect 1007 22859 1059 22911
rect 1059 22859 1061 22911
rect 1005 22857 1061 22859
rect 1525 22911 1581 22913
rect 1525 22859 1527 22911
rect 1527 22859 1579 22911
rect 1579 22859 1581 22911
rect 1525 22857 1581 22859
rect -1315 22421 -1259 22423
rect -1315 22369 -1313 22421
rect -1313 22369 -1261 22421
rect -1261 22369 -1259 22421
rect -1315 22367 -1259 22369
rect -805 22421 -749 22423
rect -805 22369 -803 22421
rect -803 22369 -751 22421
rect -751 22369 -749 22421
rect -805 22367 -749 22369
rect -285 22421 -229 22423
rect -285 22369 -283 22421
rect -283 22369 -231 22421
rect -231 22369 -229 22421
rect -285 22367 -229 22369
rect 235 22421 291 22423
rect 235 22369 237 22421
rect 237 22369 289 22421
rect 289 22369 291 22421
rect 235 22367 291 22369
rect 745 22421 801 22423
rect 745 22369 747 22421
rect 747 22369 799 22421
rect 799 22369 801 22421
rect 745 22367 801 22369
rect 1265 22421 1321 22423
rect 1265 22369 1267 22421
rect 1267 22369 1319 22421
rect 1319 22369 1321 22421
rect 1265 22367 1321 22369
rect -1315 22241 -1259 22243
rect -1315 22189 -1313 22241
rect -1313 22189 -1261 22241
rect -1261 22189 -1259 22241
rect -1315 22187 -1259 22189
rect -805 22241 -749 22243
rect -805 22189 -803 22241
rect -803 22189 -751 22241
rect -751 22189 -749 22241
rect -805 22187 -749 22189
rect -285 22241 -229 22243
rect -285 22189 -283 22241
rect -283 22189 -231 22241
rect -231 22189 -229 22241
rect -285 22187 -229 22189
rect 235 22241 291 22243
rect 235 22189 237 22241
rect 237 22189 289 22241
rect 289 22189 291 22241
rect 235 22187 291 22189
rect 745 22241 801 22243
rect 745 22189 747 22241
rect 747 22189 799 22241
rect 799 22189 801 22241
rect 745 22187 801 22189
rect 1265 22241 1321 22243
rect 1265 22189 1267 22241
rect 1267 22189 1319 22241
rect 1319 22189 1321 22241
rect 1265 22187 1321 22189
rect -105 21777 111 21993
rect -1835 21571 -1779 21573
rect -1835 21519 -1833 21571
rect -1833 21519 -1781 21571
rect -1781 21519 -1779 21571
rect -1835 21517 -1779 21519
rect -1315 21571 -1259 21573
rect -1315 21519 -1313 21571
rect -1313 21519 -1261 21571
rect -1261 21519 -1259 21571
rect -1315 21517 -1259 21519
rect -805 21571 -749 21573
rect -805 21519 -803 21571
rect -803 21519 -751 21571
rect -751 21519 -749 21571
rect -805 21517 -749 21519
rect -285 21571 -229 21573
rect -285 21519 -283 21571
rect -283 21519 -231 21571
rect -231 21519 -229 21571
rect -285 21517 -229 21519
rect 225 21571 281 21573
rect 225 21519 227 21571
rect 227 21519 279 21571
rect 279 21519 281 21571
rect 225 21517 281 21519
rect 745 21571 801 21573
rect 745 21519 747 21571
rect 747 21519 799 21571
rect 799 21519 801 21571
rect 745 21517 801 21519
rect 1265 21571 1321 21573
rect 1265 21519 1267 21571
rect 1267 21519 1319 21571
rect 1319 21519 1321 21571
rect 1265 21517 1321 21519
rect 1775 21571 1831 21573
rect 1775 21519 1777 21571
rect 1777 21519 1829 21571
rect 1829 21519 1831 21571
rect 1775 21517 1831 21519
rect -1835 21391 -1779 21393
rect -1835 21339 -1833 21391
rect -1833 21339 -1781 21391
rect -1781 21339 -1779 21391
rect -1835 21337 -1779 21339
rect -1315 21391 -1259 21393
rect -1315 21339 -1313 21391
rect -1313 21339 -1261 21391
rect -1261 21339 -1259 21391
rect -1315 21337 -1259 21339
rect -805 21391 -749 21393
rect -805 21339 -803 21391
rect -803 21339 -751 21391
rect -751 21339 -749 21391
rect -805 21337 -749 21339
rect -285 21391 -229 21393
rect -285 21339 -283 21391
rect -283 21339 -231 21391
rect -231 21339 -229 21391
rect -285 21337 -229 21339
rect 225 21391 281 21393
rect 225 21339 227 21391
rect 227 21339 279 21391
rect 279 21339 281 21391
rect 225 21337 281 21339
rect 745 21391 801 21393
rect 745 21339 747 21391
rect 747 21339 799 21391
rect 799 21339 801 21391
rect 745 21337 801 21339
rect 1265 21391 1321 21393
rect 1265 21339 1267 21391
rect 1267 21339 1319 21391
rect 1319 21339 1321 21391
rect 1265 21337 1321 21339
rect 1775 21391 1831 21393
rect 1775 21339 1777 21391
rect 1777 21339 1829 21391
rect 1829 21339 1831 21391
rect 1775 21337 1831 21339
rect 2985 23027 3041 23083
rect 2985 22867 3041 22923
rect -1575 20901 -1519 20903
rect -1575 20849 -1573 20901
rect -1573 20849 -1521 20901
rect -1521 20849 -1519 20901
rect -1575 20847 -1519 20849
rect -1065 20901 -1009 20903
rect -1065 20849 -1063 20901
rect -1063 20849 -1011 20901
rect -1011 20849 -1009 20901
rect -1065 20847 -1009 20849
rect -545 20901 -489 20903
rect -545 20849 -543 20901
rect -543 20849 -491 20901
rect -491 20849 -489 20901
rect -545 20847 -489 20849
rect -25 20901 31 20903
rect -25 20849 -23 20901
rect -23 20849 29 20901
rect 29 20849 31 20901
rect -25 20847 31 20849
rect 485 20901 541 20903
rect 485 20849 487 20901
rect 487 20849 539 20901
rect 539 20849 541 20901
rect 485 20847 541 20849
rect 1005 20901 1061 20903
rect 1005 20849 1007 20901
rect 1007 20849 1059 20901
rect 1059 20849 1061 20901
rect 1005 20847 1061 20849
rect 1515 20901 1571 20903
rect 1515 20849 1517 20901
rect 1517 20849 1569 20901
rect 1569 20849 1571 20901
rect 1515 20847 1571 20849
rect -1575 20721 -1519 20723
rect -1575 20669 -1573 20721
rect -1573 20669 -1521 20721
rect -1521 20669 -1519 20721
rect -1575 20667 -1519 20669
rect -1065 20721 -1009 20723
rect -1065 20669 -1063 20721
rect -1063 20669 -1011 20721
rect -1011 20669 -1009 20721
rect -1065 20667 -1009 20669
rect -545 20721 -489 20723
rect -545 20669 -543 20721
rect -543 20669 -491 20721
rect -491 20669 -489 20721
rect -545 20667 -489 20669
rect -25 20721 31 20723
rect -25 20669 -23 20721
rect -23 20669 29 20721
rect 29 20669 31 20721
rect -25 20667 31 20669
rect 485 20721 541 20723
rect 485 20669 487 20721
rect 487 20669 539 20721
rect 539 20669 541 20721
rect 485 20667 541 20669
rect 1005 20721 1061 20723
rect 1005 20669 1007 20721
rect 1007 20669 1059 20721
rect 1059 20669 1061 20721
rect 1005 20667 1061 20669
rect 1515 20721 1571 20723
rect 1515 20669 1517 20721
rect 1517 20669 1569 20721
rect 1569 20669 1571 20721
rect 1515 20667 1571 20669
rect 2638 21440 2878 21680
rect 2968 21440 3208 21680
rect -105 20247 111 20463
rect -3220 19480 -3060 19640
rect -2160 19480 -2000 19640
rect -700 19480 -540 19640
rect -3220 18900 -3060 19060
rect -2160 18900 -2000 19060
rect -700 18900 -540 19060
rect 520 19480 680 19640
rect 2000 19480 2160 19640
rect 3000 19480 3160 19640
rect 520 18900 680 19060
rect -840 17530 -620 17680
rect -3200 16990 -3020 17120
rect -2060 16990 -1880 17120
rect -320 17530 -100 17680
rect 100 17530 320 17680
rect -1080 17000 -900 17130
rect 2000 18900 2160 19060
rect 3000 18900 3160 19060
rect 650 17530 870 17680
rect -310 17000 -130 17130
rect 130 17000 310 17130
rect 850 16990 1030 17120
rect 1920 17000 2100 17130
rect 2920 17000 3100 17130
rect -3240 15100 -3120 15220
rect 3130 15100 3250 15220
rect -3240 12100 -3120 12220
rect 3130 12100 3250 12220
rect -3240 9100 -3120 9220
rect 3130 9100 3250 9220
rect -3240 6100 -3120 6220
rect 3130 6100 3250 6220
rect -3240 3100 -3120 3220
rect 3130 3100 3250 3220
rect -2860 1480 -1690 1890
rect -1350 1480 -180 1890
rect 170 1480 1340 1890
rect 1690 1490 2860 1900
<< metal3 >>
rect -7922 37000 -7712 37020
rect -7922 36930 -7902 37000
rect -7832 36930 -7802 37000
rect -7732 36930 -7712 37000
rect -7922 36870 -7712 36930
rect 7978 37000 8188 37020
rect 7978 36930 7998 37000
rect 8068 36930 8098 37000
rect 8168 36930 8188 37000
rect -7922 36800 -7902 36870
rect -7832 36800 -7802 36870
rect -7732 36800 -7712 36870
rect -7922 30620 -7712 36800
rect -7402 36869 -4002 36889
rect -7402 36805 -7374 36869
rect -7310 36805 -7294 36869
rect -7230 36805 -7214 36869
rect -7150 36805 -7134 36869
rect -7070 36805 -7054 36869
rect -6990 36805 -6974 36869
rect -6910 36805 -6894 36869
rect -6830 36805 -6814 36869
rect -6750 36805 -6734 36869
rect -6670 36805 -6654 36869
rect -6590 36805 -6574 36869
rect -6510 36805 -6494 36869
rect -6430 36805 -6414 36869
rect -6350 36805 -6334 36869
rect -6270 36805 -6254 36869
rect -6190 36805 -6174 36869
rect -6110 36805 -6094 36869
rect -6030 36805 -6014 36869
rect -5950 36805 -5934 36869
rect -5870 36805 -5854 36869
rect -5790 36805 -5774 36869
rect -5710 36805 -5694 36869
rect -5630 36805 -5614 36869
rect -5550 36805 -5534 36869
rect -5470 36805 -5454 36869
rect -5390 36805 -5374 36869
rect -5310 36805 -5294 36869
rect -5230 36805 -5214 36869
rect -5150 36805 -5134 36869
rect -5070 36805 -5054 36869
rect -4990 36805 -4974 36869
rect -4910 36805 -4894 36869
rect -4830 36805 -4814 36869
rect -4750 36805 -4734 36869
rect -4670 36805 -4654 36869
rect -4590 36805 -4574 36869
rect -4510 36805 -4494 36869
rect -4430 36805 -4414 36869
rect -4350 36805 -4334 36869
rect -4270 36805 -4254 36869
rect -4190 36805 -4174 36869
rect -4110 36805 -4094 36869
rect -4030 36805 -4002 36869
rect -7402 33390 -4002 36805
rect -3602 36869 -202 36889
rect -3602 36805 -3574 36869
rect -3510 36805 -3494 36869
rect -3430 36805 -3414 36869
rect -3350 36805 -3334 36869
rect -3270 36805 -3254 36869
rect -3190 36805 -3174 36869
rect -3110 36805 -3094 36869
rect -3030 36805 -3014 36869
rect -2950 36805 -2934 36869
rect -2870 36805 -2854 36869
rect -2790 36805 -2774 36869
rect -2710 36805 -2694 36869
rect -2630 36805 -2614 36869
rect -2550 36805 -2534 36869
rect -2470 36805 -2454 36869
rect -2390 36805 -2374 36869
rect -2310 36805 -2294 36869
rect -2230 36805 -2214 36869
rect -2150 36805 -2134 36869
rect -2070 36805 -2054 36869
rect -1990 36805 -1974 36869
rect -1910 36805 -1894 36869
rect -1830 36805 -1814 36869
rect -1750 36805 -1734 36869
rect -1670 36805 -1654 36869
rect -1590 36805 -1574 36869
rect -1510 36805 -1494 36869
rect -1430 36805 -1414 36869
rect -1350 36805 -1334 36869
rect -1270 36805 -1254 36869
rect -1190 36805 -1174 36869
rect -1110 36805 -1094 36869
rect -1030 36805 -1014 36869
rect -950 36805 -934 36869
rect -870 36805 -854 36869
rect -790 36805 -774 36869
rect -710 36805 -694 36869
rect -630 36805 -614 36869
rect -550 36805 -534 36869
rect -470 36805 -454 36869
rect -390 36805 -374 36869
rect -310 36805 -294 36869
rect -230 36805 -202 36869
rect -3602 33390 -202 36805
rect 198 36869 3598 36889
rect 198 36805 226 36869
rect 290 36805 306 36869
rect 370 36805 386 36869
rect 450 36805 466 36869
rect 530 36805 546 36869
rect 610 36805 626 36869
rect 690 36805 706 36869
rect 770 36805 786 36869
rect 850 36805 866 36869
rect 930 36805 946 36869
rect 1010 36805 1026 36869
rect 1090 36805 1106 36869
rect 1170 36805 1186 36869
rect 1250 36805 1266 36869
rect 1330 36805 1346 36869
rect 1410 36805 1426 36869
rect 1490 36805 1506 36869
rect 1570 36805 1586 36869
rect 1650 36805 1666 36869
rect 1730 36805 1746 36869
rect 1810 36805 1826 36869
rect 1890 36805 1906 36869
rect 1970 36805 1986 36869
rect 2050 36805 2066 36869
rect 2130 36805 2146 36869
rect 2210 36805 2226 36869
rect 2290 36805 2306 36869
rect 2370 36805 2386 36869
rect 2450 36805 2466 36869
rect 2530 36805 2546 36869
rect 2610 36805 2626 36869
rect 2690 36805 2706 36869
rect 2770 36805 2786 36869
rect 2850 36805 2866 36869
rect 2930 36805 2946 36869
rect 3010 36805 3026 36869
rect 3090 36805 3106 36869
rect 3170 36805 3186 36869
rect 3250 36805 3266 36869
rect 3330 36805 3346 36869
rect 3410 36805 3426 36869
rect 3490 36805 3506 36869
rect 3570 36805 3598 36869
rect 198 33390 3598 36805
rect 3998 36869 7398 36889
rect 3998 36805 4026 36869
rect 4090 36805 4106 36869
rect 4170 36805 4186 36869
rect 4250 36805 4266 36869
rect 4330 36805 4346 36869
rect 4410 36805 4426 36869
rect 4490 36805 4506 36869
rect 4570 36805 4586 36869
rect 4650 36805 4666 36869
rect 4730 36805 4746 36869
rect 4810 36805 4826 36869
rect 4890 36805 4906 36869
rect 4970 36805 4986 36869
rect 5050 36805 5066 36869
rect 5130 36805 5146 36869
rect 5210 36805 5226 36869
rect 5290 36805 5306 36869
rect 5370 36805 5386 36869
rect 5450 36805 5466 36869
rect 5530 36805 5546 36869
rect 5610 36805 5626 36869
rect 5690 36805 5706 36869
rect 5770 36805 5786 36869
rect 5850 36805 5866 36869
rect 5930 36805 5946 36869
rect 6010 36805 6026 36869
rect 6090 36805 6106 36869
rect 6170 36805 6186 36869
rect 6250 36805 6266 36869
rect 6330 36805 6346 36869
rect 6410 36805 6426 36869
rect 6490 36805 6506 36869
rect 6570 36805 6586 36869
rect 6650 36805 6666 36869
rect 6730 36805 6746 36869
rect 6810 36805 6826 36869
rect 6890 36805 6906 36869
rect 6970 36805 6986 36869
rect 7050 36805 7066 36869
rect 7130 36805 7146 36869
rect 7210 36805 7226 36869
rect 7290 36805 7306 36869
rect 7370 36805 7398 36869
rect 3998 33390 7398 36805
rect 7978 36870 8188 36930
rect 7978 36800 7998 36870
rect 8068 36800 8098 36870
rect 8168 36800 8188 36870
rect -652 31377 -362 31405
rect -652 31153 -619 31377
rect -395 31153 -362 31377
rect -652 31125 -362 31153
rect 398 31377 688 31405
rect 398 31153 431 31377
rect 655 31153 688 31377
rect 398 31125 688 31153
rect -3192 30925 3198 30930
rect -3202 30913 3208 30925
rect -3202 30857 -3185 30913
rect -3129 30857 -2865 30913
rect -2809 30887 -2555 30913
rect -2809 30857 -2799 30887
rect -3202 30845 -2799 30857
rect -3192 30685 -2799 30845
rect -7922 30560 -7912 30620
rect -7852 30560 -7792 30620
rect -7732 30560 -7712 30620
rect -3202 30673 -2799 30685
rect -3202 30617 -3185 30673
rect -3129 30617 -2865 30673
rect -2809 30663 -2799 30673
rect -2575 30857 -2555 30887
rect -2499 30857 -2235 30913
rect -2179 30857 -1925 30913
rect -1869 30857 -1605 30913
rect -1549 30857 -1285 30913
rect -1229 30857 -975 30913
rect -919 30877 -655 30913
rect -919 30857 -899 30877
rect -2575 30673 -899 30857
rect -2575 30663 -2555 30673
rect -2809 30617 -2555 30663
rect -2499 30617 -2235 30673
rect -2179 30617 -1925 30673
rect -1869 30617 -1605 30673
rect -1549 30617 -1285 30673
rect -1229 30617 -975 30673
rect -919 30653 -899 30673
rect -675 30857 -655 30877
rect -599 30857 -335 30913
rect -279 30857 -25 30913
rect 31 30857 295 30913
rect 351 30857 605 30913
rect 661 30877 925 30913
rect 661 30857 681 30877
rect -675 30673 681 30857
rect -675 30653 -655 30673
rect -919 30617 -655 30653
rect -599 30617 -335 30673
rect -279 30617 -25 30673
rect 31 30617 295 30673
rect 351 30617 605 30673
rect 661 30653 681 30673
rect 905 30857 925 30877
rect 981 30857 1245 30913
rect 1301 30857 1555 30913
rect 1611 30857 1875 30913
rect 1931 30857 2185 30913
rect 2241 30857 2505 30913
rect 2561 30877 2825 30913
rect 2561 30857 2581 30877
rect 905 30673 2581 30857
rect 905 30653 925 30673
rect 661 30617 925 30653
rect 981 30617 1245 30673
rect 1301 30617 1555 30673
rect 1611 30617 1875 30673
rect 1931 30617 2185 30673
rect 2241 30617 2505 30673
rect 2561 30653 2581 30673
rect 2805 30857 2825 30877
rect 2881 30857 3135 30913
rect 3191 30857 3208 30913
rect 2805 30845 3208 30857
rect 2805 30685 3198 30845
rect 2805 30673 3208 30685
rect 2805 30653 2825 30673
rect 2561 30617 2825 30653
rect 2881 30617 3135 30673
rect 3191 30617 3208 30673
rect -3202 30605 3208 30617
rect 7978 30618 8188 36800
rect -3192 30600 3198 30605
rect -7922 30520 -7712 30560
rect 7978 30562 8000 30618
rect 8056 30562 8110 30618
rect 8166 30562 8188 30618
rect 7978 30530 8188 30562
rect -3192 30303 3198 30320
rect -3192 30247 -3025 30303
rect -2969 30247 -2715 30303
rect -2659 30247 -2395 30303
rect -2339 30247 -2075 30303
rect -2019 30247 -1765 30303
rect -1709 30247 -1445 30303
rect -1389 30247 -1135 30303
rect -1079 30247 -815 30303
rect -759 30247 -495 30303
rect -439 30247 -185 30303
rect -129 30247 135 30303
rect 191 30247 455 30303
rect 511 30247 765 30303
rect 821 30247 1085 30303
rect 1141 30247 1395 30303
rect 1451 30247 1715 30303
rect 1771 30247 2035 30303
rect 2091 30247 2345 30303
rect 2401 30247 2665 30303
rect 2721 30247 2985 30303
rect 3041 30247 3198 30303
rect -3192 30063 3198 30247
rect -3192 30007 -3025 30063
rect -2969 30007 -2715 30063
rect -2659 30007 -2395 30063
rect -2339 30007 -2075 30063
rect -2019 30007 -1765 30063
rect -1709 30007 -1445 30063
rect -1389 30007 -1135 30063
rect -1079 30007 -815 30063
rect -759 30007 -495 30063
rect -439 30007 -185 30063
rect -129 30007 135 30063
rect 191 30007 455 30063
rect 511 30007 765 30063
rect 821 30007 1085 30063
rect 1141 30007 1395 30063
rect 1451 30007 1715 30063
rect 1771 30007 2035 30063
rect 2091 30007 2345 30063
rect 2401 30007 2665 30063
rect 2721 30007 2985 30063
rect 3041 30007 3198 30063
rect -3192 29990 3198 30007
rect -652 29737 -362 29765
rect -3702 29697 -2932 29730
rect -3702 29633 -3669 29697
rect -3605 29693 -2932 29697
rect -3605 29637 -3025 29693
rect -2969 29637 -2932 29693
rect -3605 29633 -2932 29637
rect -3702 29600 -2932 29633
rect -652 29513 -619 29737
rect -395 29513 -362 29737
rect -652 29485 -362 29513
rect 398 29737 688 29765
rect 398 29513 431 29737
rect 655 29513 688 29737
rect 2948 29697 3478 29730
rect 2948 29693 3381 29697
rect 2948 29637 2985 29693
rect 3041 29637 3381 29693
rect 2948 29633 3381 29637
rect 3445 29633 3478 29697
rect 2948 29600 3478 29633
rect 398 29485 688 29513
rect -1692 29255 1698 29260
rect -1702 29243 1698 29255
rect -1702 29187 -1685 29243
rect -1629 29187 -1365 29243
rect -1309 29222 -1055 29243
rect -1309 29187 -1294 29222
rect -1702 29175 -1294 29187
rect -1692 29045 -1294 29175
rect -1702 29033 -1294 29045
rect -1702 28977 -1685 29033
rect -1629 28977 -1365 29033
rect -1309 28998 -1294 29033
rect -1070 29187 -1055 29222
rect -999 29187 -735 29243
rect -679 29187 -415 29243
rect -359 29187 -105 29243
rect -49 29222 215 29243
rect -49 29187 -24 29222
rect -1070 29033 -24 29187
rect -1070 28998 -1055 29033
rect -1309 28977 -1055 28998
rect -999 28977 -735 29033
rect -679 28977 -415 29033
rect -359 28977 -105 29033
rect -49 28998 -24 29033
rect 200 29187 215 29222
rect 271 29187 535 29243
rect 591 29187 845 29243
rect 901 29187 1165 29243
rect 1221 29222 1475 29243
rect 1221 29187 1236 29222
rect 200 29033 1236 29187
rect 200 28998 215 29033
rect -49 28977 215 28998
rect 271 28977 535 29033
rect 591 28977 845 29033
rect 901 28977 1165 29033
rect 1221 28998 1236 29033
rect 1460 29187 1475 29222
rect 1531 29187 1698 29243
rect 1460 29033 1698 29187
rect 1460 28998 1475 29033
rect 1221 28977 1475 28998
rect 1531 28977 1698 29033
rect -1702 28965 1698 28977
rect -1692 28960 1698 28965
rect -2112 28603 2108 28620
rect -2112 28588 -1525 28603
rect -2112 28532 -2060 28588
rect -2004 28547 -1525 28588
rect -1469 28547 -1205 28603
rect -1149 28547 -895 28603
rect -839 28547 -575 28603
rect -519 28547 -255 28603
rect -199 28547 55 28603
rect 111 28547 375 28603
rect 431 28547 685 28603
rect 741 28547 1005 28603
rect 1061 28547 1325 28603
rect 1381 28547 1635 28603
rect 1691 28588 2108 28603
rect 1691 28547 2000 28588
rect -2004 28532 2000 28547
rect 2056 28532 2108 28588
rect -2112 28408 2108 28532
rect -2112 28352 -2060 28408
rect -2004 28393 2000 28408
rect -2004 28352 -1525 28393
rect -2112 28337 -1525 28352
rect -1469 28337 -1205 28393
rect -1149 28337 -895 28393
rect -839 28337 -575 28393
rect -519 28337 -255 28393
rect -199 28337 55 28393
rect 111 28337 375 28393
rect 431 28337 685 28393
rect 741 28337 1005 28393
rect 1061 28337 1325 28393
rect 1381 28337 1635 28393
rect 1691 28352 2000 28393
rect 2056 28352 2108 28408
rect 1691 28337 2108 28352
rect -2112 28320 2108 28337
rect -882 28132 -602 28155
rect -882 27908 -854 28132
rect -630 27908 -602 28132
rect -882 27885 -602 27908
rect 618 28132 898 28155
rect 618 27908 646 28132
rect 870 27908 898 28132
rect 618 27885 898 27908
rect -1692 27705 1698 27710
rect -1702 27693 1698 27705
rect -1702 27637 -1685 27693
rect -1629 27637 -1365 27693
rect -1309 27672 -1055 27693
rect -1309 27637 -1294 27672
rect -1702 27625 -1294 27637
rect -1692 27495 -1294 27625
rect -1702 27483 -1294 27495
rect -1702 27427 -1685 27483
rect -1629 27427 -1365 27483
rect -1309 27448 -1294 27483
rect -1070 27637 -1055 27672
rect -999 27637 -735 27693
rect -679 27637 -415 27693
rect -359 27637 -105 27693
rect -49 27672 215 27693
rect -49 27637 -24 27672
rect -1070 27483 -24 27637
rect -1070 27448 -1055 27483
rect -1309 27427 -1055 27448
rect -999 27427 -735 27483
rect -679 27427 -415 27483
rect -359 27427 -105 27483
rect -49 27448 -24 27483
rect 200 27637 215 27672
rect 271 27637 525 27693
rect 581 27637 845 27693
rect 901 27637 1165 27693
rect 1221 27672 1475 27693
rect 1221 27637 1236 27672
rect 200 27483 1236 27637
rect 200 27448 215 27483
rect -49 27427 215 27448
rect 271 27427 525 27483
rect 581 27427 845 27483
rect 901 27427 1165 27483
rect 1221 27448 1236 27483
rect 1460 27637 1475 27672
rect 1531 27637 1698 27693
rect 1460 27483 1698 27637
rect 1460 27448 1475 27483
rect 1221 27427 1475 27448
rect 1531 27427 1698 27483
rect -1702 27415 1698 27427
rect -1692 27410 1698 27415
rect -1692 27075 1698 27080
rect -1692 27063 1708 27075
rect -1692 27007 -1525 27063
rect -1469 27007 -1205 27063
rect -1149 27007 -895 27063
rect -839 27007 -575 27063
rect -519 27007 -265 27063
rect -209 27007 55 27063
rect 111 27007 375 27063
rect 431 27007 685 27063
rect 741 27007 1005 27063
rect 1061 27007 1315 27063
rect 1371 27007 1635 27063
rect 1691 27007 1708 27063
rect -1692 26995 1708 27007
rect -1692 26865 1698 26995
rect -1692 26853 1708 26865
rect -1692 26797 -1525 26853
rect -1469 26797 -1205 26853
rect -1149 26797 -895 26853
rect -839 26797 -575 26853
rect -519 26797 -265 26853
rect -209 26797 55 26853
rect 111 26797 375 26853
rect 431 26797 685 26853
rect 741 26797 1005 26853
rect 1061 26797 1315 26853
rect 1371 26797 1635 26853
rect 1691 26797 1708 26853
rect -1692 26785 1708 26797
rect -1692 26780 1698 26785
rect -2112 26133 2108 26150
rect -2112 26098 -585 26133
rect -2112 26042 -2060 26098
rect -2004 26077 -585 26098
rect -529 26077 -265 26133
rect -209 26077 45 26133
rect 101 26077 365 26133
rect 421 26098 2108 26133
rect 421 26077 2000 26098
rect -2004 26042 2000 26077
rect 2056 26042 2108 26098
rect -2112 25878 2108 26042
rect -2112 25822 -2060 25878
rect -2004 25843 2000 25878
rect -2004 25822 -585 25843
rect -2112 25787 -585 25822
rect -529 25787 -265 25843
rect -209 25787 45 25843
rect 101 25787 365 25843
rect 421 25822 2000 25843
rect 2056 25822 2108 25878
rect 421 25787 2108 25822
rect -2112 25770 2108 25787
rect -1872 25573 1868 25590
rect -1872 25538 -425 25573
rect -1872 25482 -1820 25538
rect -1764 25517 -425 25538
rect -369 25517 -115 25573
rect -59 25517 205 25573
rect 261 25517 525 25573
rect 581 25538 1868 25573
rect 581 25517 1760 25538
rect -1764 25482 1760 25517
rect 1816 25482 1868 25538
rect -1872 25318 1868 25482
rect -1872 25262 -1820 25318
rect -1764 25283 1760 25318
rect -1764 25262 -425 25283
rect -1872 25227 -425 25262
rect -369 25227 -115 25283
rect -59 25227 205 25283
rect 261 25227 525 25283
rect 581 25262 1760 25283
rect 1816 25262 1868 25318
rect 581 25227 1868 25262
rect -1872 25210 1868 25227
rect -142 25032 138 25055
rect -142 24808 -114 25032
rect 110 24808 138 25032
rect -142 24785 138 24808
rect -1872 24613 1868 24630
rect -1872 24578 -585 24613
rect -1872 24522 -1820 24578
rect -1764 24557 -585 24578
rect -529 24557 -265 24613
rect -209 24557 45 24613
rect 101 24557 365 24613
rect 421 24578 1868 24613
rect 421 24557 1760 24578
rect -1764 24522 1760 24557
rect 1816 24522 1868 24578
rect -1872 24358 1868 24522
rect -1872 24302 -1820 24358
rect -1764 24323 1760 24358
rect -1764 24302 -585 24323
rect -1872 24267 -585 24302
rect -529 24267 -265 24323
rect -209 24267 45 24323
rect 101 24267 365 24323
rect 421 24302 1760 24323
rect 1816 24302 1868 24358
rect 421 24267 1868 24302
rect -1872 24250 1868 24267
rect -1242 24053 1408 24070
rect -1242 24033 -425 24053
rect -1242 23977 -1205 24033
rect -1149 23997 -425 24033
rect -369 23997 -115 24053
rect -59 23997 205 24053
rect 261 23997 525 24053
rect 581 24033 1408 24053
rect 581 23997 1315 24033
rect -1149 23977 1315 23997
rect 1371 23977 1408 24033
rect -1242 23783 1408 23977
rect -1242 23727 -1205 23783
rect -1149 23763 1315 23783
rect -1149 23727 -425 23763
rect -1242 23707 -425 23727
rect -369 23707 -115 23763
rect -59 23707 205 23763
rect 261 23707 525 23763
rect 581 23727 1315 23763
rect 1371 23727 1408 23783
rect 581 23707 1408 23727
rect -1242 23690 1408 23707
rect -142 23512 138 23535
rect -142 23288 -114 23512
rect 110 23288 138 23512
rect -142 23265 138 23288
rect -3062 23093 3078 23110
rect -3062 23083 -1575 23093
rect -3062 23027 -3025 23083
rect -2969 23037 -1575 23083
rect -1519 23037 -1055 23093
rect -999 23037 -545 23093
rect -489 23037 -25 23093
rect 31 23037 485 23093
rect 541 23037 1005 23093
rect 1061 23037 1525 23093
rect 1581 23083 3078 23093
rect 1581 23037 2985 23083
rect -2969 23027 2985 23037
rect 3041 23027 3078 23083
rect -3062 22923 3078 23027
rect -3062 22867 -3025 22923
rect -2969 22913 2985 22923
rect -2969 22867 -1575 22913
rect -3062 22857 -1575 22867
rect -1519 22857 -1055 22913
rect -999 22857 -545 22913
rect -489 22857 -25 22913
rect 31 22857 485 22913
rect 541 22857 1005 22913
rect 1061 22857 1525 22913
rect 1581 22867 2985 22913
rect 3041 22867 3078 22923
rect 1581 22857 3078 22867
rect -3062 22840 3078 22857
rect -1582 22423 1588 22440
rect -1582 22367 -1315 22423
rect -1259 22417 -805 22423
rect -1259 22367 -1139 22417
rect -1582 22243 -1139 22367
rect -1582 22187 -1315 22243
rect -1259 22193 -1139 22243
rect -915 22367 -805 22417
rect -749 22367 -285 22423
rect -229 22367 235 22423
rect 291 22367 745 22423
rect 801 22417 1265 22423
rect 801 22367 921 22417
rect -915 22243 921 22367
rect -915 22193 -805 22243
rect -1259 22187 -805 22193
rect -749 22187 -285 22243
rect -229 22187 235 22243
rect 291 22187 745 22243
rect 801 22193 921 22243
rect 1145 22367 1265 22417
rect 1321 22367 1588 22423
rect 1145 22243 1588 22367
rect 1145 22193 1265 22243
rect 801 22187 1265 22193
rect 1321 22187 1588 22243
rect -1582 22170 1588 22187
rect -132 21997 138 22015
rect -132 21773 -109 21997
rect 115 21773 138 21997
rect -132 21755 138 21773
rect -3272 21722 -2662 21745
rect -3272 21338 -3239 21722
rect -2695 21338 -2662 21722
rect 2628 21680 2888 21685
rect -1842 21585 1838 21590
rect -1852 21573 1848 21585
rect -1852 21517 -1835 21573
rect -1779 21517 -1315 21573
rect -1259 21517 -805 21573
rect -749 21517 -285 21573
rect -229 21517 225 21573
rect 281 21517 745 21573
rect 801 21517 1265 21573
rect 1321 21517 1775 21573
rect 1831 21517 1848 21573
rect -1852 21505 1848 21517
rect -1842 21405 1838 21505
rect 2628 21440 2638 21680
rect 2878 21440 2888 21680
rect 2628 21435 2888 21440
rect 2958 21680 3218 21685
rect 2958 21440 2968 21680
rect 3208 21440 3218 21680
rect 2958 21435 3218 21440
rect -3272 21315 -2662 21338
rect -1852 21393 1848 21405
rect -1852 21337 -1835 21393
rect -1779 21337 -1315 21393
rect -1259 21337 -805 21393
rect -749 21337 -285 21393
rect -229 21337 225 21393
rect 281 21337 745 21393
rect 801 21337 1265 21393
rect 1321 21337 1775 21393
rect 1831 21337 1848 21393
rect -1852 21325 1848 21337
rect -1842 21320 1838 21325
rect -1842 20903 1838 20920
rect -1842 20847 -1575 20903
rect -1519 20897 -1065 20903
rect -1519 20847 -1399 20897
rect -1842 20723 -1399 20847
rect -1842 20667 -1575 20723
rect -1519 20673 -1399 20723
rect -1175 20847 -1065 20897
rect -1009 20847 -545 20903
rect -489 20847 -25 20903
rect 31 20847 485 20903
rect 541 20847 1005 20903
rect 1061 20897 1515 20903
rect 1061 20847 1181 20897
rect -1175 20723 1181 20847
rect -1175 20673 -1065 20723
rect -1519 20667 -1065 20673
rect -1009 20667 -545 20723
rect -489 20667 -25 20723
rect 31 20667 485 20723
rect 541 20667 1005 20723
rect 1061 20673 1181 20723
rect 1405 20847 1515 20897
rect 1571 20847 1838 20903
rect 1405 20723 1838 20847
rect 1405 20673 1515 20723
rect 1061 20667 1515 20673
rect 1571 20667 1838 20723
rect -1842 20650 1838 20667
rect -132 20467 138 20485
rect -132 20243 -109 20467
rect 115 20243 138 20467
rect -132 20225 138 20243
rect -3280 19690 3220 19700
rect -3280 19670 -2210 19690
rect -3280 19450 -3250 19670
rect -3030 19450 -2210 19670
rect -3280 19430 -2210 19450
rect -1950 19430 -750 19690
rect -490 19430 470 19690
rect 730 19430 1950 19690
rect 2210 19430 2950 19690
rect 3210 19430 3220 19690
rect -3280 19060 3220 19430
rect -3280 18900 -3220 19060
rect -3060 18900 -2160 19060
rect -2000 18900 -700 19060
rect -540 18900 520 19060
rect 680 18900 2000 19060
rect 2160 18900 3000 19060
rect 3160 18900 3220 19060
rect -3280 18880 3220 18900
rect -3310 17680 3310 17720
rect -3310 17570 -840 17680
rect -3310 17310 -3230 17570
rect -2970 17310 -2270 17570
rect -2010 17310 -1280 17570
rect -1020 17530 -840 17570
rect -620 17530 -320 17680
rect -100 17530 100 17680
rect 320 17530 650 17680
rect 870 17570 3310 17680
rect 870 17530 960 17570
rect -1020 17310 960 17530
rect 1220 17310 1980 17570
rect 2240 17310 2970 17570
rect 3230 17310 3310 17570
rect -3310 17130 3310 17310
rect -3310 17120 -1080 17130
rect -3310 16990 -3200 17120
rect -3020 16990 -2060 17120
rect -1880 17000 -1080 17120
rect -900 17000 -310 17130
rect -130 17000 130 17130
rect 310 17120 1920 17130
rect 310 17000 850 17120
rect -1880 16990 850 17000
rect 1030 17000 1920 17120
rect 2100 17000 2920 17130
rect 3100 17000 3310 17130
rect 1030 16990 3310 17000
rect -3310 16960 3310 16990
rect -3310 15220 -2990 16960
rect -3310 15100 -3240 15220
rect -3120 15100 -2990 15220
rect -3310 12220 -2990 15100
rect -3310 12100 -3240 12220
rect -3120 12100 -2990 12220
rect -3310 9220 -2990 12100
rect -3310 9100 -3240 9220
rect -3120 9100 -2990 9220
rect -3310 6220 -2990 9100
rect -3310 6100 -3240 6220
rect -3120 6100 -2990 6220
rect -3310 3220 -2990 6100
rect -3310 3100 -3240 3220
rect -3120 3100 -2990 3220
rect -3310 1920 -2990 3100
rect 2990 15220 3310 16960
rect 2990 15100 3130 15220
rect 3250 15100 3310 15220
rect 2990 12220 3310 15100
rect 2990 12100 3130 12220
rect 3250 12100 3310 12220
rect 2990 9220 3310 12100
rect 2990 9100 3130 9220
rect 3250 9100 3310 9220
rect 2990 6220 3310 9100
rect 2990 6100 3130 6220
rect 3250 6100 3310 6220
rect 2990 3220 3310 6100
rect 2990 3100 3130 3220
rect 3250 3100 3310 3220
rect 2990 1920 3310 3100
rect -3310 1900 3310 1920
rect -3310 1890 1690 1900
rect -3310 1480 -2860 1890
rect -1690 1480 -1350 1890
rect -180 1480 170 1890
rect 1340 1490 1690 1890
rect 2860 1490 3310 1900
rect 1340 1480 3310 1490
rect -3310 1440 3310 1480
<< via3 >>
rect -7902 36930 -7832 37000
rect -7802 36930 -7732 37000
rect 7998 36930 8068 37000
rect 8098 36930 8168 37000
rect -7902 36800 -7832 36870
rect -7802 36800 -7732 36870
rect -7374 36805 -7310 36869
rect -7294 36805 -7230 36869
rect -7214 36805 -7150 36869
rect -7134 36805 -7070 36869
rect -7054 36805 -6990 36869
rect -6974 36805 -6910 36869
rect -6894 36805 -6830 36869
rect -6814 36805 -6750 36869
rect -6734 36805 -6670 36869
rect -6654 36805 -6590 36869
rect -6574 36805 -6510 36869
rect -6494 36805 -6430 36869
rect -6414 36805 -6350 36869
rect -6334 36805 -6270 36869
rect -6254 36805 -6190 36869
rect -6174 36805 -6110 36869
rect -6094 36805 -6030 36869
rect -6014 36805 -5950 36869
rect -5934 36805 -5870 36869
rect -5854 36805 -5790 36869
rect -5774 36805 -5710 36869
rect -5694 36805 -5630 36869
rect -5614 36805 -5550 36869
rect -5534 36805 -5470 36869
rect -5454 36805 -5390 36869
rect -5374 36805 -5310 36869
rect -5294 36805 -5230 36869
rect -5214 36805 -5150 36869
rect -5134 36805 -5070 36869
rect -5054 36805 -4990 36869
rect -4974 36805 -4910 36869
rect -4894 36805 -4830 36869
rect -4814 36805 -4750 36869
rect -4734 36805 -4670 36869
rect -4654 36805 -4590 36869
rect -4574 36805 -4510 36869
rect -4494 36805 -4430 36869
rect -4414 36805 -4350 36869
rect -4334 36805 -4270 36869
rect -4254 36805 -4190 36869
rect -4174 36805 -4110 36869
rect -4094 36805 -4030 36869
rect -3574 36805 -3510 36869
rect -3494 36805 -3430 36869
rect -3414 36805 -3350 36869
rect -3334 36805 -3270 36869
rect -3254 36805 -3190 36869
rect -3174 36805 -3110 36869
rect -3094 36805 -3030 36869
rect -3014 36805 -2950 36869
rect -2934 36805 -2870 36869
rect -2854 36805 -2790 36869
rect -2774 36805 -2710 36869
rect -2694 36805 -2630 36869
rect -2614 36805 -2550 36869
rect -2534 36805 -2470 36869
rect -2454 36805 -2390 36869
rect -2374 36805 -2310 36869
rect -2294 36805 -2230 36869
rect -2214 36805 -2150 36869
rect -2134 36805 -2070 36869
rect -2054 36805 -1990 36869
rect -1974 36805 -1910 36869
rect -1894 36805 -1830 36869
rect -1814 36805 -1750 36869
rect -1734 36805 -1670 36869
rect -1654 36805 -1590 36869
rect -1574 36805 -1510 36869
rect -1494 36805 -1430 36869
rect -1414 36805 -1350 36869
rect -1334 36805 -1270 36869
rect -1254 36805 -1190 36869
rect -1174 36805 -1110 36869
rect -1094 36805 -1030 36869
rect -1014 36805 -950 36869
rect -934 36805 -870 36869
rect -854 36805 -790 36869
rect -774 36805 -710 36869
rect -694 36805 -630 36869
rect -614 36805 -550 36869
rect -534 36805 -470 36869
rect -454 36805 -390 36869
rect -374 36805 -310 36869
rect -294 36805 -230 36869
rect 226 36805 290 36869
rect 306 36805 370 36869
rect 386 36805 450 36869
rect 466 36805 530 36869
rect 546 36805 610 36869
rect 626 36805 690 36869
rect 706 36805 770 36869
rect 786 36805 850 36869
rect 866 36805 930 36869
rect 946 36805 1010 36869
rect 1026 36805 1090 36869
rect 1106 36805 1170 36869
rect 1186 36805 1250 36869
rect 1266 36805 1330 36869
rect 1346 36805 1410 36869
rect 1426 36805 1490 36869
rect 1506 36805 1570 36869
rect 1586 36805 1650 36869
rect 1666 36805 1730 36869
rect 1746 36805 1810 36869
rect 1826 36805 1890 36869
rect 1906 36805 1970 36869
rect 1986 36805 2050 36869
rect 2066 36805 2130 36869
rect 2146 36805 2210 36869
rect 2226 36805 2290 36869
rect 2306 36805 2370 36869
rect 2386 36805 2450 36869
rect 2466 36805 2530 36869
rect 2546 36805 2610 36869
rect 2626 36805 2690 36869
rect 2706 36805 2770 36869
rect 2786 36805 2850 36869
rect 2866 36805 2930 36869
rect 2946 36805 3010 36869
rect 3026 36805 3090 36869
rect 3106 36805 3170 36869
rect 3186 36805 3250 36869
rect 3266 36805 3330 36869
rect 3346 36805 3410 36869
rect 3426 36805 3490 36869
rect 3506 36805 3570 36869
rect 4026 36805 4090 36869
rect 4106 36805 4170 36869
rect 4186 36805 4250 36869
rect 4266 36805 4330 36869
rect 4346 36805 4410 36869
rect 4426 36805 4490 36869
rect 4506 36805 4570 36869
rect 4586 36805 4650 36869
rect 4666 36805 4730 36869
rect 4746 36805 4810 36869
rect 4826 36805 4890 36869
rect 4906 36805 4970 36869
rect 4986 36805 5050 36869
rect 5066 36805 5130 36869
rect 5146 36805 5210 36869
rect 5226 36805 5290 36869
rect 5306 36805 5370 36869
rect 5386 36805 5450 36869
rect 5466 36805 5530 36869
rect 5546 36805 5610 36869
rect 5626 36805 5690 36869
rect 5706 36805 5770 36869
rect 5786 36805 5850 36869
rect 5866 36805 5930 36869
rect 5946 36805 6010 36869
rect 6026 36805 6090 36869
rect 6106 36805 6170 36869
rect 6186 36805 6250 36869
rect 6266 36805 6330 36869
rect 6346 36805 6410 36869
rect 6426 36805 6490 36869
rect 6506 36805 6570 36869
rect 6586 36805 6650 36869
rect 6666 36805 6730 36869
rect 6746 36805 6810 36869
rect 6826 36805 6890 36869
rect 6906 36805 6970 36869
rect 6986 36805 7050 36869
rect 7066 36805 7130 36869
rect 7146 36805 7210 36869
rect 7226 36805 7290 36869
rect 7306 36805 7370 36869
rect 7998 36800 8068 36870
rect 8098 36800 8168 36870
rect -619 31373 -395 31377
rect -619 31157 -615 31373
rect -615 31157 -399 31373
rect -399 31157 -395 31373
rect -619 31153 -395 31157
rect 431 31373 655 31377
rect 431 31157 435 31373
rect 435 31157 651 31373
rect 651 31157 655 31373
rect 431 31153 655 31157
rect -2799 30663 -2575 30887
rect -899 30653 -675 30877
rect 681 30653 905 30877
rect 2581 30653 2805 30877
rect -3669 29633 -3605 29697
rect -619 29733 -395 29737
rect -619 29517 -615 29733
rect -615 29517 -399 29733
rect -399 29517 -395 29733
rect -619 29513 -395 29517
rect 431 29733 655 29737
rect 431 29517 435 29733
rect 435 29517 651 29733
rect 651 29517 655 29733
rect 431 29513 655 29517
rect 3381 29633 3445 29697
rect -1294 28998 -1070 29222
rect -24 28998 200 29222
rect 1236 28998 1460 29222
rect -854 28128 -630 28132
rect -854 27912 -850 28128
rect -850 27912 -634 28128
rect -634 27912 -630 28128
rect -854 27908 -630 27912
rect 646 28128 870 28132
rect 646 27912 650 28128
rect 650 27912 866 28128
rect 866 27912 870 28128
rect 646 27908 870 27912
rect -1294 27448 -1070 27672
rect -24 27448 200 27672
rect 1236 27448 1460 27672
rect -114 25028 110 25032
rect -114 24812 -110 25028
rect -110 24812 106 25028
rect 106 24812 110 25028
rect -114 24808 110 24812
rect -114 23508 110 23512
rect -114 23292 -110 23508
rect -110 23292 106 23508
rect 106 23292 110 23508
rect -114 23288 110 23292
rect -1139 22193 -915 22417
rect 921 22193 1145 22417
rect -109 21993 115 21997
rect -109 21777 -105 21993
rect -105 21777 111 21993
rect 111 21777 115 21993
rect -109 21773 115 21777
rect -3239 21718 -2695 21722
rect -3239 21342 -3235 21718
rect -3235 21342 -2699 21718
rect -2699 21342 -2695 21718
rect -3239 21338 -2695 21342
rect 2638 21440 2878 21680
rect 2968 21440 3208 21680
rect -1399 20673 -1175 20897
rect 1181 20673 1405 20897
rect -109 20463 115 20467
rect -109 20247 -105 20463
rect -105 20247 111 20463
rect 111 20247 115 20463
rect -109 20243 115 20247
rect -3250 19640 -3030 19670
rect -3250 19480 -3220 19640
rect -3220 19480 -3060 19640
rect -3060 19480 -3030 19640
rect -3250 19450 -3030 19480
rect -2210 19640 -1950 19690
rect -2210 19480 -2160 19640
rect -2160 19480 -2000 19640
rect -2000 19480 -1950 19640
rect -2210 19430 -1950 19480
rect -750 19640 -490 19690
rect -750 19480 -700 19640
rect -700 19480 -540 19640
rect -540 19480 -490 19640
rect -750 19430 -490 19480
rect 470 19640 730 19690
rect 470 19480 520 19640
rect 520 19480 680 19640
rect 680 19480 730 19640
rect 470 19430 730 19480
rect 1950 19640 2210 19690
rect 1950 19480 2000 19640
rect 2000 19480 2160 19640
rect 2160 19480 2210 19640
rect 1950 19430 2210 19480
rect 2950 19640 3210 19690
rect 2950 19480 3000 19640
rect 3000 19480 3160 19640
rect 3160 19480 3210 19640
rect 2950 19430 3210 19480
rect -3230 17310 -2970 17570
rect -2270 17310 -2010 17570
rect -1280 17310 -1020 17570
rect 960 17310 1220 17570
rect 1980 17310 2240 17570
rect 2970 17310 3230 17570
<< mimcap >>
rect -7302 36642 -4102 36690
rect -7302 33538 -7254 36642
rect -4150 33538 -4102 36642
rect -7302 33490 -4102 33538
rect -3502 36642 -302 36690
rect -3502 33538 -3454 36642
rect -350 33538 -302 36642
rect -3502 33490 -302 33538
rect 298 36642 3498 36690
rect 298 33538 346 36642
rect 3450 33538 3498 36642
rect 298 33490 3498 33538
rect 4098 36642 7298 36690
rect 4098 33538 4146 36642
rect 7250 33538 7298 36642
rect 4098 33490 7298 33538
<< mimcapcontact >>
rect -7254 33538 -4150 36642
rect -3454 33538 -350 36642
rect 346 33538 3450 36642
rect 4146 33538 7250 36642
<< metal4 >>
rect -7922 37000 8188 37020
rect -7922 36930 -7902 37000
rect -7832 36930 -7802 37000
rect -7732 36930 7998 37000
rect 8068 36930 8098 37000
rect 8168 36930 8188 37000
rect -7922 36870 8188 36930
rect -7922 36800 -7902 36870
rect -7832 36800 -7802 36870
rect -7732 36869 7998 36870
rect -7732 36805 -7374 36869
rect -7310 36805 -7294 36869
rect -7230 36805 -7214 36869
rect -7150 36805 -7134 36869
rect -7070 36805 -7054 36869
rect -6990 36805 -6974 36869
rect -6910 36805 -6894 36869
rect -6830 36805 -6814 36869
rect -6750 36805 -6734 36869
rect -6670 36805 -6654 36869
rect -6590 36805 -6574 36869
rect -6510 36805 -6494 36869
rect -6430 36805 -6414 36869
rect -6350 36805 -6334 36869
rect -6270 36805 -6254 36869
rect -6190 36805 -6174 36869
rect -6110 36805 -6094 36869
rect -6030 36805 -6014 36869
rect -5950 36805 -5934 36869
rect -5870 36805 -5854 36869
rect -5790 36805 -5774 36869
rect -5710 36805 -5694 36869
rect -5630 36805 -5614 36869
rect -5550 36805 -5534 36869
rect -5470 36805 -5454 36869
rect -5390 36805 -5374 36869
rect -5310 36805 -5294 36869
rect -5230 36805 -5214 36869
rect -5150 36805 -5134 36869
rect -5070 36805 -5054 36869
rect -4990 36805 -4974 36869
rect -4910 36805 -4894 36869
rect -4830 36805 -4814 36869
rect -4750 36805 -4734 36869
rect -4670 36805 -4654 36869
rect -4590 36805 -4574 36869
rect -4510 36805 -4494 36869
rect -4430 36805 -4414 36869
rect -4350 36805 -4334 36869
rect -4270 36805 -4254 36869
rect -4190 36805 -4174 36869
rect -4110 36805 -4094 36869
rect -4030 36805 -3574 36869
rect -3510 36805 -3494 36869
rect -3430 36805 -3414 36869
rect -3350 36805 -3334 36869
rect -3270 36805 -3254 36869
rect -3190 36805 -3174 36869
rect -3110 36805 -3094 36869
rect -3030 36805 -3014 36869
rect -2950 36805 -2934 36869
rect -2870 36805 -2854 36869
rect -2790 36805 -2774 36869
rect -2710 36805 -2694 36869
rect -2630 36805 -2614 36869
rect -2550 36805 -2534 36869
rect -2470 36805 -2454 36869
rect -2390 36805 -2374 36869
rect -2310 36805 -2294 36869
rect -2230 36805 -2214 36869
rect -2150 36805 -2134 36869
rect -2070 36805 -2054 36869
rect -1990 36805 -1974 36869
rect -1910 36805 -1894 36869
rect -1830 36805 -1814 36869
rect -1750 36805 -1734 36869
rect -1670 36805 -1654 36869
rect -1590 36805 -1574 36869
rect -1510 36805 -1494 36869
rect -1430 36805 -1414 36869
rect -1350 36805 -1334 36869
rect -1270 36805 -1254 36869
rect -1190 36805 -1174 36869
rect -1110 36805 -1094 36869
rect -1030 36805 -1014 36869
rect -950 36805 -934 36869
rect -870 36805 -854 36869
rect -790 36805 -774 36869
rect -710 36805 -694 36869
rect -630 36805 -614 36869
rect -550 36805 -534 36869
rect -470 36805 -454 36869
rect -390 36805 -374 36869
rect -310 36805 -294 36869
rect -230 36805 226 36869
rect 290 36805 306 36869
rect 370 36805 386 36869
rect 450 36805 466 36869
rect 530 36805 546 36869
rect 610 36805 626 36869
rect 690 36805 706 36869
rect 770 36805 786 36869
rect 850 36805 866 36869
rect 930 36805 946 36869
rect 1010 36805 1026 36869
rect 1090 36805 1106 36869
rect 1170 36805 1186 36869
rect 1250 36805 1266 36869
rect 1330 36805 1346 36869
rect 1410 36805 1426 36869
rect 1490 36805 1506 36869
rect 1570 36805 1586 36869
rect 1650 36805 1666 36869
rect 1730 36805 1746 36869
rect 1810 36805 1826 36869
rect 1890 36805 1906 36869
rect 1970 36805 1986 36869
rect 2050 36805 2066 36869
rect 2130 36805 2146 36869
rect 2210 36805 2226 36869
rect 2290 36805 2306 36869
rect 2370 36805 2386 36869
rect 2450 36805 2466 36869
rect 2530 36805 2546 36869
rect 2610 36805 2626 36869
rect 2690 36805 2706 36869
rect 2770 36805 2786 36869
rect 2850 36805 2866 36869
rect 2930 36805 2946 36869
rect 3010 36805 3026 36869
rect 3090 36805 3106 36869
rect 3170 36805 3186 36869
rect 3250 36805 3266 36869
rect 3330 36805 3346 36869
rect 3410 36805 3426 36869
rect 3490 36805 3506 36869
rect 3570 36805 4026 36869
rect 4090 36805 4106 36869
rect 4170 36805 4186 36869
rect 4250 36805 4266 36869
rect 4330 36805 4346 36869
rect 4410 36805 4426 36869
rect 4490 36805 4506 36869
rect 4570 36805 4586 36869
rect 4650 36805 4666 36869
rect 4730 36805 4746 36869
rect 4810 36805 4826 36869
rect 4890 36805 4906 36869
rect 4970 36805 4986 36869
rect 5050 36805 5066 36869
rect 5130 36805 5146 36869
rect 5210 36805 5226 36869
rect 5290 36805 5306 36869
rect 5370 36805 5386 36869
rect 5450 36805 5466 36869
rect 5530 36805 5546 36869
rect 5610 36805 5626 36869
rect 5690 36805 5706 36869
rect 5770 36805 5786 36869
rect 5850 36805 5866 36869
rect 5930 36805 5946 36869
rect 6010 36805 6026 36869
rect 6090 36805 6106 36869
rect 6170 36805 6186 36869
rect 6250 36805 6266 36869
rect 6330 36805 6346 36869
rect 6410 36805 6426 36869
rect 6490 36805 6506 36869
rect 6570 36805 6586 36869
rect 6650 36805 6666 36869
rect 6730 36805 6746 36869
rect 6810 36805 6826 36869
rect 6890 36805 6906 36869
rect 6970 36805 6986 36869
rect 7050 36805 7066 36869
rect 7130 36805 7146 36869
rect 7210 36805 7226 36869
rect 7290 36805 7306 36869
rect 7370 36805 7998 36869
rect -7732 36800 7998 36805
rect 8068 36800 8098 36870
rect 8168 36800 8188 36870
rect -7922 36780 8188 36800
rect -7263 36642 -4141 36651
rect -7263 33538 -7254 36642
rect -4150 35310 -4141 36642
rect -3463 36642 -341 36651
rect -3463 35310 -3454 36642
rect -4150 34950 -3454 35310
rect -4150 33538 -4141 34950
rect -7263 33529 -4141 33538
rect -3962 32162 -3642 34950
rect -3463 33538 -3454 34950
rect -350 35310 -341 36642
rect 337 36642 3459 36651
rect 337 35310 346 36642
rect -350 34950 346 35310
rect -350 33538 -341 34950
rect -3463 33529 -341 33538
rect 337 33538 346 34950
rect 3450 35310 3459 36642
rect 4137 36642 7259 36651
rect 4137 35310 4146 36642
rect 3450 34950 4146 35310
rect 3450 33538 3459 34950
rect 337 33529 3459 33538
rect -10700 31400 -9200 31500
rect -10700 31100 -10600 31400
rect -10300 31100 -9600 31400
rect -9300 31100 -9200 31400
rect -10700 30700 -9200 31100
rect -10700 30400 -10600 30700
rect -10300 30400 -9600 30700
rect -9300 30400 -9200 30700
rect -10700 28400 -9200 30400
rect -3960 29730 -3642 32162
rect -643 31383 -371 31401
rect -643 31147 -625 31383
rect -389 31147 -371 31383
rect -643 31129 -371 31147
rect 407 31383 679 31401
rect 407 31147 425 31383
rect 661 31147 679 31383
rect 407 31129 679 31147
rect -2813 30893 -2561 30901
rect -2813 30657 -2805 30893
rect -2569 30657 -2561 30893
rect -2813 30649 -2561 30657
rect -913 30883 -661 30891
rect -913 30647 -905 30883
rect -669 30647 -661 30883
rect -913 30639 -661 30647
rect 667 30883 919 30891
rect 667 30647 675 30883
rect 911 30647 919 30883
rect 667 30639 919 30647
rect 2567 30883 2819 30891
rect 2567 30647 2575 30883
rect 2811 30647 2819 30883
rect 2567 30639 2819 30647
rect -643 29743 -371 29761
rect -3960 29697 -3562 29730
rect -3960 29633 -3669 29697
rect -3605 29633 -3562 29697
rect -3960 29600 -3562 29633
rect -643 29507 -625 29743
rect -389 29507 -371 29743
rect -643 29489 -371 29507
rect 407 29743 679 29761
rect 407 29507 425 29743
rect 661 29507 679 29743
rect 3648 29730 3968 34950
rect 4137 33538 4146 34950
rect 7250 33538 7259 36642
rect 4137 33529 7259 33538
rect 3338 29697 3968 29730
rect 3338 29633 3381 29697
rect 3445 29633 3968 29697
rect 3338 29600 3968 29633
rect 407 29489 679 29507
rect -1313 29228 -1051 29241
rect -1313 28992 -1300 29228
rect -1064 28992 -1051 29228
rect -1313 28979 -1051 28992
rect -43 29228 219 29241
rect -43 28992 -30 29228
rect 206 28992 219 29228
rect -43 28979 219 28992
rect 1217 29228 1479 29241
rect 1217 28992 1230 29228
rect 1466 28992 1479 29228
rect 1217 28979 1479 28992
rect -10700 28100 -10600 28400
rect -10300 28100 -9600 28400
rect -9300 28100 -9200 28400
rect -10700 27800 -9200 28100
rect -873 28138 -611 28151
rect -873 27902 -860 28138
rect -624 27902 -611 28138
rect -873 27889 -611 27902
rect 627 28138 889 28151
rect 627 27902 640 28138
rect 876 27902 889 28138
rect 627 27889 889 27902
rect -10700 27500 -10600 27800
rect -10300 27500 -9600 27800
rect -9300 27500 -9200 27800
rect -10700 19700 -9200 27500
rect -1313 27678 -1051 27691
rect -1313 27442 -1300 27678
rect -1064 27442 -1051 27678
rect -1313 27429 -1051 27442
rect -43 27678 219 27691
rect -43 27442 -30 27678
rect 206 27442 219 27678
rect -43 27429 219 27442
rect 1217 27678 1479 27691
rect 1217 27442 1230 27678
rect 1466 27442 1479 27678
rect 1217 27429 1479 27442
rect -133 25038 129 25051
rect -133 24802 -120 25038
rect 116 24802 129 25038
rect -133 24789 129 24802
rect -133 23518 129 23531
rect -133 23282 -120 23518
rect 116 23282 129 23518
rect -133 23269 129 23282
rect -1153 22423 -901 22431
rect -1153 22187 -1145 22423
rect -909 22187 -901 22423
rect -1153 22179 -901 22187
rect 907 22423 1159 22431
rect 907 22187 915 22423
rect 1151 22187 1159 22423
rect 907 22179 1159 22187
rect 7600 22400 9100 22500
rect 7600 22100 7700 22400
rect 8000 22100 8700 22400
rect 9000 22100 9100 22400
rect -123 22003 129 22011
rect -123 21767 -115 22003
rect 121 21767 129 22003
rect -123 21759 129 21767
rect -3263 21722 -2671 21741
rect -3263 21648 -3239 21722
rect -2695 21648 -2671 21722
rect 7600 21700 9100 22100
rect -3263 21412 -3245 21648
rect -2689 21412 -2671 21648
rect 2637 21680 2879 21681
rect 2637 21440 2638 21680
rect 2878 21440 2879 21680
rect 2637 21439 2879 21440
rect 2967 21680 3209 21681
rect 2967 21440 2968 21680
rect 3208 21440 3209 21680
rect 2967 21439 3209 21440
rect -3263 21338 -3239 21412
rect -2695 21338 -2671 21412
rect -3263 21319 -2671 21338
rect 7600 21400 7700 21700
rect 8000 21400 8700 21700
rect 9000 21400 9100 21700
rect 7600 21000 9100 21400
rect -1413 20903 -1161 20911
rect -1413 20667 -1405 20903
rect -1169 20667 -1161 20903
rect -1413 20659 -1161 20667
rect 1167 20903 1419 20911
rect 1167 20667 1175 20903
rect 1411 20667 1419 20903
rect 1167 20659 1419 20667
rect 7600 20700 7700 21000
rect 8000 20700 8700 21000
rect 9000 20700 9100 21000
rect -123 20473 129 20481
rect -123 20237 -115 20473
rect 121 20237 129 20473
rect -123 20229 129 20237
rect -10700 19400 -10600 19700
rect -10300 19400 -9600 19700
rect -9300 19400 -9200 19700
rect -2211 19690 -1949 19691
rect -2211 19430 -2210 19690
rect -1950 19430 -1949 19690
rect -2211 19429 -1949 19430
rect -751 19690 -489 19691
rect -751 19430 -750 19690
rect -490 19430 -489 19690
rect -751 19429 -489 19430
rect 469 19690 731 19691
rect 469 19430 470 19690
rect 730 19430 731 19690
rect 469 19429 731 19430
rect 1949 19690 2211 19691
rect 1949 19430 1950 19690
rect 2210 19430 2211 19690
rect 1949 19429 2211 19430
rect 2949 19690 3211 19691
rect 2949 19430 2950 19690
rect 3210 19430 3211 19690
rect 2949 19429 3211 19430
rect -10700 19200 -9200 19400
rect -10700 18900 -10600 19200
rect -10300 18900 -9600 19200
rect -9300 18900 -9200 19200
rect -10700 18800 -9200 18900
rect 7600 17700 9100 20700
rect -3231 17570 -2969 17571
rect -3231 17310 -3230 17570
rect -2970 17310 -2969 17570
rect -3231 17309 -2969 17310
rect -2271 17570 -2009 17571
rect -2271 17310 -2270 17570
rect -2010 17310 -2009 17570
rect -2271 17309 -2009 17310
rect -1281 17570 -1019 17571
rect -1281 17310 -1280 17570
rect -1020 17310 -1019 17570
rect -1281 17309 -1019 17310
rect 959 17570 1221 17571
rect 959 17310 960 17570
rect 1220 17310 1221 17570
rect 959 17309 1221 17310
rect 1979 17570 2241 17571
rect 1979 17310 1980 17570
rect 2240 17310 2241 17570
rect 1979 17309 2241 17310
rect 2969 17570 3231 17571
rect 2969 17310 2970 17570
rect 3230 17310 3231 17570
rect 2969 17309 3231 17310
rect 7600 17400 7700 17700
rect 8000 17400 8700 17700
rect 9000 17400 9100 17700
rect 7600 17200 9100 17400
rect 7600 16900 7700 17200
rect 8000 16900 8700 17200
rect 9000 16900 9100 17200
rect 7600 16800 9100 16900
<< via4 >>
rect -10600 31100 -10300 31400
rect -9600 31100 -9300 31400
rect -10600 30400 -10300 30700
rect -9600 30400 -9300 30700
rect -625 31377 -389 31383
rect -625 31153 -619 31377
rect -619 31153 -395 31377
rect -395 31153 -389 31377
rect -625 31147 -389 31153
rect 425 31377 661 31383
rect 425 31153 431 31377
rect 431 31153 655 31377
rect 655 31153 661 31377
rect 425 31147 661 31153
rect -2805 30887 -2569 30893
rect -2805 30663 -2799 30887
rect -2799 30663 -2575 30887
rect -2575 30663 -2569 30887
rect -2805 30657 -2569 30663
rect -905 30877 -669 30883
rect -905 30653 -899 30877
rect -899 30653 -675 30877
rect -675 30653 -669 30877
rect -905 30647 -669 30653
rect 675 30877 911 30883
rect 675 30653 681 30877
rect 681 30653 905 30877
rect 905 30653 911 30877
rect 675 30647 911 30653
rect 2575 30877 2811 30883
rect 2575 30653 2581 30877
rect 2581 30653 2805 30877
rect 2805 30653 2811 30877
rect 2575 30647 2811 30653
rect -625 29737 -389 29743
rect -625 29513 -619 29737
rect -619 29513 -395 29737
rect -395 29513 -389 29737
rect -625 29507 -389 29513
rect 425 29737 661 29743
rect 425 29513 431 29737
rect 431 29513 655 29737
rect 655 29513 661 29737
rect 425 29507 661 29513
rect -1300 29222 -1064 29228
rect -1300 28998 -1294 29222
rect -1294 28998 -1070 29222
rect -1070 28998 -1064 29222
rect -1300 28992 -1064 28998
rect -30 29222 206 29228
rect -30 28998 -24 29222
rect -24 28998 200 29222
rect 200 28998 206 29222
rect -30 28992 206 28998
rect 1230 29222 1466 29228
rect 1230 28998 1236 29222
rect 1236 28998 1460 29222
rect 1460 28998 1466 29222
rect 1230 28992 1466 28998
rect -10600 28100 -10300 28400
rect -9600 28100 -9300 28400
rect -860 28132 -624 28138
rect -860 27908 -854 28132
rect -854 27908 -630 28132
rect -630 27908 -624 28132
rect -860 27902 -624 27908
rect 640 28132 876 28138
rect 640 27908 646 28132
rect 646 27908 870 28132
rect 870 27908 876 28132
rect 640 27902 876 27908
rect -10600 27500 -10300 27800
rect -9600 27500 -9300 27800
rect -1300 27672 -1064 27678
rect -1300 27448 -1294 27672
rect -1294 27448 -1070 27672
rect -1070 27448 -1064 27672
rect -1300 27442 -1064 27448
rect -30 27672 206 27678
rect -30 27448 -24 27672
rect -24 27448 200 27672
rect 200 27448 206 27672
rect -30 27442 206 27448
rect 1230 27672 1466 27678
rect 1230 27448 1236 27672
rect 1236 27448 1460 27672
rect 1460 27448 1466 27672
rect 1230 27442 1466 27448
rect -120 25032 116 25038
rect -120 24808 -114 25032
rect -114 24808 110 25032
rect 110 24808 116 25032
rect -120 24802 116 24808
rect -120 23512 116 23518
rect -120 23288 -114 23512
rect -114 23288 110 23512
rect 110 23288 116 23512
rect -120 23282 116 23288
rect -1145 22417 -909 22423
rect -1145 22193 -1139 22417
rect -1139 22193 -915 22417
rect -915 22193 -909 22417
rect -1145 22187 -909 22193
rect 915 22417 1151 22423
rect 915 22193 921 22417
rect 921 22193 1145 22417
rect 1145 22193 1151 22417
rect 915 22187 1151 22193
rect 7700 22100 8000 22400
rect 8700 22100 9000 22400
rect -115 21997 121 22003
rect -115 21773 -109 21997
rect -109 21773 115 21997
rect 115 21773 121 21997
rect -115 21767 121 21773
rect -3245 21412 -3239 21648
rect -3239 21412 -3009 21648
rect -2925 21412 -2695 21648
rect -2695 21412 -2689 21648
rect 2638 21440 2878 21680
rect 2968 21440 3208 21680
rect 7700 21400 8000 21700
rect 8700 21400 9000 21700
rect -1405 20897 -1169 20903
rect -1405 20673 -1399 20897
rect -1399 20673 -1175 20897
rect -1175 20673 -1169 20897
rect -1405 20667 -1169 20673
rect 1175 20897 1411 20903
rect 1175 20673 1181 20897
rect 1181 20673 1405 20897
rect 1405 20673 1411 20897
rect 1175 20667 1411 20673
rect 7700 20700 8000 21000
rect 8700 20700 9000 21000
rect -115 20467 121 20473
rect -115 20243 -109 20467
rect -109 20243 115 20467
rect 115 20243 121 20467
rect -115 20237 121 20243
rect -10600 19400 -10300 19700
rect -9600 19400 -9300 19700
rect -3270 19670 -3010 19690
rect -3270 19450 -3250 19670
rect -3250 19450 -3030 19670
rect -3030 19450 -3010 19670
rect -3270 19430 -3010 19450
rect -2210 19430 -1950 19690
rect -750 19430 -490 19690
rect 470 19430 730 19690
rect 1950 19430 2210 19690
rect 2950 19430 3210 19690
rect -10600 18900 -10300 19200
rect -9600 18900 -9300 19200
rect -3230 17310 -2970 17570
rect -2270 17310 -2010 17570
rect -1280 17310 -1020 17570
rect 960 17310 1220 17570
rect 1980 17310 2240 17570
rect 2970 17310 3230 17570
rect 7700 17400 8000 17700
rect 8700 17400 9000 17700
rect 7700 16900 8000 17200
rect 8700 16900 9000 17200
<< metal5 >>
rect -10700 31400 9100 31500
rect -10700 31100 -10600 31400
rect -10300 31100 -9600 31400
rect -9300 31383 9100 31400
rect -9300 31147 -625 31383
rect -389 31147 425 31383
rect 661 31147 9100 31383
rect -9300 31100 9100 31147
rect -10700 30893 9100 31100
rect -10700 30700 -2805 30893
rect -10700 30400 -10600 30700
rect -10300 30400 -9600 30700
rect -9300 30657 -2805 30700
rect -2569 30883 9100 30893
rect -2569 30657 -905 30883
rect -9300 30647 -905 30657
rect -669 30647 675 30883
rect 911 30647 2575 30883
rect 2811 30647 9100 30883
rect -9300 30400 9100 30647
rect -10700 29743 9100 30400
rect -10700 29507 -625 29743
rect -389 29507 425 29743
rect 661 29507 9100 29743
rect -10700 29228 9100 29507
rect -10700 28992 -1300 29228
rect -1064 28992 -30 29228
rect 206 28992 1230 29228
rect 1466 28992 9100 29228
rect -10700 28400 9100 28992
rect -10700 28100 -10600 28400
rect -10300 28100 -9600 28400
rect -9300 28138 9100 28400
rect -9300 28100 -860 28138
rect -10700 27902 -860 28100
rect -624 27902 640 28138
rect 876 27902 9100 28138
rect -10700 27800 9100 27902
rect -10700 27500 -10600 27800
rect -10300 27500 -9600 27800
rect -9300 27678 9100 27800
rect -9300 27500 -1300 27678
rect -10700 27442 -1300 27500
rect -1064 27442 -30 27678
rect 206 27442 1230 27678
rect 1466 27442 9100 27678
rect -10700 27400 9100 27442
rect -222 25038 218 25090
rect -222 24802 -120 25038
rect 116 24802 218 25038
rect -222 23518 218 24802
rect -222 23282 -120 23518
rect 116 23282 218 23518
rect -222 22500 218 23282
rect -10700 22423 9100 22500
rect -10700 22187 -1145 22423
rect -909 22187 915 22423
rect 1151 22400 9100 22423
rect 1151 22187 7700 22400
rect -10700 22100 7700 22187
rect 8000 22100 8700 22400
rect 9000 22100 9100 22400
rect -10700 22003 9100 22100
rect -10700 21767 -115 22003
rect 121 21767 9100 22003
rect -10700 21700 9100 21767
rect -10700 21680 7700 21700
rect -10700 21648 2638 21680
rect -10700 21412 -3245 21648
rect -3009 21412 -2925 21648
rect -2689 21440 2638 21648
rect 2878 21440 2968 21680
rect 3208 21440 7700 21680
rect -2689 21412 7700 21440
rect -10700 21400 7700 21412
rect 8000 21400 8700 21700
rect 9000 21400 9100 21700
rect -10700 21000 9100 21400
rect -10700 20903 7700 21000
rect -10700 20667 -1405 20903
rect -1169 20667 1175 20903
rect 1411 20700 7700 20903
rect 8000 20700 8700 21000
rect 9000 20700 9100 21000
rect 1411 20667 9100 20700
rect -10700 20600 9100 20667
rect -212 20473 228 20600
rect -212 20237 -115 20473
rect 121 20237 228 20473
rect -212 20160 228 20237
rect -10700 19700 9100 19800
rect -10700 19400 -10600 19700
rect -10300 19400 -9600 19700
rect -9300 19690 9100 19700
rect -9300 19430 -3270 19690
rect -3010 19430 -2210 19690
rect -1950 19430 -750 19690
rect -490 19430 470 19690
rect 730 19430 1950 19690
rect 2210 19430 2950 19690
rect 3210 19430 9100 19690
rect -9300 19400 9100 19430
rect -10700 19200 9100 19400
rect -10700 18900 -10600 19200
rect -10300 18900 -9600 19200
rect -9300 18900 9100 19200
rect -10700 18800 9100 18900
rect -10700 17700 9100 17800
rect -10700 17570 7700 17700
rect -10700 17310 -3230 17570
rect -2970 17310 -2270 17570
rect -2010 17310 -1280 17570
rect -1020 17310 960 17570
rect 1220 17310 1980 17570
rect 2240 17310 2970 17570
rect 3230 17400 7700 17570
rect 8000 17400 8700 17700
rect 9000 17400 9100 17700
rect 3230 17310 9100 17400
rect -10700 17200 9100 17310
rect -10700 16900 7700 17200
rect 8000 16900 8700 17200
rect 9000 16900 9100 17200
rect -10700 16800 9100 16900
<< res5p73 >>
rect -6704 30794 -4700 31944
rect -6704 29294 -4700 30444
rect -2845 1930 -1695 15734
rect -1325 1930 -175 15734
rect 185 1936 1335 15740
rect 1695 1936 2845 15740
<< labels >>
rlabel metal2 880 20190 1200 20350 1 Vmirror
port 1 n
rlabel metal1 -3580 30390 -3420 30560 1 Vmid
port 2 n
rlabel metal4 3700 30810 3920 31170 1 Vout
port 3 n
rlabel metal1 710 25600 760 25760 1 Vp
port 4 n
rlabel metal1 710 24080 760 24240 1 Vn
port 5 n
rlabel metal5 -8800 27800 -7600 28400 1 Vdd
port 6 n
rlabel metal5 -8400 20900 -7300 21600 1 Vss
port 7 n
<< end >>
