magic
tech sky130A
magscale 1 2
timestamp 1679690840
<< metal1 >>
rect 3844 30396 4126 30622
rect 1738 28844 1816 29002
rect 690 25652 770 25778
rect 690 24160 770 24230
<< metal2 >>
rect -2420 20370 -2020 20410
rect 1980 20370 2380 20480
rect -2420 20170 -330 20370
rect -480 18830 -330 20170
rect 330 20170 2380 20370
rect 330 18830 480 20170
rect -580 18570 -360 18830
rect 360 18570 580 18830
<< metal3 >>
rect -3010 19100 -3000 19400
rect -2700 19100 -2690 19400
rect -1410 19100 -1400 19400
rect -1100 19100 -1090 19400
rect 400 19380 980 19680
rect 1090 19100 1100 19400
rect 1400 19100 1410 19400
rect 2590 19100 2600 19400
rect 2900 19100 2910 19400
rect 1260 17500 1840 17570
rect -3110 17200 -3100 17500
rect -2800 17200 -2790 17500
rect -2210 17200 -2200 17500
rect -1900 17200 -1890 17500
rect -1310 17200 -1300 17500
rect -1000 17200 -990 17500
rect 990 17200 1000 17500
rect 1300 17270 1840 17500
rect 1300 17200 1310 17270
rect 1890 17200 1900 17500
rect 2200 17200 2210 17500
rect 2790 17200 2800 17500
rect 3100 17200 3110 17500
<< via3 >>
rect -3000 19100 -2700 19400
rect -1400 19100 -1100 19400
rect 1100 19100 1400 19400
rect 2600 19100 2900 19400
rect -3100 17200 -2800 17500
rect -2200 17200 -1900 17500
rect -1300 17200 -1000 17500
rect 1000 17200 1300 17500
rect 1900 17200 2200 17500
rect 2800 17200 3100 17500
<< metal4 >>
rect 3716 32514 3902 32770
rect 6710 28340 7380 28370
rect -7450 28240 -6780 28270
rect -7450 28000 -7420 28240
rect -7180 28000 -7050 28240
rect -6810 28000 -6780 28240
rect -7450 27670 -6780 28000
rect -7450 27430 -7420 27670
rect -7180 27430 -7050 27670
rect -6810 27430 -6780 27670
rect -7450 19770 -6780 27430
rect 6710 28100 6740 28340
rect 6980 28100 7110 28340
rect 7350 28100 7380 28340
rect 6710 27670 7380 28100
rect 6710 27430 6740 27670
rect 6980 27430 7110 27670
rect 7350 27430 7380 27670
rect -7450 19530 -7420 19770
rect -7180 19530 -7050 19770
rect -6810 19530 -6780 19770
rect -7450 18570 -6780 19530
rect -7450 18330 -7420 18570
rect -7180 18330 -7050 18570
rect -6810 18330 -6780 18570
rect -7450 18300 -6780 18330
rect -5990 17670 -5330 21750
rect -3001 19400 -2699 19401
rect -3001 19100 -3000 19400
rect -2700 19100 -2699 19400
rect -3001 19099 -2699 19100
rect -1401 19400 -1099 19401
rect -1401 19100 -1400 19400
rect -1100 19100 -1099 19400
rect -1401 19099 -1099 19100
rect 1099 19400 1401 19401
rect 1099 19100 1100 19400
rect 1400 19100 1401 19400
rect 1099 19099 1401 19100
rect 2599 19400 2901 19401
rect 2599 19100 2600 19400
rect 2900 19100 2901 19400
rect 2599 19099 2901 19100
rect -5990 17430 -5960 17670
rect -5720 17430 -5600 17670
rect -5360 17430 -5330 17670
rect 5260 17670 5920 23440
rect 6710 19770 7380 27430
rect 6710 19530 6740 19770
rect 6980 19530 7110 19770
rect 7350 19530 7380 19770
rect 6710 18570 7380 19530
rect 6710 18330 6740 18570
rect 6980 18330 7110 18570
rect 7350 18330 7380 18570
rect 6710 18300 7380 18330
rect -5990 16370 -5330 17430
rect -3101 17500 -2799 17501
rect -3101 17200 -3100 17500
rect -2800 17200 -2799 17500
rect -3101 17199 -2799 17200
rect -2201 17500 -1899 17501
rect -2201 17200 -2200 17500
rect -1900 17200 -1899 17500
rect -2201 17199 -1899 17200
rect -1301 17500 -999 17501
rect -1301 17200 -1300 17500
rect -1000 17200 -999 17500
rect -1301 17199 -999 17200
rect 999 17500 1301 17501
rect 999 17200 1000 17500
rect 1300 17200 1301 17500
rect 999 17199 1301 17200
rect 1899 17500 2201 17501
rect 1899 17200 1900 17500
rect 2200 17200 2201 17500
rect 1899 17199 2201 17200
rect 2799 17500 3101 17501
rect 2799 17200 2800 17500
rect 3100 17200 3101 17500
rect 2799 17199 3101 17200
rect 5260 17430 5290 17670
rect 5530 17430 5650 17670
rect 5890 17430 5920 17670
rect -5990 16130 -5960 16370
rect -5720 16130 -5600 16370
rect -5360 16130 -5330 16370
rect -5990 16100 -5330 16130
rect 5260 16370 5920 17430
rect 5260 16130 5290 16370
rect 5530 16130 5650 16370
rect 5890 16130 5920 16370
rect 5260 16100 5920 16130
<< via4 >>
rect -7420 28000 -7180 28240
rect -7050 28000 -6810 28240
rect -7420 27430 -7180 27670
rect -7050 27430 -6810 27670
rect 6740 28100 6980 28340
rect 7110 28100 7350 28340
rect 6740 27430 6980 27670
rect 7110 27430 7350 27670
rect -7420 19530 -7180 19770
rect -7050 19530 -6810 19770
rect -7420 18330 -7180 18570
rect -7050 18330 -6810 18570
rect -3000 19100 -2700 19400
rect -1400 19100 -1100 19400
rect 1100 19100 1400 19400
rect 2600 19100 2900 19400
rect -5960 17430 -5720 17670
rect -5600 17430 -5360 17670
rect 6740 19530 6980 19770
rect 7110 19530 7350 19770
rect 6740 18330 6980 18570
rect 7110 18330 7350 18570
rect -3100 17200 -2800 17500
rect -2200 17200 -1900 17500
rect -1300 17200 -1000 17500
rect 1000 17200 1300 17500
rect 1900 17200 2200 17500
rect 2800 17200 3100 17500
rect 5290 17430 5530 17670
rect 5650 17430 5890 17670
rect -5960 16130 -5720 16370
rect -5600 16130 -5360 16370
rect 5290 16130 5530 16370
rect 5650 16130 5890 16370
<< metal5 >>
rect -8300 28340 8900 31500
rect -8300 28240 6740 28340
rect -8300 28000 -7420 28240
rect -7180 28000 -7050 28240
rect -6810 28100 6740 28240
rect 6980 28100 7110 28340
rect 7350 28100 8900 28340
rect -6810 28000 8900 28100
rect -8300 27670 8900 28000
rect -8300 27430 -7420 27670
rect -7180 27430 -7050 27670
rect -6810 27430 6740 27670
rect 6980 27430 7110 27670
rect 7350 27430 8900 27670
rect -8300 27400 8900 27430
rect -7700 20660 7380 22520
rect -7700 19770 7380 19800
rect -7700 19530 -7420 19770
rect -7180 19530 -7050 19770
rect -6810 19530 6740 19770
rect 6980 19530 7110 19770
rect 7350 19530 7380 19770
rect -7700 19400 7380 19530
rect -7700 19100 -3000 19400
rect -2700 19100 -1400 19400
rect -1100 19100 1100 19400
rect 1400 19100 2600 19400
rect 2900 19100 7380 19400
rect -7700 18570 7380 19100
rect -7700 18330 -7420 18570
rect -7180 18330 -7050 18570
rect -6810 18330 6740 18570
rect 6980 18330 7110 18570
rect 7350 18330 7380 18570
rect -7700 18300 7380 18330
rect -7700 17670 7380 17700
rect -7700 17430 -5960 17670
rect -5720 17430 -5600 17670
rect -5360 17500 5290 17670
rect -5360 17430 -3100 17500
rect -7700 17200 -3100 17430
rect -2800 17200 -2200 17500
rect -1900 17200 -1300 17500
rect -1000 17200 1000 17500
rect 1300 17200 1900 17500
rect 2200 17200 2800 17500
rect 3100 17430 5290 17500
rect 5530 17430 5650 17670
rect 5890 17430 7380 17670
rect 3100 17200 7380 17430
rect -7700 16370 7380 17200
rect -7700 16130 -5960 16370
rect -5720 16130 -5600 16370
rect -5360 16130 5290 16370
rect 5530 16130 5650 16370
rect 5890 16130 7380 16370
rect -7700 16100 7380 16130
use OTA_fingers_031123_NON_FLAT  OTA_fingers_031123_NON_FLAT_0
timestamp 1679690840
transform 1 0 -1920 0 1 20510
box -5940 -310 9780 16550
use constant_gm_local_030423  constant_gm_local_030423_0
timestamp 1679690840
transform 1 0 0 0 1 16460
box -3840 -15020 3830 3300
<< labels >>
rlabel metal1 3866 30438 4092 30598 1 Vmid
port 1 n
rlabel metal4 3732 32548 3876 32728 1 Vout
port 2 n
rlabel metal1 700 25690 760 25750 1 Vp
port 3 n
rlabel metal1 700 24170 760 24220 1 Vn
port 4 n
rlabel metal2 920 20220 1070 20330 1 Vmirror
port 5 n
rlabel metal5 -4810 16660 -4030 17140 1 Vss
port 6 n
rlabel metal5 -4870 18860 -4090 19340 1 Vdd
port 7 n
<< end >>
