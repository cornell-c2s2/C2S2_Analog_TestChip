magic
tech sky130A
magscale 1 2
timestamp 1683391037
<< nwell >>
rect -4170 1941 4040 3182
rect -3810 1940 3808 1941
<< pwell >>
rect -1040 1150 1034 1742
rect -820 625 818 1117
rect -3755 0 3755 592
rect -3290 -6320 3290 -1008
rect -3290 -13822 3280 -6320
<< nmos >>
rect -830 1346 -580 1546
rect -362 1346 -112 1546
rect 106 1346 356 1546
rect 574 1346 824 1546
rect -610 821 -110 921
rect 108 821 608 921
rect -3545 196 -2545 396
rect -2327 196 -1327 396
rect -1109 196 -109 396
rect 109 196 1109 396
rect 1327 196 2327 396
rect 2545 196 3545 396
<< pmos >>
rect -3591 2726 -2591 2926
rect -2355 2726 -1355 2926
rect -1119 2726 -119 2926
rect 117 2726 1117 2926
rect 1353 2726 2353 2926
rect 2589 2726 3589 2926
rect -3591 2136 -2591 2336
rect -2355 2136 -1355 2336
rect -1119 2136 -119 2336
rect 117 2136 1117 2336
rect 1353 2136 2353 2336
rect 2589 2136 3589 2336
<< ndiff >>
rect -830 1592 -580 1604
rect -830 1558 -818 1592
rect -592 1558 -580 1592
rect -830 1546 -580 1558
rect -362 1592 -112 1604
rect -362 1558 -350 1592
rect -124 1558 -112 1592
rect -362 1546 -112 1558
rect 106 1592 356 1604
rect 106 1558 118 1592
rect 344 1558 356 1592
rect 106 1546 356 1558
rect 574 1592 824 1604
rect 574 1558 586 1592
rect 812 1558 824 1592
rect 574 1546 824 1558
rect -830 1334 -580 1346
rect -830 1300 -818 1334
rect -592 1300 -580 1334
rect -830 1288 -580 1300
rect -362 1334 -112 1346
rect -362 1300 -350 1334
rect -124 1300 -112 1334
rect -362 1288 -112 1300
rect 106 1334 356 1346
rect 106 1300 118 1334
rect 344 1300 356 1334
rect 106 1288 356 1300
rect 574 1334 824 1346
rect 574 1300 586 1334
rect 812 1300 824 1334
rect 574 1288 824 1300
rect -610 967 -110 979
rect -610 933 -598 967
rect -122 933 -110 967
rect -610 921 -110 933
rect 108 967 608 979
rect 108 933 120 967
rect 596 933 608 967
rect 108 921 608 933
rect -610 809 -110 821
rect -610 775 -598 809
rect -122 775 -110 809
rect -610 763 -110 775
rect 108 809 608 821
rect 108 775 120 809
rect 596 775 608 809
rect 108 763 608 775
rect -3545 442 -2545 454
rect -3545 408 -3533 442
rect -2557 408 -2545 442
rect -3545 396 -2545 408
rect -2327 442 -1327 454
rect -2327 408 -2315 442
rect -1339 408 -1327 442
rect -2327 396 -1327 408
rect -1109 442 -109 454
rect -1109 408 -1097 442
rect -121 408 -109 442
rect -1109 396 -109 408
rect 109 442 1109 454
rect 109 408 121 442
rect 1097 408 1109 442
rect 109 396 1109 408
rect 1327 442 2327 454
rect 1327 408 1339 442
rect 2315 408 2327 442
rect 1327 396 2327 408
rect 2545 442 3545 454
rect 2545 408 2557 442
rect 3533 408 3545 442
rect 2545 396 3545 408
rect -3545 184 -2545 196
rect -3545 150 -3533 184
rect -2557 150 -2545 184
rect -3545 138 -2545 150
rect -2327 184 -1327 196
rect -2327 150 -2315 184
rect -1339 150 -1327 184
rect -2327 138 -1327 150
rect -1109 184 -109 196
rect -1109 150 -1097 184
rect -121 150 -109 184
rect -1109 138 -109 150
rect 109 184 1109 196
rect 109 150 121 184
rect 1097 150 1109 184
rect 109 138 1109 150
rect 1327 184 2327 196
rect 1327 150 1339 184
rect 2315 150 2327 184
rect 1327 138 2327 150
rect 2545 184 3545 196
rect 2545 150 2557 184
rect 3533 150 3545 184
rect 2545 138 3545 150
<< pdiff >>
rect -3591 2972 -2591 2984
rect -3591 2938 -3579 2972
rect -2603 2938 -2591 2972
rect -3591 2926 -2591 2938
rect -2355 2972 -1355 2984
rect -2355 2938 -2343 2972
rect -1367 2938 -1355 2972
rect -2355 2926 -1355 2938
rect -1119 2972 -119 2984
rect -1119 2938 -1107 2972
rect -131 2938 -119 2972
rect -1119 2926 -119 2938
rect 117 2972 1117 2984
rect 117 2938 129 2972
rect 1105 2938 1117 2972
rect 117 2926 1117 2938
rect 1353 2972 2353 2984
rect 1353 2938 1365 2972
rect 2341 2938 2353 2972
rect 1353 2926 2353 2938
rect 2589 2972 3589 2984
rect 2589 2938 2601 2972
rect 3577 2938 3589 2972
rect 2589 2926 3589 2938
rect -3591 2714 -2591 2726
rect -3591 2680 -3579 2714
rect -2603 2680 -2591 2714
rect -3591 2668 -2591 2680
rect -2355 2714 -1355 2726
rect -2355 2680 -2343 2714
rect -1367 2680 -1355 2714
rect -2355 2668 -1355 2680
rect -1119 2714 -119 2726
rect -1119 2680 -1107 2714
rect -131 2680 -119 2714
rect -1119 2668 -119 2680
rect 117 2714 1117 2726
rect 117 2680 129 2714
rect 1105 2680 1117 2714
rect 117 2668 1117 2680
rect 1353 2714 2353 2726
rect 1353 2680 1365 2714
rect 2341 2680 2353 2714
rect 1353 2668 2353 2680
rect 2589 2714 3589 2726
rect 2589 2680 2601 2714
rect 3577 2680 3589 2714
rect 2589 2668 3589 2680
rect -3591 2382 -2591 2394
rect -3591 2348 -3579 2382
rect -2603 2348 -2591 2382
rect -3591 2336 -2591 2348
rect -2355 2382 -1355 2394
rect -2355 2348 -2343 2382
rect -1367 2348 -1355 2382
rect -2355 2336 -1355 2348
rect -1119 2382 -119 2394
rect -1119 2348 -1107 2382
rect -131 2348 -119 2382
rect -1119 2336 -119 2348
rect 117 2382 1117 2394
rect 117 2348 129 2382
rect 1105 2348 1117 2382
rect 117 2336 1117 2348
rect 1353 2382 2353 2394
rect 1353 2348 1365 2382
rect 2341 2348 2353 2382
rect 1353 2336 2353 2348
rect 2589 2382 3589 2394
rect 2589 2348 2601 2382
rect 3577 2348 3589 2382
rect 2589 2336 3589 2348
rect -3591 2124 -2591 2136
rect -3591 2090 -3579 2124
rect -2603 2090 -2591 2124
rect -3591 2078 -2591 2090
rect -2355 2124 -1355 2136
rect -2355 2090 -2343 2124
rect -1367 2090 -1355 2124
rect -2355 2078 -1355 2090
rect -1119 2124 -119 2136
rect -1119 2090 -1107 2124
rect -131 2090 -119 2124
rect -1119 2078 -119 2090
rect 117 2124 1117 2136
rect 117 2090 129 2124
rect 1105 2090 1117 2124
rect 117 2078 1117 2090
rect 1353 2124 2353 2136
rect 1353 2090 1365 2124
rect 2341 2090 2353 2124
rect 1353 2078 2353 2090
rect 2589 2124 3589 2136
rect 2589 2090 2601 2124
rect 3577 2090 3589 2124
rect 2589 2078 3589 2090
<< ndiffc >>
rect -818 1558 -592 1592
rect -350 1558 -124 1592
rect 118 1558 344 1592
rect 586 1558 812 1592
rect -818 1300 -592 1334
rect -350 1300 -124 1334
rect 118 1300 344 1334
rect 586 1300 812 1334
rect -598 933 -122 967
rect 120 933 596 967
rect -598 775 -122 809
rect 120 775 596 809
rect -3533 408 -2557 442
rect -2315 408 -1339 442
rect -1097 408 -121 442
rect 121 408 1097 442
rect 1339 408 2315 442
rect 2557 408 3533 442
rect -3533 150 -2557 184
rect -2315 150 -1339 184
rect -1097 150 -121 184
rect 121 150 1097 184
rect 1339 150 2315 184
rect 2557 150 3533 184
<< pdiffc >>
rect -3579 2938 -2603 2972
rect -2343 2938 -1367 2972
rect -1107 2938 -131 2972
rect 129 2938 1105 2972
rect 1365 2938 2341 2972
rect 2601 2938 3577 2972
rect -3579 2680 -2603 2714
rect -2343 2680 -1367 2714
rect -1107 2680 -131 2714
rect 129 2680 1105 2714
rect 1365 2680 2341 2714
rect 2601 2680 3577 2714
rect -3579 2348 -2603 2382
rect -2343 2348 -1367 2382
rect -1107 2348 -131 2382
rect 129 2348 1105 2382
rect 1365 2348 2341 2382
rect 2601 2348 3577 2382
rect -3579 2090 -2603 2124
rect -2343 2090 -1367 2124
rect -1107 2090 -131 2124
rect 129 2090 1105 2124
rect 1365 2090 2341 2124
rect 2601 2090 3577 2124
<< psubdiff >>
rect -1004 1672 -908 1706
rect 902 1672 998 1706
rect -1004 1610 -970 1672
rect 964 1610 998 1672
rect -1004 1220 -970 1282
rect 964 1220 998 1282
rect -1004 1186 -908 1220
rect 902 1186 998 1220
rect -784 1047 -688 1081
rect 686 1047 782 1081
rect -784 985 -750 1047
rect 748 985 782 1047
rect -784 695 -750 757
rect 748 695 782 757
rect -784 661 -688 695
rect 686 661 782 695
rect -3719 522 -3623 556
rect 3623 522 3719 556
rect -3719 460 -3685 522
rect 3685 460 3719 522
rect -3719 70 -3685 132
rect 3685 70 3719 132
rect -3719 36 -3623 70
rect 3623 36 3719 70
rect -3240 -1240 -3120 -1216
rect -3240 -1384 -3120 -1360
rect -3240 -4240 -3120 -4216
rect -3240 -4384 -3120 -4360
rect -3240 -7240 -3120 -7216
rect -3240 -7384 -3120 -7360
rect -3240 -10240 -3120 -10216
rect -3240 -10384 -3120 -10360
rect -3240 -13240 -3120 -13216
rect -3240 -13384 -3120 -13360
rect 3130 -1240 3250 -1216
rect 3130 -1384 3250 -1360
rect 3130 -4240 3250 -4216
rect 3130 -4384 3250 -4360
rect 3130 -7240 3250 -7216
rect 3130 -7384 3250 -7360
rect 3130 -10240 3250 -10216
rect 3130 -10384 3250 -10360
rect 3130 -13240 3250 -13216
rect 3130 -13384 3250 -13360
<< nsubdiff >>
rect -3774 3052 -3678 3086
rect 3676 3052 3772 3086
rect -3774 2990 -3740 3052
rect 3738 2990 3772 3052
rect -3774 2600 -3740 2662
rect 3738 2600 3772 2662
rect -3774 2566 -3678 2600
rect 3676 2566 3772 2600
rect -3774 2462 -3678 2496
rect 3676 2462 3772 2496
rect -3774 2400 -3740 2462
rect 3738 2400 3772 2462
rect -3774 2010 -3740 2072
rect 3738 2010 3772 2072
rect -3774 1976 -3678 2010
rect 3676 1976 3772 2010
<< psubdiffcont >>
rect -908 1672 902 1706
rect -1004 1282 -970 1610
rect 964 1282 998 1610
rect -908 1186 902 1220
rect -688 1047 686 1081
rect -784 757 -750 985
rect 748 757 782 985
rect -688 661 686 695
rect -3623 522 3623 556
rect -3719 132 -3685 460
rect 3685 132 3719 460
rect -3623 36 3623 70
rect -3240 -1360 -3120 -1240
rect -3240 -4360 -3120 -4240
rect -3240 -7360 -3120 -7240
rect -3240 -10360 -3120 -10240
rect -3240 -13360 -3120 -13240
rect 3130 -1360 3250 -1240
rect 3130 -4360 3250 -4240
rect 3130 -7360 3250 -7240
rect 3130 -10360 3250 -10240
rect 3130 -13360 3250 -13240
<< nsubdiffcont >>
rect -3678 3052 3676 3086
rect -3774 2662 -3740 2990
rect 3738 2662 3772 2990
rect -3678 2566 3676 2600
rect -3678 2462 3676 2496
rect -3774 2072 -3740 2400
rect 3738 2072 3772 2400
rect -3678 1976 3676 2010
<< poly >>
rect -3688 2910 -3591 2926
rect -3688 2742 -3672 2910
rect -3638 2742 -3591 2910
rect -3688 2726 -3591 2742
rect -2591 2910 -2494 2926
rect -2591 2742 -2544 2910
rect -2510 2742 -2494 2910
rect -2591 2726 -2494 2742
rect -2452 2910 -2355 2926
rect -2452 2742 -2436 2910
rect -2402 2742 -2355 2910
rect -2452 2726 -2355 2742
rect -1355 2910 -1258 2926
rect -1355 2742 -1308 2910
rect -1274 2742 -1258 2910
rect -1355 2726 -1258 2742
rect -1216 2910 -1119 2926
rect -1216 2742 -1200 2910
rect -1166 2742 -1119 2910
rect -1216 2726 -1119 2742
rect -119 2910 -22 2926
rect -119 2742 -72 2910
rect -38 2742 -22 2910
rect -119 2726 -22 2742
rect 20 2910 117 2926
rect 20 2742 36 2910
rect 70 2742 117 2910
rect 20 2726 117 2742
rect 1117 2910 1214 2926
rect 1117 2742 1164 2910
rect 1198 2742 1214 2910
rect 1117 2726 1214 2742
rect 1256 2910 1353 2926
rect 1256 2742 1272 2910
rect 1306 2742 1353 2910
rect 1256 2726 1353 2742
rect 2353 2910 2450 2926
rect 2353 2742 2400 2910
rect 2434 2742 2450 2910
rect 2353 2726 2450 2742
rect 2492 2910 2589 2926
rect 2492 2742 2508 2910
rect 2542 2742 2589 2910
rect 2492 2726 2589 2742
rect 3589 2910 3686 2926
rect 3589 2742 3636 2910
rect 3670 2742 3686 2910
rect 3589 2726 3686 2742
rect -3688 2320 -3591 2336
rect -3688 2152 -3672 2320
rect -3638 2152 -3591 2320
rect -3688 2136 -3591 2152
rect -2591 2320 -2494 2336
rect -2591 2152 -2544 2320
rect -2510 2152 -2494 2320
rect -2591 2136 -2494 2152
rect -2452 2320 -2355 2336
rect -2452 2152 -2436 2320
rect -2402 2152 -2355 2320
rect -2452 2136 -2355 2152
rect -1355 2320 -1258 2336
rect -1355 2152 -1308 2320
rect -1274 2152 -1258 2320
rect -1355 2136 -1258 2152
rect -1216 2320 -1119 2336
rect -1216 2152 -1200 2320
rect -1166 2152 -1119 2320
rect -1216 2136 -1119 2152
rect -119 2320 -22 2336
rect -119 2152 -72 2320
rect -38 2152 -22 2320
rect -119 2136 -22 2152
rect 20 2320 117 2336
rect 20 2152 36 2320
rect 70 2152 117 2320
rect 20 2136 117 2152
rect 1117 2320 1214 2336
rect 1117 2152 1164 2320
rect 1198 2152 1214 2320
rect 1117 2136 1214 2152
rect 1256 2320 1353 2336
rect 1256 2152 1272 2320
rect 1306 2152 1353 2320
rect 1256 2136 1353 2152
rect 2353 2320 2450 2336
rect 2353 2152 2400 2320
rect 2434 2152 2450 2320
rect 2353 2136 2450 2152
rect 2492 2320 2589 2336
rect 2492 2152 2508 2320
rect 2542 2152 2589 2320
rect 2492 2136 2589 2152
rect 3589 2320 3686 2336
rect 3589 2152 3636 2320
rect 3670 2152 3686 2320
rect 3589 2136 3686 2152
rect -918 1530 -830 1546
rect -918 1362 -902 1530
rect -868 1362 -830 1530
rect -918 1346 -830 1362
rect -580 1530 -492 1546
rect -580 1362 -542 1530
rect -508 1362 -492 1530
rect -580 1346 -492 1362
rect -450 1530 -362 1546
rect -450 1362 -434 1530
rect -400 1362 -362 1530
rect -450 1346 -362 1362
rect -112 1530 -24 1546
rect -112 1362 -74 1530
rect -40 1362 -24 1530
rect -112 1346 -24 1362
rect 18 1530 106 1546
rect 18 1362 34 1530
rect 68 1362 106 1530
rect 18 1346 106 1362
rect 356 1530 444 1546
rect 356 1362 394 1530
rect 428 1362 444 1530
rect 356 1346 444 1362
rect 486 1530 574 1546
rect 486 1362 502 1530
rect 536 1362 574 1530
rect 486 1346 574 1362
rect 824 1530 912 1546
rect 824 1362 862 1530
rect 896 1362 912 1530
rect 824 1346 912 1362
rect -698 905 -610 921
rect -698 837 -682 905
rect -648 837 -610 905
rect -698 821 -610 837
rect -110 905 -22 921
rect -110 837 -72 905
rect -38 837 -22 905
rect -110 821 -22 837
rect 20 905 108 921
rect 20 837 36 905
rect 70 837 108 905
rect 20 821 108 837
rect 608 905 696 921
rect 608 837 646 905
rect 680 837 696 905
rect 608 821 696 837
rect -3633 380 -3545 396
rect -3633 212 -3617 380
rect -3583 212 -3545 380
rect -3633 196 -3545 212
rect -2545 380 -2457 396
rect -2545 212 -2507 380
rect -2473 212 -2457 380
rect -2545 196 -2457 212
rect -2415 380 -2327 396
rect -2415 212 -2399 380
rect -2365 212 -2327 380
rect -2415 196 -2327 212
rect -1327 380 -1239 396
rect -1327 212 -1289 380
rect -1255 212 -1239 380
rect -1327 196 -1239 212
rect -1197 380 -1109 396
rect -1197 212 -1181 380
rect -1147 212 -1109 380
rect -1197 196 -1109 212
rect -109 380 -21 396
rect -109 212 -71 380
rect -37 212 -21 380
rect -109 196 -21 212
rect 21 380 109 396
rect 21 212 37 380
rect 71 212 109 380
rect 21 196 109 212
rect 1109 380 1197 396
rect 1109 212 1147 380
rect 1181 212 1197 380
rect 1109 196 1197 212
rect 1239 380 1327 396
rect 1239 212 1255 380
rect 1289 212 1327 380
rect 1239 196 1327 212
rect 2327 380 2415 396
rect 2327 212 2365 380
rect 2399 212 2415 380
rect 2327 196 2415 212
rect 2457 380 2545 396
rect 2457 212 2473 380
rect 2507 212 2545 380
rect 2457 196 2545 212
rect 3545 380 3633 396
rect 3545 212 3583 380
rect 3617 212 3633 380
rect 3545 196 3633 212
<< polycont >>
rect -3672 2742 -3638 2910
rect -2544 2742 -2510 2910
rect -2436 2742 -2402 2910
rect -1308 2742 -1274 2910
rect -1200 2742 -1166 2910
rect -72 2742 -38 2910
rect 36 2742 70 2910
rect 1164 2742 1198 2910
rect 1272 2742 1306 2910
rect 2400 2742 2434 2910
rect 2508 2742 2542 2910
rect 3636 2742 3670 2910
rect -3672 2152 -3638 2320
rect -2544 2152 -2510 2320
rect -2436 2152 -2402 2320
rect -1308 2152 -1274 2320
rect -1200 2152 -1166 2320
rect -72 2152 -38 2320
rect 36 2152 70 2320
rect 1164 2152 1198 2320
rect 1272 2152 1306 2320
rect 2400 2152 2434 2320
rect 2508 2152 2542 2320
rect 3636 2152 3670 2320
rect -902 1362 -868 1530
rect -542 1362 -508 1530
rect -434 1362 -400 1530
rect -74 1362 -40 1530
rect 34 1362 68 1530
rect 394 1362 428 1530
rect 502 1362 536 1530
rect 862 1362 896 1530
rect -682 837 -648 905
rect -72 837 -38 905
rect 36 837 70 905
rect 646 837 680 905
rect -3617 212 -3583 380
rect -2507 212 -2473 380
rect -2399 212 -2365 380
rect -1289 212 -1255 380
rect -1181 212 -1147 380
rect -71 212 -37 380
rect 37 212 71 380
rect 1147 212 1181 380
rect 1255 212 1289 380
rect 2365 212 2399 380
rect 2473 212 2507 380
rect 3583 212 3617 380
<< xpolycontact >>
rect -2843 -728 -1697 -296
rect -2843 -14960 -1697 -14528
rect -1323 -728 -177 -296
rect -1323 -14960 -177 -14528
rect 187 -722 1333 -290
rect 187 -14954 1333 -14522
rect 1697 -722 2843 -290
rect 1697 -14954 2843 -14522
<< xpolyres >>
rect -2843 -14528 -1697 -728
rect -1323 -14528 -177 -728
rect 187 -14522 1333 -722
rect 1697 -14522 2843 -722
<< locali >>
rect -3774 3052 -3678 3086
rect 3676 3052 3772 3086
rect -3774 2990 -3740 3052
rect 3738 2990 3772 3052
rect -3595 2938 -3579 2972
rect -2603 2938 -2587 2972
rect -2359 2938 -2343 2972
rect -1367 2938 -1351 2972
rect -1123 2938 -1107 2972
rect -131 2938 -115 2972
rect 113 2938 129 2972
rect 1105 2938 1121 2972
rect 1349 2938 1365 2972
rect 2341 2938 2357 2972
rect 2585 2938 2601 2972
rect 3577 2938 3593 2972
rect -3672 2910 -3638 2926
rect -3672 2726 -3638 2742
rect -2544 2910 -2510 2926
rect -2544 2726 -2510 2742
rect -2436 2910 -2402 2926
rect -2436 2726 -2402 2742
rect -1308 2910 -1274 2926
rect -1308 2726 -1274 2742
rect -1200 2910 -1166 2926
rect -1200 2726 -1166 2742
rect -72 2910 -38 2926
rect -72 2726 -38 2742
rect 36 2910 70 2926
rect 36 2726 70 2742
rect 1164 2910 1198 2926
rect 1164 2726 1198 2742
rect 1272 2910 1306 2926
rect 1272 2726 1306 2742
rect 2400 2910 2434 2926
rect 2400 2726 2434 2742
rect 2508 2910 2542 2926
rect 2508 2726 2542 2742
rect 3636 2910 3670 2926
rect 3636 2726 3670 2742
rect -3595 2680 -3579 2714
rect -2603 2680 -2587 2714
rect -2359 2680 -2343 2714
rect -1367 2680 -1351 2714
rect -1123 2680 -1107 2714
rect -131 2680 -115 2714
rect 113 2680 129 2714
rect 1105 2680 1121 2714
rect 1349 2680 1365 2714
rect 2341 2680 2357 2714
rect 2585 2680 2601 2714
rect 3577 2680 3593 2714
rect -3774 2600 -3740 2662
rect 3738 2600 3772 2662
rect -3774 2566 -3678 2600
rect 3676 2566 3772 2600
rect -3774 2462 -3678 2496
rect 3676 2462 3772 2496
rect -3774 2400 -3740 2462
rect 3738 2400 3772 2462
rect -3595 2348 -3579 2382
rect -2603 2348 -2587 2382
rect -2359 2348 -2343 2382
rect -1367 2348 -1351 2382
rect -1123 2348 -1107 2382
rect -131 2348 -115 2382
rect 113 2348 129 2382
rect 1105 2348 1121 2382
rect 1349 2348 1365 2382
rect 2341 2348 2357 2382
rect 2585 2348 2601 2382
rect 3577 2348 3593 2382
rect -3672 2320 -3638 2336
rect -3672 2136 -3638 2152
rect -2544 2320 -2510 2336
rect -2544 2136 -2510 2152
rect -2436 2320 -2402 2336
rect -2436 2136 -2402 2152
rect -1308 2320 -1274 2336
rect -1308 2136 -1274 2152
rect -1200 2320 -1166 2336
rect -1200 2136 -1166 2152
rect -72 2320 -38 2336
rect -72 2136 -38 2152
rect 36 2320 70 2336
rect 36 2136 70 2152
rect 1164 2320 1198 2336
rect 1164 2136 1198 2152
rect 1272 2320 1306 2336
rect 1272 2136 1306 2152
rect 2400 2320 2434 2336
rect 2400 2136 2434 2152
rect 2508 2320 2542 2336
rect 2508 2136 2542 2152
rect 3636 2320 3670 2336
rect 3636 2136 3670 2152
rect -3595 2090 -3579 2124
rect -2603 2090 -2587 2124
rect -2359 2090 -2343 2124
rect -1367 2090 -1351 2124
rect -1123 2090 -1107 2124
rect -131 2090 -115 2124
rect 113 2090 129 2124
rect 1105 2090 1121 2124
rect 1349 2090 1365 2124
rect 2341 2090 2357 2124
rect 2585 2090 2601 2124
rect 3577 2090 3593 2124
rect -3774 2010 -3740 2072
rect 3738 2010 3772 2072
rect -3774 1976 -3678 2010
rect 3676 1976 3772 2010
rect -1004 1672 -908 1706
rect 902 1672 998 1706
rect -1004 1610 -970 1672
rect 964 1610 998 1672
rect -834 1558 -818 1592
rect -592 1558 -576 1592
rect -366 1558 -350 1592
rect -124 1558 -108 1592
rect 102 1558 118 1592
rect 344 1558 360 1592
rect 570 1558 586 1592
rect 812 1558 828 1592
rect -902 1530 -868 1546
rect -902 1346 -868 1362
rect -542 1530 -508 1546
rect -542 1346 -508 1362
rect -434 1530 -400 1546
rect -434 1346 -400 1362
rect -74 1530 -40 1546
rect -74 1346 -40 1362
rect 34 1530 68 1546
rect 34 1346 68 1362
rect 394 1530 428 1546
rect 394 1346 428 1362
rect 502 1530 536 1546
rect 502 1346 536 1362
rect 862 1530 896 1546
rect 862 1346 896 1362
rect -834 1300 -818 1334
rect -592 1300 -576 1334
rect -366 1300 -350 1334
rect -124 1300 -108 1334
rect 102 1300 118 1334
rect 344 1300 360 1334
rect 570 1300 586 1334
rect 812 1300 828 1334
rect -1004 1220 -970 1282
rect 964 1220 998 1282
rect -1004 1186 -908 1220
rect 902 1186 998 1220
rect -784 1047 -688 1070
rect 686 1047 782 1070
rect -784 985 -750 1047
rect 748 985 782 1047
rect -614 933 -598 967
rect -122 933 -106 967
rect 104 933 120 967
rect 596 933 612 967
rect -682 905 -648 921
rect -682 821 -648 837
rect -72 905 -38 921
rect -72 821 -38 837
rect 36 905 70 921
rect 36 821 70 837
rect 646 905 680 921
rect 646 821 680 837
rect -614 775 -598 809
rect -122 775 -106 809
rect 104 775 120 809
rect 596 775 612 809
rect -784 695 -750 757
rect 748 695 782 757
rect -784 661 -688 695
rect 686 661 782 695
rect -3719 522 -3623 556
rect 3623 522 3719 556
rect -3719 460 -3685 522
rect 3685 460 3719 522
rect -3549 408 -3533 442
rect -2557 408 -2541 442
rect -2331 408 -2315 442
rect -1339 408 -1323 442
rect -1113 408 -1097 442
rect -121 408 -105 442
rect 105 408 121 442
rect 1097 408 1113 442
rect 1323 408 1339 442
rect 2315 408 2331 442
rect 2541 408 2557 442
rect 3533 408 3549 442
rect -3617 380 -3583 396
rect -3617 196 -3583 212
rect -2507 380 -2473 396
rect -2507 196 -2473 212
rect -2399 380 -2365 396
rect -2399 196 -2365 212
rect -1289 380 -1255 396
rect -1289 196 -1255 212
rect -1181 380 -1147 396
rect -1181 196 -1147 212
rect -71 380 -37 396
rect -71 196 -37 212
rect 37 380 71 396
rect 37 196 71 212
rect 1147 380 1181 396
rect 1147 196 1181 212
rect 1255 380 1289 396
rect 1255 196 1289 212
rect 2365 380 2399 396
rect 2365 196 2399 212
rect 2473 380 2507 396
rect 2473 196 2507 212
rect 3583 380 3617 396
rect 3583 196 3617 212
rect -3549 150 -3533 184
rect -2557 150 -2541 184
rect -2331 150 -2315 184
rect -1339 150 -1323 184
rect -1113 150 -1097 184
rect -121 150 -105 184
rect 105 150 121 184
rect 1097 150 1113 184
rect 1323 150 1339 184
rect 2315 150 2331 184
rect 2541 150 2557 184
rect 3533 150 3549 184
rect -3719 70 -3685 132
rect 3685 70 3719 132
rect -3719 36 -3623 70
rect 3623 36 3719 70
rect -3240 -1240 -3120 -1224
rect -3240 -1376 -3120 -1360
rect 3130 -1240 3250 -1224
rect 3130 -1376 3250 -1360
rect -3240 -4240 -3120 -4224
rect -3240 -4376 -3120 -4360
rect 3130 -4240 3250 -4224
rect 3130 -4376 3250 -4360
rect -3240 -7240 -3120 -7224
rect -3240 -7376 -3120 -7360
rect 3130 -7240 3250 -7224
rect 3130 -7376 3250 -7360
rect -3240 -10240 -3120 -10224
rect -3240 -10376 -3120 -10360
rect 3130 -10240 3250 -10224
rect 3130 -10376 3250 -10360
rect -3240 -13240 -3120 -13224
rect -3240 -13376 -3120 -13360
rect 3130 -13240 3250 -13224
rect 3130 -13376 3250 -13360
<< viali >>
rect -3220 3086 -3060 3180
rect -2160 3086 -2000 3180
rect -700 3086 -540 3180
rect 520 3086 680 3180
rect 2000 3086 2160 3180
rect 3000 3086 3160 3180
rect -3220 3052 -3060 3086
rect -2160 3052 -2000 3086
rect -700 3052 -540 3086
rect 520 3052 680 3086
rect 2000 3052 2160 3086
rect 3000 3052 3160 3086
rect -3220 3020 -3060 3052
rect -2160 3020 -2000 3052
rect -700 3020 -540 3052
rect 520 3020 680 3052
rect 2000 3020 2160 3052
rect 3000 3020 3160 3052
rect -3579 2938 -2603 2972
rect -2343 2938 -1367 2972
rect -1107 2938 -131 2972
rect 129 2938 1105 2972
rect 1365 2938 2341 2972
rect 2601 2938 3577 2972
rect -3672 2742 -3638 2910
rect -2544 2742 -2510 2910
rect -2436 2742 -2402 2910
rect -1308 2742 -1274 2910
rect -1200 2742 -1166 2910
rect -72 2742 -38 2910
rect 36 2742 70 2910
rect 1164 2742 1198 2910
rect 1272 2742 1306 2910
rect 2400 2742 2434 2910
rect 2508 2742 2542 2910
rect 3636 2742 3670 2910
rect -3579 2680 -2603 2714
rect -2343 2680 -1367 2714
rect -1107 2680 -131 2714
rect 129 2680 1105 2714
rect 1365 2680 2341 2714
rect 2601 2680 3577 2714
rect -3220 2566 -3060 2600
rect -2160 2566 -2000 2600
rect -700 2566 -540 2600
rect 520 2566 680 2600
rect 2000 2566 2160 2600
rect 3000 2566 3160 2600
rect -3220 2496 -3060 2566
rect -2160 2496 -2000 2566
rect -700 2496 -540 2566
rect 520 2496 680 2566
rect 2000 2496 2160 2566
rect 3000 2496 3160 2566
rect -3220 2462 -3060 2496
rect -2160 2462 -2000 2496
rect -700 2462 -540 2496
rect 520 2462 680 2496
rect 2000 2462 2160 2496
rect 3000 2462 3160 2496
rect -3220 2440 -3060 2462
rect -2160 2440 -2000 2462
rect -700 2440 -540 2462
rect 520 2440 680 2462
rect 2000 2440 2160 2462
rect 3000 2440 3160 2462
rect -3579 2348 -2603 2382
rect -2343 2348 -1367 2382
rect -1107 2348 -131 2382
rect 129 2348 1105 2382
rect 1365 2348 2341 2382
rect 2601 2348 3577 2382
rect -3672 2152 -3638 2320
rect -2544 2152 -2510 2320
rect -2436 2152 -2402 2320
rect -1308 2152 -1274 2320
rect -1200 2152 -1166 2320
rect -72 2152 -38 2320
rect 36 2152 70 2320
rect 1164 2152 1198 2320
rect 1272 2152 1306 2320
rect 2400 2152 2434 2320
rect 2508 2152 2542 2320
rect 3636 2152 3670 2320
rect -3579 2090 -2603 2124
rect -2343 2090 -1367 2124
rect -1107 2090 -131 2124
rect 129 2090 1105 2124
rect 1365 2090 2341 2124
rect 2601 2090 3577 2124
rect -818 1558 -592 1592
rect -350 1558 -124 1592
rect 118 1558 344 1592
rect 586 1558 812 1592
rect -902 1362 -868 1530
rect -542 1362 -508 1530
rect -434 1362 -400 1530
rect -74 1362 -40 1530
rect 34 1362 68 1530
rect 394 1362 428 1530
rect 502 1362 536 1530
rect 862 1362 896 1530
rect -818 1300 -592 1334
rect -350 1300 -124 1334
rect 118 1300 344 1334
rect 586 1300 812 1334
rect -840 1186 -620 1220
rect -320 1186 -100 1220
rect 100 1186 320 1220
rect 650 1186 870 1220
rect -840 1081 -620 1186
rect -320 1081 -100 1186
rect 100 1081 320 1186
rect 650 1081 870 1186
rect -840 1070 -688 1081
rect -688 1070 -620 1081
rect -320 1070 -100 1081
rect 100 1070 320 1081
rect 650 1070 686 1081
rect 686 1070 870 1081
rect -598 933 -122 967
rect 120 933 596 967
rect -682 837 -648 905
rect -72 837 -38 905
rect 36 837 70 905
rect 646 837 680 905
rect -598 775 -122 809
rect 120 775 596 809
rect -3200 556 -3020 660
rect -2060 556 -1880 660
rect -1080 556 -900 670
rect -310 661 -130 670
rect 130 661 310 670
rect -310 556 -130 661
rect 130 556 310 661
rect 850 556 1030 660
rect 1920 556 2100 670
rect 2920 556 3100 670
rect -3200 530 -3020 556
rect -2060 530 -1880 556
rect -1080 540 -900 556
rect -310 540 -130 556
rect 130 540 310 556
rect 850 530 1030 556
rect 1920 540 2100 556
rect 2920 540 3100 556
rect -3533 408 -2557 442
rect -2315 408 -1339 442
rect -1097 408 -121 442
rect 121 408 1097 442
rect 1339 408 2315 442
rect 2557 408 3533 442
rect -3617 212 -3583 380
rect -2507 212 -2473 380
rect -2399 212 -2365 380
rect -1289 212 -1255 380
rect -1181 212 -1147 380
rect -71 212 -37 380
rect 37 212 71 380
rect 1147 212 1181 380
rect 1255 212 1289 380
rect 2365 212 2399 380
rect 2473 212 2507 380
rect 3583 212 3617 380
rect -3533 150 -2557 184
rect -2315 150 -1339 184
rect -1097 150 -121 184
rect 121 150 1097 184
rect 1339 150 2315 184
rect 2557 150 3533 184
rect -2827 -711 -1713 -314
rect -1307 -711 -193 -314
rect 203 -705 1317 -308
rect 1713 -705 2827 -308
rect -3240 -1360 -3120 -1240
rect 3130 -1360 3250 -1240
rect -3240 -4360 -3120 -4240
rect 3130 -4360 3250 -4240
rect -3240 -7360 -3120 -7240
rect 3130 -7360 3250 -7240
rect -3240 -10360 -3120 -10240
rect 3130 -10360 3250 -10240
rect -3240 -13360 -3120 -13240
rect 3130 -13360 3250 -13240
rect -2827 -14942 -1713 -14545
rect -1307 -14942 -193 -14545
rect 203 -14936 1317 -14539
rect 1713 -14936 2827 -14539
<< metal1 >>
rect -3232 3180 -3048 3186
rect -2172 3180 -1988 3186
rect -712 3180 -528 3186
rect 508 3180 692 3186
rect 1988 3180 2172 3186
rect 2988 3180 3172 3186
rect -3600 3020 -3220 3180
rect -3060 3020 -2160 3180
rect -2000 3020 -700 3180
rect -540 3020 520 3180
rect 680 3020 2000 3180
rect 2160 3020 3000 3180
rect 3160 3020 3600 3180
rect -3600 2972 3600 3020
rect -3600 2938 -3579 2972
rect -2603 2960 -2343 2972
rect -2603 2938 -2580 2960
rect -3678 2910 -3632 2922
rect -3600 2920 -2580 2938
rect -2360 2938 -2343 2960
rect -1367 2960 -1107 2972
rect -1367 2938 -1355 2960
rect -2360 2932 -1355 2938
rect -1120 2938 -1107 2960
rect -131 2960 129 2972
rect -131 2938 -119 2960
rect -1120 2932 -119 2938
rect 117 2938 129 2960
rect 1105 2960 1365 2972
rect 1105 2938 1120 2960
rect 117 2932 1120 2938
rect -3678 2742 -3672 2910
rect -3638 2870 -3632 2910
rect -2550 2910 -2504 2922
rect -2550 2870 -2544 2910
rect -3638 2742 -2544 2870
rect -2510 2870 -2504 2910
rect -2442 2910 -2396 2922
rect -2360 2920 -1360 2932
rect -2442 2870 -2436 2910
rect -2510 2742 -2436 2870
rect -2402 2870 -2396 2910
rect -1314 2910 -1268 2922
rect -1314 2870 -1308 2910
rect -2402 2860 -1308 2870
rect -2402 2790 -1720 2860
rect -1650 2790 -1500 2860
rect -1430 2790 -1308 2860
rect -2402 2742 -1308 2790
rect -1274 2870 -1268 2910
rect -1206 2910 -1160 2922
rect -1120 2920 -120 2932
rect -1206 2870 -1200 2910
rect -1274 2742 -1200 2870
rect -1166 2870 -1160 2910
rect -78 2910 -32 2922
rect -78 2870 -72 2910
rect -1166 2742 -72 2870
rect -38 2870 -32 2910
rect 30 2910 76 2922
rect 120 2920 1120 2932
rect 1340 2938 1365 2960
rect 2341 2960 2601 2972
rect 2341 2938 2360 2960
rect 30 2870 36 2910
rect -38 2742 36 2870
rect 70 2870 76 2910
rect 1158 2910 1204 2922
rect 1158 2870 1164 2910
rect 70 2742 1164 2870
rect 1198 2870 1204 2910
rect 1266 2910 1312 2922
rect 1340 2920 2360 2938
rect 2580 2938 2601 2960
rect 3577 2938 3600 2972
rect 1266 2870 1272 2910
rect 1198 2742 1272 2870
rect 1306 2870 1312 2910
rect 2394 2910 2440 2922
rect 2394 2870 2400 2910
rect 1306 2860 2400 2870
rect 1306 2790 1460 2860
rect 1530 2790 1700 2860
rect 1770 2790 2400 2860
rect 1306 2742 2400 2790
rect 2434 2870 2440 2910
rect 2502 2910 2548 2922
rect 2580 2920 3600 2938
rect 2502 2870 2508 2910
rect 2434 2742 2508 2870
rect 2542 2870 2548 2910
rect 3630 2910 3676 2922
rect 3630 2870 3636 2910
rect 2542 2742 3636 2870
rect 3670 2742 3676 2910
rect -3678 2730 3676 2742
rect -3678 2714 3670 2730
rect -3678 2680 -3579 2714
rect -2603 2680 -2343 2714
rect -1367 2680 -1107 2714
rect -131 2680 129 2714
rect 1105 2680 1365 2714
rect 2341 2680 2601 2714
rect 3577 2680 3670 2714
rect -3678 2658 3670 2680
rect -3232 2600 -3048 2606
rect -2172 2600 -1988 2606
rect -712 2600 -528 2606
rect 508 2600 692 2606
rect 1988 2600 2172 2606
rect 2988 2600 3172 2606
rect -3600 2440 -3220 2600
rect -3060 2440 -2160 2600
rect -2000 2440 -700 2600
rect -540 2440 520 2600
rect 680 2440 2000 2600
rect 2160 2440 3000 2600
rect 3160 2440 3600 2600
rect -3600 2382 3600 2440
rect -3600 2360 -3579 2382
rect -3591 2348 -3579 2360
rect -2603 2370 -2343 2382
rect -2603 2348 -2591 2370
rect -3591 2342 -2591 2348
rect -2355 2348 -2343 2370
rect -1367 2370 -1107 2382
rect -1367 2348 -1355 2370
rect -2355 2342 -1355 2348
rect -1119 2348 -1107 2370
rect -131 2370 129 2382
rect -131 2348 -119 2370
rect -1119 2342 -119 2348
rect 117 2348 129 2370
rect 1105 2370 1365 2382
rect 1105 2348 1117 2370
rect 117 2342 1117 2348
rect 1353 2348 1365 2370
rect 2341 2370 2601 2382
rect 2341 2348 2353 2370
rect 1353 2342 2353 2348
rect 2589 2348 2601 2370
rect 3577 2360 3600 2382
rect 3577 2348 3589 2360
rect 2589 2342 3589 2348
rect -3678 2320 -3632 2332
rect -3678 2280 -3672 2320
rect -3680 2190 -3672 2280
rect -3678 2152 -3672 2190
rect -3638 2280 -3632 2320
rect -2550 2320 -2504 2332
rect -2550 2280 -2544 2320
rect -3638 2190 -2544 2280
rect -3638 2152 -3632 2190
rect -3678 2140 -3632 2152
rect -2550 2152 -2544 2190
rect -2510 2280 -2504 2320
rect -2442 2320 -2396 2332
rect -2442 2280 -2436 2320
rect -2510 2190 -2436 2280
rect -2510 2152 -2504 2190
rect -2550 2140 -2504 2152
rect -2442 2152 -2436 2190
rect -2402 2280 -2396 2320
rect -1314 2320 -1268 2332
rect -1314 2280 -1308 2320
rect -2402 2270 -1308 2280
rect -2402 2200 -1720 2270
rect -1650 2200 -1500 2270
rect -1430 2200 -1308 2270
rect -2402 2190 -1308 2200
rect -2402 2152 -2396 2190
rect -2442 2140 -2396 2152
rect -1314 2152 -1308 2190
rect -1274 2280 -1268 2320
rect -1206 2320 -1160 2332
rect -1206 2280 -1200 2320
rect -1274 2190 -1200 2280
rect -1274 2152 -1268 2190
rect -1314 2140 -1268 2152
rect -1206 2152 -1200 2190
rect -1166 2280 -1160 2320
rect -78 2320 -32 2332
rect -78 2280 -72 2320
rect -1166 2190 -72 2280
rect -1166 2152 -1160 2190
rect -1206 2140 -1160 2152
rect -78 2152 -72 2190
rect -38 2280 -32 2320
rect 30 2320 76 2332
rect 30 2280 36 2320
rect -38 2190 36 2280
rect -38 2152 -32 2190
rect -78 2140 -32 2152
rect 30 2152 36 2190
rect 70 2280 76 2320
rect 1158 2320 1204 2332
rect 1158 2280 1164 2320
rect 70 2190 1164 2280
rect 70 2152 76 2190
rect 30 2140 76 2152
rect 1158 2152 1164 2190
rect 1198 2280 1204 2320
rect 1266 2320 1312 2332
rect 1266 2280 1272 2320
rect 1198 2190 1272 2280
rect 1198 2152 1204 2190
rect 1158 2140 1204 2152
rect 1266 2152 1272 2190
rect 1306 2280 1312 2320
rect 2394 2320 2440 2332
rect 2394 2280 2400 2320
rect 1306 2270 2400 2280
rect 1306 2200 1460 2270
rect 1530 2200 1700 2270
rect 1770 2200 2400 2270
rect 1306 2190 2400 2200
rect 1306 2152 1312 2190
rect 1266 2140 1312 2152
rect 2394 2152 2400 2190
rect 2434 2280 2440 2320
rect 2502 2320 2548 2332
rect 2502 2280 2508 2320
rect 2434 2190 2508 2280
rect 2434 2152 2440 2190
rect 2394 2140 2440 2152
rect 2502 2152 2508 2190
rect 2542 2280 2548 2320
rect 3630 2320 3676 2332
rect 3630 2280 3636 2320
rect 2542 2190 3636 2280
rect 2542 2152 2548 2190
rect 2502 2140 2548 2152
rect 3630 2152 3636 2190
rect 3670 2152 3676 2320
rect 3630 2140 3676 2152
rect -3600 2124 -2591 2130
rect -3600 2090 -3579 2124
rect -2603 2110 -2591 2124
rect -2355 2124 -1355 2130
rect -2355 2110 -2343 2124
rect -2603 2090 -2343 2110
rect -1367 2110 -1355 2124
rect -1119 2124 -119 2130
rect -1119 2110 -1107 2124
rect -131 2110 -119 2124
rect 117 2124 1117 2130
rect 117 2110 129 2124
rect 1105 2110 1117 2124
rect 1353 2124 2353 2130
rect 1353 2110 1365 2124
rect -1367 2090 -1107 2110
rect -131 2090 129 2110
rect 1105 2090 1365 2110
rect 2341 2110 2353 2124
rect 2589 2124 3594 2130
rect 2589 2110 2601 2124
rect 2341 2090 2601 2110
rect 3577 2090 3594 2124
rect -3600 2040 -560 2090
rect -490 2040 -450 2090
rect -380 2040 380 2090
rect 450 2040 490 2090
rect 560 2040 3594 2090
rect -3600 2030 3594 2040
rect -920 1592 900 1620
rect -920 1558 -818 1592
rect -592 1558 -350 1592
rect -124 1558 118 1592
rect 344 1558 586 1592
rect 812 1558 900 1592
rect -920 1550 900 1558
rect -920 1540 380 1550
rect -920 1530 -560 1540
rect -920 1470 -902 1530
rect -908 1362 -902 1470
rect -868 1470 -560 1530
rect -490 1470 -450 1540
rect -380 1530 380 1540
rect -380 1470 -74 1530
rect -868 1390 -542 1470
rect -868 1362 -862 1390
rect -908 1350 -862 1362
rect -550 1362 -542 1390
rect -508 1362 -434 1470
rect -400 1390 -74 1470
rect -400 1362 -390 1390
rect -550 1350 -390 1362
rect -80 1362 -74 1390
rect -40 1362 34 1530
rect 68 1480 380 1530
rect 450 1480 490 1550
rect 560 1542 900 1550
rect 560 1530 902 1542
rect 560 1480 862 1530
rect 68 1390 394 1480
rect 68 1362 75 1390
rect -80 1350 75 1362
rect 388 1362 394 1390
rect 428 1362 502 1480
rect 536 1390 862 1480
rect 536 1362 545 1390
rect 388 1350 545 1362
rect 856 1362 862 1390
rect 896 1362 902 1530
rect 856 1350 902 1362
rect -830 1334 -580 1340
rect -830 1320 -818 1334
rect -840 1300 -818 1320
rect -592 1320 -580 1334
rect -362 1334 -112 1340
rect -362 1320 -350 1334
rect -592 1300 -350 1320
rect -124 1320 -112 1334
rect 106 1334 356 1340
rect 106 1320 118 1334
rect -124 1300 118 1320
rect 344 1320 356 1334
rect 574 1334 824 1340
rect 574 1320 586 1334
rect 344 1300 586 1320
rect 812 1320 824 1334
rect 812 1300 830 1320
rect -840 1280 830 1300
rect -840 1226 870 1280
rect -852 1220 882 1226
rect -852 1070 -840 1220
rect -620 1210 -320 1220
rect -620 1070 -608 1210
rect -852 1064 -608 1070
rect -332 1070 -320 1210
rect -100 1210 100 1220
rect -100 1070 -88 1210
rect -332 1064 -88 1070
rect 88 1070 100 1210
rect 320 1210 650 1220
rect 320 1070 332 1210
rect 88 1064 332 1070
rect 638 1070 650 1210
rect 870 1070 882 1220
rect 638 1064 882 1070
rect 1440 1030 1790 1050
rect -1740 1010 1460 1030
rect -1740 940 -1720 1010
rect -1650 940 -1510 1010
rect -1440 967 1460 1010
rect -1440 940 -598 967
rect -1740 933 -598 940
rect -122 933 120 967
rect 596 960 1460 967
rect 1530 960 1700 1030
rect 1770 960 1790 1030
rect 596 940 1790 960
rect 596 933 1460 940
rect -1740 920 1460 933
rect -1740 850 -1720 920
rect -1650 850 -1510 920
rect -1440 905 1460 920
rect -1440 850 -682 905
rect -1740 820 -1410 850
rect -688 837 -682 850
rect -648 850 -72 905
rect -648 837 -642 850
rect -688 825 -642 837
rect -78 837 -72 850
rect -38 850 36 905
rect -38 837 -32 850
rect -78 825 -32 837
rect 30 837 36 850
rect 70 850 646 905
rect 70 837 76 850
rect 30 825 76 837
rect 640 837 646 850
rect 680 870 1460 905
rect 1530 870 1700 940
rect 1770 870 1790 940
rect 680 850 1790 870
rect 680 837 686 850
rect 640 825 686 837
rect -610 809 -110 815
rect -610 795 -598 809
rect -615 780 -598 795
rect -122 795 -110 809
rect 108 809 608 815
rect 108 795 120 809
rect -620 775 -598 780
rect -122 775 120 795
rect 596 795 608 809
rect 596 780 620 795
rect 596 775 630 780
rect -620 720 -560 775
rect -490 720 -450 775
rect -380 720 380 775
rect 450 720 490 775
rect 560 720 630 775
rect -620 710 630 720
rect -1092 670 -888 676
rect -3212 660 -3008 666
rect -3212 530 -3200 660
rect -3020 530 -3008 660
rect -3212 524 -3008 530
rect -2072 660 -1868 666
rect -2072 530 -2060 660
rect -1880 530 -1868 660
rect -1092 540 -1080 670
rect -900 540 -888 670
rect -1092 534 -888 540
rect -322 670 -118 676
rect -322 540 -310 670
rect -130 540 -118 670
rect -322 534 -118 540
rect 118 670 322 676
rect 118 540 130 670
rect 310 540 322 670
rect 1908 670 2112 676
rect 118 534 322 540
rect 838 660 1042 666
rect -2072 524 -1868 530
rect 838 530 850 660
rect 1030 530 1042 660
rect 1908 540 1920 670
rect 2100 540 2112 670
rect 1908 534 2112 540
rect 2908 670 3112 676
rect 2908 540 2920 670
rect 3100 540 3112 670
rect 2908 534 3112 540
rect 838 524 1042 530
rect -3550 490 3540 495
rect -3550 442 -1720 490
rect -1650 442 -1500 490
rect -1430 442 1460 490
rect 1530 442 1700 490
rect 1770 448 3540 490
rect 1770 442 3545 448
rect -3550 420 -3533 442
rect -3545 408 -3533 420
rect -2557 420 -2315 442
rect -1339 420 -1097 442
rect -2557 408 -2545 420
rect -3545 402 -2545 408
rect -2327 408 -2315 420
rect -1339 408 -1327 420
rect -2327 402 -1327 408
rect -1109 408 -1097 420
rect -121 420 121 442
rect -121 408 -109 420
rect -1109 402 -109 408
rect 109 408 121 420
rect 1097 420 1339 442
rect 2315 420 2557 442
rect 1097 408 1109 420
rect 109 402 1109 408
rect 1327 408 1339 420
rect 2315 408 2327 420
rect 1327 402 2327 408
rect 2545 408 2557 420
rect 3533 408 3545 442
rect 2545 402 3545 408
rect -3623 380 -3577 392
rect -3623 212 -3617 380
rect -3583 345 -3577 380
rect -2513 380 -2467 392
rect -2513 345 -2507 380
rect -3583 260 -2507 345
rect -3583 212 -3577 260
rect -3623 200 -3577 212
rect -2513 212 -2507 260
rect -2473 345 -2467 380
rect -2405 380 -2359 392
rect -2405 345 -2399 380
rect -2473 260 -2399 345
rect -2473 212 -2467 260
rect -2513 200 -2467 212
rect -2405 212 -2399 260
rect -2365 345 -2359 380
rect -1295 380 -1249 392
rect -1295 345 -1289 380
rect -2365 260 -1289 345
rect -2365 212 -2359 260
rect -2405 200 -2359 212
rect -1295 212 -1289 260
rect -1255 345 -1249 380
rect -1187 380 -1141 392
rect -1187 345 -1181 380
rect -1255 260 -1181 345
rect -1255 212 -1249 260
rect -1295 200 -1249 212
rect -1187 212 -1181 260
rect -1147 345 -1141 380
rect -77 380 -31 392
rect -77 345 -71 380
rect -1147 340 -71 345
rect -1147 270 -560 340
rect -490 270 -450 340
rect -380 270 -71 340
rect -1147 260 -71 270
rect -1147 212 -1141 260
rect -1187 200 -1141 212
rect -77 212 -71 260
rect -37 345 -31 380
rect 31 380 77 392
rect 31 345 37 380
rect -37 260 37 345
rect -37 212 -31 260
rect -77 200 -31 212
rect 31 212 37 260
rect 71 345 77 380
rect 1141 380 1187 392
rect 1141 345 1147 380
rect 71 340 1147 345
rect 71 270 380 340
rect 450 270 490 340
rect 560 270 1147 340
rect 71 260 1147 270
rect 71 212 77 260
rect 31 200 77 212
rect 1141 212 1147 260
rect 1181 345 1187 380
rect 1249 380 1295 392
rect 1249 345 1255 380
rect 1181 260 1255 345
rect 1181 212 1187 260
rect 1141 200 1187 212
rect 1249 212 1255 260
rect 1289 345 1295 380
rect 2359 380 2405 392
rect 2359 345 2365 380
rect 1289 260 2365 345
rect 1289 212 1295 260
rect 1249 200 1295 212
rect 2359 212 2365 260
rect 2399 345 2405 380
rect 2467 380 2513 392
rect 2467 345 2473 380
rect 2399 260 2473 345
rect 2399 212 2405 260
rect 2359 200 2405 212
rect 2467 212 2473 260
rect 2507 345 2513 380
rect 3577 380 3623 392
rect 3577 345 3583 380
rect 2507 260 3583 345
rect 2507 212 2513 260
rect 2467 200 2513 212
rect 3577 212 3583 260
rect 3617 212 3623 380
rect 3577 200 3623 212
rect -3545 184 -2545 190
rect -3545 170 -3533 184
rect -3550 150 -3533 170
rect -2557 170 -2545 184
rect -2327 184 -1327 190
rect -2327 170 -2315 184
rect -2557 150 -2315 170
rect -1339 170 -1327 184
rect -1109 184 -109 190
rect -1109 170 -1097 184
rect -1339 150 -1097 170
rect -121 170 -109 184
rect 109 184 1109 190
rect 109 170 121 184
rect -121 150 121 170
rect 1097 170 1109 184
rect 1327 184 2327 190
rect 1327 170 1339 184
rect 1097 150 1339 170
rect 2315 170 2327 184
rect 2545 184 3545 190
rect 2545 170 2557 184
rect 2315 150 2557 170
rect 3533 150 3545 184
rect -3550 144 3545 150
rect -3550 95 3540 144
rect -2200 -200 -1800 95
rect -800 -200 -400 95
rect 500 -200 900 95
rect 1790 -200 2200 95
rect -3000 -308 3000 -200
rect -3000 -314 203 -308
rect -3000 -711 -2827 -314
rect -1713 -711 -1307 -314
rect -193 -705 203 -314
rect 1317 -705 1713 -308
rect 2827 -705 3000 -308
rect -193 -711 3000 -705
rect -3000 -800 3000 -711
rect -3252 -1240 -3108 -1234
rect -3252 -1360 -3240 -1240
rect -3120 -1360 -3108 -1240
rect -3252 -1366 -3108 -1360
rect 3118 -1240 3262 -1234
rect 3118 -1360 3130 -1240
rect 3250 -1360 3262 -1240
rect 3118 -1366 3262 -1360
rect -3252 -4240 -3108 -4234
rect -3252 -4360 -3240 -4240
rect -3120 -4360 -3108 -4240
rect -3252 -4366 -3108 -4360
rect 3118 -4240 3262 -4234
rect 3118 -4360 3130 -4240
rect 3250 -4360 3262 -4240
rect 3118 -4366 3262 -4360
rect -3252 -7240 -3108 -7234
rect -3252 -7360 -3240 -7240
rect -3120 -7360 -3108 -7240
rect -3252 -7366 -3108 -7360
rect 3118 -7240 3262 -7234
rect 3118 -7360 3130 -7240
rect 3250 -7360 3262 -7240
rect 3118 -7366 3262 -7360
rect -3252 -10240 -3108 -10234
rect -3252 -10360 -3240 -10240
rect -3120 -10360 -3108 -10240
rect -3252 -10366 -3108 -10360
rect 3118 -10240 3262 -10234
rect 3118 -10360 3130 -10240
rect 3250 -10360 3262 -10240
rect 3118 -10366 3262 -10360
rect -3252 -13240 -3108 -13234
rect -3252 -13360 -3240 -13240
rect -3120 -13360 -3108 -13240
rect -3252 -13366 -3108 -13360
rect 3118 -13240 3262 -13234
rect 3118 -13360 3130 -13240
rect 3250 -13360 3262 -13240
rect 3118 -13366 3262 -13360
rect -3000 -14539 3000 -14500
rect -3000 -14545 203 -14539
rect -3000 -14570 -2827 -14545
rect -1713 -14570 -1307 -14545
rect -193 -14570 203 -14545
rect 1317 -14560 1713 -14539
rect 2827 -14560 3000 -14539
rect 1317 -14570 1690 -14560
rect -3000 -14980 -2860 -14570
rect -1690 -14980 -1350 -14570
rect -180 -14980 170 -14570
rect 1340 -14970 1690 -14570
rect 2860 -14970 3000 -14560
rect 1340 -14980 3000 -14970
rect -3000 -15000 3000 -14980
<< via1 >>
rect -3220 3020 -3060 3180
rect -2160 3020 -2000 3180
rect -700 3020 -540 3180
rect 520 3020 680 3180
rect 2000 3020 2160 3180
rect 3000 3020 3160 3180
rect -1720 2790 -1650 2860
rect -1500 2790 -1430 2860
rect 1460 2790 1530 2860
rect 1700 2790 1770 2860
rect -3220 2440 -3060 2600
rect -2160 2440 -2000 2600
rect -700 2440 -540 2600
rect 520 2440 680 2600
rect 2000 2440 2160 2600
rect 3000 2440 3160 2600
rect -1720 2200 -1650 2270
rect -1500 2200 -1430 2270
rect 1460 2200 1530 2270
rect 1700 2200 1770 2270
rect -560 2090 -490 2110
rect -450 2090 -380 2110
rect 380 2090 450 2110
rect 490 2090 560 2110
rect -560 2040 -490 2090
rect -450 2040 -380 2090
rect 380 2040 450 2090
rect 490 2040 560 2090
rect -560 1530 -490 1540
rect -560 1470 -542 1530
rect -542 1470 -508 1530
rect -508 1470 -490 1530
rect -450 1530 -380 1540
rect 380 1530 450 1550
rect -450 1470 -434 1530
rect -434 1470 -400 1530
rect -400 1470 -380 1530
rect 380 1480 394 1530
rect 394 1480 428 1530
rect 428 1480 450 1530
rect 490 1530 560 1550
rect 490 1480 502 1530
rect 502 1480 536 1530
rect 536 1480 560 1530
rect -840 1070 -620 1220
rect -320 1070 -100 1220
rect 100 1070 320 1220
rect 650 1070 870 1220
rect -1720 940 -1650 1010
rect -1510 940 -1440 1010
rect 1460 960 1530 1030
rect 1700 960 1770 1030
rect -1720 850 -1650 920
rect -1510 850 -1440 920
rect 1460 870 1530 940
rect 1700 870 1770 940
rect -560 775 -490 790
rect -450 775 -380 790
rect 380 775 450 790
rect 490 775 560 790
rect -560 720 -490 775
rect -450 720 -380 775
rect 380 720 450 775
rect 490 720 560 775
rect -3200 530 -3020 660
rect -2060 530 -1880 660
rect -1080 540 -900 670
rect -310 540 -130 670
rect 130 540 310 670
rect 850 530 1030 660
rect 1920 540 2100 670
rect 2920 540 3100 670
rect -1720 442 -1650 490
rect -1500 442 -1430 490
rect 1460 442 1530 490
rect 1700 442 1770 490
rect -1720 420 -1650 442
rect -1500 420 -1430 442
rect 1460 420 1530 442
rect 1700 420 1770 442
rect -560 270 -490 340
rect -450 270 -380 340
rect 380 270 450 340
rect 490 270 560 340
rect -3240 -1360 -3120 -1240
rect 3130 -1360 3250 -1240
rect -3240 -4360 -3120 -4240
rect 3130 -4360 3250 -4240
rect -3240 -7360 -3120 -7240
rect 3130 -7360 3250 -7240
rect -3240 -10360 -3120 -10240
rect 3130 -10360 3250 -10240
rect -3240 -13360 -3120 -13240
rect 3130 -13360 3250 -13240
rect -2860 -14942 -2827 -14570
rect -2827 -14942 -1713 -14570
rect -1713 -14942 -1690 -14570
rect -2860 -14980 -1690 -14942
rect -1350 -14942 -1307 -14570
rect -1307 -14942 -193 -14570
rect -193 -14942 -180 -14570
rect -1350 -14980 -180 -14942
rect 170 -14936 203 -14570
rect 203 -14936 1317 -14570
rect 1317 -14936 1340 -14570
rect 170 -14980 1340 -14936
rect 1690 -14936 1713 -14560
rect 1713 -14936 2827 -14560
rect 2827 -14936 2860 -14560
rect 1690 -14970 2860 -14936
<< metal2 >>
rect -3220 3180 -3060 3190
rect -3220 3010 -3060 3020
rect -2160 3180 -2000 3190
rect -2160 3010 -2000 3020
rect -700 3180 -540 3190
rect -700 3010 -540 3020
rect 520 3180 680 3190
rect 520 3010 680 3020
rect 2000 3180 2160 3190
rect 2000 3010 2160 3020
rect 3000 3180 3160 3190
rect 3000 3010 3160 3020
rect 1440 2860 1790 2870
rect -1740 2790 -1720 2860
rect -1650 2790 -1500 2860
rect -1430 2790 -1410 2860
rect -3220 2600 -3060 2610
rect -3220 2430 -3060 2440
rect -2160 2600 -2000 2610
rect -2160 2430 -2000 2440
rect -1740 2270 -1410 2790
rect 1440 2790 1460 2860
rect 1530 2790 1700 2860
rect 1770 2790 1790 2860
rect -700 2600 -540 2610
rect -700 2430 -540 2440
rect 520 2600 680 2610
rect 520 2430 680 2440
rect -1740 2200 -1720 2270
rect -1650 2200 -1500 2270
rect -1430 2200 -1410 2270
rect -1740 1010 -1410 2200
rect 1440 2270 1790 2790
rect 2000 2600 2160 2610
rect 2000 2430 2160 2440
rect 3000 2600 3160 2610
rect 3000 2430 3160 2440
rect 1440 2200 1460 2270
rect 1530 2200 1700 2270
rect 1770 2200 1790 2270
rect -580 2110 -360 2120
rect -580 2040 -560 2110
rect -490 2040 -450 2110
rect -380 2040 -360 2110
rect -580 1540 -360 2040
rect -580 1470 -560 1540
rect -490 1470 -450 1540
rect -380 1470 -360 1540
rect -840 1220 -620 1230
rect -840 1060 -620 1070
rect -1740 940 -1720 1010
rect -1650 940 -1510 1010
rect -1440 940 -1410 1010
rect -1740 920 -1410 940
rect -1740 850 -1720 920
rect -1650 850 -1510 920
rect -1440 850 -1410 920
rect -3200 660 -3020 670
rect -3200 520 -3020 530
rect -2060 660 -1880 670
rect -2060 520 -1880 530
rect -1740 490 -1410 850
rect -580 790 -360 1470
rect 360 2110 580 2130
rect 360 2040 380 2110
rect 450 2040 490 2110
rect 560 2040 580 2110
rect 360 1550 580 2040
rect 360 1480 380 1550
rect 450 1480 490 1550
rect 560 1480 580 1550
rect -320 1220 -100 1230
rect -320 1060 -100 1070
rect 100 1220 320 1230
rect 100 1060 320 1070
rect -580 720 -560 790
rect -490 720 -450 790
rect -380 720 -360 790
rect -1080 670 -900 680
rect -1080 530 -900 540
rect -1740 420 -1720 490
rect -1650 420 -1500 490
rect -1430 420 -1410 490
rect -1740 410 -1410 420
rect -580 340 -360 720
rect 360 790 580 1480
rect 650 1220 870 1230
rect 650 1060 870 1070
rect 360 720 380 790
rect 450 720 490 790
rect 560 720 580 790
rect -310 670 -130 680
rect -310 530 -130 540
rect 130 670 310 680
rect 130 530 310 540
rect -580 270 -560 340
rect -490 270 -450 340
rect -380 270 -360 340
rect -580 200 -360 270
rect 360 340 580 720
rect 1440 1030 1790 2200
rect 1440 960 1460 1030
rect 1530 960 1700 1030
rect 1770 960 1790 1030
rect 1440 940 1790 960
rect 1440 870 1460 940
rect 1530 870 1700 940
rect 1770 870 1790 940
rect 850 660 1030 670
rect 850 520 1030 530
rect 1440 490 1790 870
rect 1920 670 2100 680
rect 1920 530 2100 540
rect 2920 670 3100 680
rect 2920 530 3100 540
rect 1440 420 1460 490
rect 1530 420 1700 490
rect 1770 420 1790 490
rect 1440 390 1790 420
rect 360 270 380 340
rect 450 270 490 340
rect 560 270 580 340
rect 360 210 580 270
rect -3240 -1240 -3120 -1230
rect -3240 -1370 -3120 -1360
rect 3130 -1240 3250 -1230
rect 3130 -1370 3250 -1360
rect -3240 -4240 -3120 -4230
rect -3240 -4370 -3120 -4360
rect 3130 -4240 3250 -4230
rect 3130 -4370 3250 -4360
rect -3240 -7240 -3120 -7230
rect -3240 -7370 -3120 -7360
rect 3130 -7240 3250 -7230
rect 3130 -7370 3250 -7360
rect -3240 -10240 -3120 -10230
rect -3240 -10370 -3120 -10360
rect 3130 -10240 3250 -10230
rect 3130 -10370 3250 -10360
rect -3240 -13240 -3120 -13230
rect -3240 -13370 -3120 -13360
rect 3130 -13240 3250 -13230
rect 3130 -13370 3250 -13360
rect 1690 -14560 2860 -14550
rect -2860 -14570 -1690 -14560
rect -2860 -14990 -1690 -14980
rect -1350 -14570 -180 -14560
rect -1350 -14990 -180 -14980
rect 170 -14570 1340 -14560
rect 1690 -14980 2860 -14970
rect 170 -14990 1340 -14980
<< via2 >>
rect -3220 3020 -3060 3180
rect -2160 3020 -2000 3180
rect -700 3020 -540 3180
rect 520 3020 680 3180
rect 2000 3020 2160 3180
rect 3000 3020 3160 3180
rect -3220 2440 -3060 2600
rect -2160 2440 -2000 2600
rect -700 2440 -540 2600
rect 520 2440 680 2600
rect 2000 2440 2160 2600
rect 3000 2440 3160 2600
rect -840 1070 -620 1220
rect -3200 530 -3020 660
rect -2060 530 -1880 660
rect -320 1070 -100 1220
rect 100 1070 320 1220
rect -1080 540 -900 670
rect 650 1070 870 1220
rect -310 540 -130 670
rect 130 540 310 670
rect 850 530 1030 660
rect 1920 540 2100 670
rect 2920 540 3100 670
rect -3240 -1360 -3120 -1240
rect 3130 -1360 3250 -1240
rect -3240 -4360 -3120 -4240
rect 3130 -4360 3250 -4240
rect -3240 -7360 -3120 -7240
rect 3130 -7360 3250 -7240
rect -3240 -10360 -3120 -10240
rect 3130 -10360 3250 -10240
rect -3240 -13360 -3120 -13240
rect 3130 -13360 3250 -13240
rect -2860 -14980 -1690 -14570
rect -1350 -14980 -180 -14570
rect 170 -14980 1340 -14570
rect 1690 -14970 2860 -14560
<< metal3 >>
rect -3260 3180 3200 3640
rect -3260 3020 -3220 3180
rect -3060 3020 -2160 3180
rect -2000 3020 -700 3180
rect -540 3020 520 3180
rect 680 3020 2000 3180
rect 2160 3020 3000 3180
rect 3160 3020 3200 3180
rect -3260 2600 3200 3020
rect -3260 2440 -3220 2600
rect -3060 2440 -2160 2600
rect -2000 2440 -700 2600
rect -540 2440 520 2600
rect 680 2440 2000 2600
rect 2160 2440 3000 2600
rect 3160 2440 3200 2600
rect -3260 2420 3200 2440
rect -3710 1220 3310 1260
rect -3710 1080 -840 1220
rect -3310 1070 -840 1080
rect -620 1070 -320 1220
rect -100 1070 100 1220
rect 320 1070 650 1220
rect 870 1070 3310 1220
rect -3310 670 3310 1070
rect -3310 660 -1080 670
rect -3310 530 -3200 660
rect -3020 530 -2060 660
rect -1880 540 -1080 660
rect -900 540 -310 670
rect -130 540 130 670
rect 310 660 1920 670
rect 310 540 850 660
rect -1880 530 850 540
rect 1030 540 1920 660
rect 2100 540 2920 670
rect 3100 540 3310 670
rect 1030 530 3310 540
rect -3310 500 3310 530
rect -3310 -1240 -2990 500
rect -3310 -1360 -3240 -1240
rect -3120 -1360 -2990 -1240
rect -3310 -4240 -2990 -1360
rect -3310 -4360 -3240 -4240
rect -3120 -4360 -2990 -4240
rect -3310 -7240 -2990 -4360
rect -3310 -7360 -3240 -7240
rect -3120 -7360 -2990 -7240
rect -3310 -10240 -2990 -7360
rect -3310 -10360 -3240 -10240
rect -3120 -10360 -2990 -10240
rect -3310 -13240 -2990 -10360
rect -3310 -13360 -3240 -13240
rect -3120 -13360 -2990 -13240
rect -3310 -14540 -2990 -13360
rect 2990 -1240 3310 500
rect 2990 -1360 3130 -1240
rect 3250 -1360 3310 -1240
rect 2990 -4240 3310 -1360
rect 2990 -4360 3130 -4240
rect 3250 -4360 3310 -4240
rect 2990 -7240 3310 -4360
rect 2990 -7360 3130 -7240
rect 3250 -7360 3310 -7240
rect 2990 -10240 3310 -7360
rect 2990 -10360 3130 -10240
rect 3250 -10360 3310 -10240
rect 2990 -13240 3310 -10360
rect 2990 -13360 3130 -13240
rect 3250 -13360 3310 -13240
rect 2990 -14540 3310 -13360
rect -3310 -14560 3310 -14540
rect -3310 -14570 1690 -14560
rect -3310 -14980 -2860 -14570
rect -1690 -14980 -1350 -14570
rect -180 -14980 170 -14570
rect 1340 -14970 1690 -14570
rect 2860 -14970 3310 -14560
rect 1340 -14980 3310 -14970
rect -3310 -15020 3310 -14980
<< res5p73 >>
rect -2845 -14530 -1695 -726
rect -1325 -14530 -175 -726
rect 185 -14524 1335 -720
rect 1695 -14524 2845 -720
<< end >>
