magic
tech sky130A
magscale 1 2
timestamp 1683391037
<< pwell >>
rect -720 -710 720 710
<< nmos >>
rect -524 -500 -424 500
rect -366 -500 -266 500
rect -208 -500 -108 500
rect -50 -500 50 500
rect 108 -500 208 500
rect 266 -500 366 500
rect 424 -500 524 500
<< ndiff >>
rect -582 488 -524 500
rect -582 -488 -570 488
rect -536 -488 -524 488
rect -582 -500 -524 -488
rect -424 488 -366 500
rect -424 -488 -412 488
rect -378 -488 -366 488
rect -424 -500 -366 -488
rect -266 488 -208 500
rect -266 -488 -254 488
rect -220 -488 -208 488
rect -266 -500 -208 -488
rect -108 488 -50 500
rect -108 -488 -96 488
rect -62 -488 -50 488
rect -108 -500 -50 -488
rect 50 488 108 500
rect 50 -488 62 488
rect 96 -488 108 488
rect 50 -500 108 -488
rect 208 488 266 500
rect 208 -488 220 488
rect 254 -488 266 488
rect 208 -500 266 -488
rect 366 488 424 500
rect 366 -488 378 488
rect 412 -488 424 488
rect 366 -500 424 -488
rect 524 488 582 500
rect 524 -488 536 488
rect 570 -488 582 488
rect 524 -500 582 -488
<< ndiffc >>
rect -570 -488 -536 488
rect -412 -488 -378 488
rect -254 -488 -220 488
rect -96 -488 -62 488
rect 62 -488 96 488
rect 220 -488 254 488
rect 378 -488 412 488
rect 536 -488 570 488
<< psubdiff >>
rect -684 640 -588 674
rect 588 640 684 674
rect -684 578 -650 640
rect 650 578 684 640
rect -684 -640 -650 -578
rect 650 -640 684 -578
rect -684 -674 -588 -640
rect 588 -674 684 -640
<< psubdiffcont >>
rect -588 640 588 674
rect -684 -578 -650 578
rect 650 -578 684 578
rect -588 -674 588 -640
<< poly >>
rect -524 572 -424 588
rect -524 538 -508 572
rect -440 538 -424 572
rect -524 500 -424 538
rect -366 572 -266 588
rect -366 538 -350 572
rect -282 538 -266 572
rect -366 500 -266 538
rect -208 572 -108 588
rect -208 538 -192 572
rect -124 538 -108 572
rect -208 500 -108 538
rect -50 572 50 588
rect -50 538 -34 572
rect 34 538 50 572
rect -50 500 50 538
rect 108 572 208 588
rect 108 538 124 572
rect 192 538 208 572
rect 108 500 208 538
rect 266 572 366 588
rect 266 538 282 572
rect 350 538 366 572
rect 266 500 366 538
rect 424 572 524 588
rect 424 538 440 572
rect 508 538 524 572
rect 424 500 524 538
rect -524 -538 -424 -500
rect -524 -572 -508 -538
rect -440 -572 -424 -538
rect -524 -588 -424 -572
rect -366 -538 -266 -500
rect -366 -572 -350 -538
rect -282 -572 -266 -538
rect -366 -588 -266 -572
rect -208 -538 -108 -500
rect -208 -572 -192 -538
rect -124 -572 -108 -538
rect -208 -588 -108 -572
rect -50 -538 50 -500
rect -50 -572 -34 -538
rect 34 -572 50 -538
rect -50 -588 50 -572
rect 108 -538 208 -500
rect 108 -572 124 -538
rect 192 -572 208 -538
rect 108 -588 208 -572
rect 266 -538 366 -500
rect 266 -572 282 -538
rect 350 -572 366 -538
rect 266 -588 366 -572
rect 424 -538 524 -500
rect 424 -572 440 -538
rect 508 -572 524 -538
rect 424 -588 524 -572
<< polycont >>
rect -508 538 -440 572
rect -350 538 -282 572
rect -192 538 -124 572
rect -34 538 34 572
rect 124 538 192 572
rect 282 538 350 572
rect 440 538 508 572
rect -508 -572 -440 -538
rect -350 -572 -282 -538
rect -192 -572 -124 -538
rect -34 -572 34 -538
rect 124 -572 192 -538
rect 282 -572 350 -538
rect 440 -572 508 -538
<< locali >>
rect -684 640 -588 674
rect 588 640 684 674
rect -684 578 -650 640
rect 650 578 684 640
rect -524 538 -508 572
rect -440 538 -424 572
rect -366 538 -350 572
rect -282 538 -266 572
rect -208 538 -192 572
rect -124 538 -108 572
rect -50 538 -34 572
rect 34 538 50 572
rect 108 538 124 572
rect 192 538 208 572
rect 266 538 282 572
rect 350 538 366 572
rect 424 538 440 572
rect 508 538 524 572
rect -570 488 -536 504
rect -570 -504 -536 -488
rect -412 488 -378 504
rect -412 -504 -378 -488
rect -254 488 -220 504
rect -254 -504 -220 -488
rect -96 488 -62 504
rect -96 -504 -62 -488
rect 62 488 96 504
rect 62 -504 96 -488
rect 220 488 254 504
rect 220 -504 254 -488
rect 378 488 412 504
rect 378 -504 412 -488
rect 536 488 570 504
rect 536 -504 570 -488
rect -524 -572 -508 -538
rect -440 -572 -424 -538
rect -366 -572 -350 -538
rect -282 -572 -266 -538
rect -208 -572 -192 -538
rect -124 -572 -108 -538
rect -50 -572 -34 -538
rect 34 -572 50 -538
rect 108 -572 124 -538
rect 192 -572 208 -538
rect 266 -572 282 -538
rect 350 -572 366 -538
rect 424 -572 440 -538
rect 508 -572 524 -538
rect -684 -640 -650 -578
rect 650 -640 684 -578
rect -684 -674 -588 -640
rect 588 -674 684 -640
<< viali >>
rect -325 640 325 674
rect -508 538 -440 572
rect -350 538 -282 572
rect -192 538 -124 572
rect -34 538 34 572
rect 124 538 192 572
rect 282 538 350 572
rect 440 538 508 572
rect -570 -488 -536 488
rect -412 -488 -378 488
rect -254 -488 -220 488
rect -96 -488 -62 488
rect 62 -488 96 488
rect 220 -488 254 488
rect 378 -488 412 488
rect 536 -488 570 488
rect -508 -572 -440 -538
rect -350 -572 -282 -538
rect -192 -572 -124 -538
rect -34 -572 34 -538
rect 124 -572 192 -538
rect 282 -572 350 -538
rect 440 -572 508 -538
rect -325 -674 325 -640
<< metal1 >>
rect -337 674 337 680
rect -337 640 -325 674
rect 325 640 337 674
rect -337 634 337 640
rect -520 572 -428 578
rect -520 538 -508 572
rect -440 538 -428 572
rect -520 532 -428 538
rect -362 572 -270 578
rect -362 538 -350 572
rect -282 538 -270 572
rect -362 532 -270 538
rect -204 572 -112 578
rect -204 538 -192 572
rect -124 538 -112 572
rect -204 532 -112 538
rect -46 572 46 578
rect -46 538 -34 572
rect 34 538 46 572
rect -46 532 46 538
rect 112 572 204 578
rect 112 538 124 572
rect 192 538 204 572
rect 112 532 204 538
rect 270 572 362 578
rect 270 538 282 572
rect 350 538 362 572
rect 270 532 362 538
rect 428 572 520 578
rect 428 538 440 572
rect 508 538 520 572
rect 428 532 520 538
rect -576 488 -530 500
rect -576 -488 -570 488
rect -536 -488 -530 488
rect -576 -500 -530 -488
rect -418 488 -372 500
rect -418 -488 -412 488
rect -378 -488 -372 488
rect -418 -500 -372 -488
rect -260 488 -214 500
rect -260 -488 -254 488
rect -220 -488 -214 488
rect -260 -500 -214 -488
rect -102 488 -56 500
rect -102 -488 -96 488
rect -62 -488 -56 488
rect -102 -500 -56 -488
rect 56 488 102 500
rect 56 -488 62 488
rect 96 -488 102 488
rect 56 -500 102 -488
rect 214 488 260 500
rect 214 -488 220 488
rect 254 -488 260 488
rect 214 -500 260 -488
rect 372 488 418 500
rect 372 -488 378 488
rect 412 -488 418 488
rect 372 -500 418 -488
rect 530 488 576 500
rect 530 -488 536 488
rect 570 -488 576 488
rect 530 -500 576 -488
rect -520 -538 -428 -532
rect -520 -572 -508 -538
rect -440 -572 -428 -538
rect -520 -578 -428 -572
rect -362 -538 -270 -532
rect -362 -572 -350 -538
rect -282 -572 -270 -538
rect -362 -578 -270 -572
rect -204 -538 -112 -532
rect -204 -572 -192 -538
rect -124 -572 -112 -538
rect -204 -578 -112 -572
rect -46 -538 46 -532
rect -46 -572 -34 -538
rect 34 -572 46 -538
rect -46 -578 46 -572
rect 112 -538 204 -532
rect 112 -572 124 -538
rect 192 -572 204 -538
rect 112 -578 204 -572
rect 270 -538 362 -532
rect 270 -572 282 -538
rect 350 -572 362 -538
rect 270 -578 362 -572
rect 428 -538 520 -532
rect 428 -572 440 -538
rect 508 -572 520 -538
rect 428 -578 520 -572
rect -337 -640 337 -634
rect -337 -674 -325 -640
rect 325 -674 337 -640
rect -337 -680 337 -674
<< properties >>
string FIXED_BBOX -667 -657 667 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.5 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 50 viagr 0 viagl 0 viagt 50
<< end >>
