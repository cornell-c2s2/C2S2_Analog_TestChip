magic
tech sky130A
magscale 1 2
timestamp 1683391037
<< nwell >>
rect -246 -4427 246 4427
<< pmos >>
rect -50 3208 50 4208
rect -50 1972 50 2972
rect -50 736 50 1736
rect -50 -500 50 500
rect -50 -1736 50 -736
rect -50 -2972 50 -1972
rect -50 -4208 50 -3208
<< pdiff >>
rect -108 4196 -50 4208
rect -108 3220 -96 4196
rect -62 3220 -50 4196
rect -108 3208 -50 3220
rect 50 4196 108 4208
rect 50 3220 62 4196
rect 96 3220 108 4196
rect 50 3208 108 3220
rect -108 2960 -50 2972
rect -108 1984 -96 2960
rect -62 1984 -50 2960
rect -108 1972 -50 1984
rect 50 2960 108 2972
rect 50 1984 62 2960
rect 96 1984 108 2960
rect 50 1972 108 1984
rect -108 1724 -50 1736
rect -108 748 -96 1724
rect -62 748 -50 1724
rect -108 736 -50 748
rect 50 1724 108 1736
rect 50 748 62 1724
rect 96 748 108 1724
rect 50 736 108 748
rect -108 488 -50 500
rect -108 -488 -96 488
rect -62 -488 -50 488
rect -108 -500 -50 -488
rect 50 488 108 500
rect 50 -488 62 488
rect 96 -488 108 488
rect 50 -500 108 -488
rect -108 -748 -50 -736
rect -108 -1724 -96 -748
rect -62 -1724 -50 -748
rect -108 -1736 -50 -1724
rect 50 -748 108 -736
rect 50 -1724 62 -748
rect 96 -1724 108 -748
rect 50 -1736 108 -1724
rect -108 -1984 -50 -1972
rect -108 -2960 -96 -1984
rect -62 -2960 -50 -1984
rect -108 -2972 -50 -2960
rect 50 -1984 108 -1972
rect 50 -2960 62 -1984
rect 96 -2960 108 -1984
rect 50 -2972 108 -2960
rect -108 -3220 -50 -3208
rect -108 -4196 -96 -3220
rect -62 -4196 -50 -3220
rect -108 -4208 -50 -4196
rect 50 -3220 108 -3208
rect 50 -4196 62 -3220
rect 96 -4196 108 -3220
rect 50 -4208 108 -4196
<< pdiffc >>
rect -96 3220 -62 4196
rect 62 3220 96 4196
rect -96 1984 -62 2960
rect 62 1984 96 2960
rect -96 748 -62 1724
rect 62 748 96 1724
rect -96 -488 -62 488
rect 62 -488 96 488
rect -96 -1724 -62 -748
rect 62 -1724 96 -748
rect -96 -2960 -62 -1984
rect 62 -2960 96 -1984
rect -96 -4196 -62 -3220
rect 62 -4196 96 -3220
<< nsubdiff >>
rect -210 4357 -114 4391
rect 114 4357 210 4391
rect -210 4295 -176 4357
rect 176 4295 210 4357
rect -210 -4357 -176 -4295
rect 176 -4357 210 -4295
rect -210 -4391 -114 -4357
rect 114 -4391 210 -4357
<< nsubdiffcont >>
rect -114 4357 114 4391
rect -210 -4295 -176 4295
rect 176 -4295 210 4295
rect -114 -4391 114 -4357
<< poly >>
rect -50 4289 50 4305
rect -50 4255 -34 4289
rect 34 4255 50 4289
rect -50 4208 50 4255
rect -50 3161 50 3208
rect -50 3127 -34 3161
rect 34 3127 50 3161
rect -50 3111 50 3127
rect -50 3053 50 3069
rect -50 3019 -34 3053
rect 34 3019 50 3053
rect -50 2972 50 3019
rect -50 1925 50 1972
rect -50 1891 -34 1925
rect 34 1891 50 1925
rect -50 1875 50 1891
rect -50 1817 50 1833
rect -50 1783 -34 1817
rect 34 1783 50 1817
rect -50 1736 50 1783
rect -50 689 50 736
rect -50 655 -34 689
rect 34 655 50 689
rect -50 639 50 655
rect -50 581 50 597
rect -50 547 -34 581
rect 34 547 50 581
rect -50 500 50 547
rect -50 -547 50 -500
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -50 -597 50 -581
rect -50 -655 50 -639
rect -50 -689 -34 -655
rect 34 -689 50 -655
rect -50 -736 50 -689
rect -50 -1783 50 -1736
rect -50 -1817 -34 -1783
rect 34 -1817 50 -1783
rect -50 -1833 50 -1817
rect -50 -1891 50 -1875
rect -50 -1925 -34 -1891
rect 34 -1925 50 -1891
rect -50 -1972 50 -1925
rect -50 -3019 50 -2972
rect -50 -3053 -34 -3019
rect 34 -3053 50 -3019
rect -50 -3069 50 -3053
rect -50 -3127 50 -3111
rect -50 -3161 -34 -3127
rect 34 -3161 50 -3127
rect -50 -3208 50 -3161
rect -50 -4255 50 -4208
rect -50 -4289 -34 -4255
rect 34 -4289 50 -4255
rect -50 -4305 50 -4289
<< polycont >>
rect -34 4255 34 4289
rect -34 3127 34 3161
rect -34 3019 34 3053
rect -34 1891 34 1925
rect -34 1783 34 1817
rect -34 655 34 689
rect -34 547 34 581
rect -34 -581 34 -547
rect -34 -689 34 -655
rect -34 -1817 34 -1783
rect -34 -1925 34 -1891
rect -34 -3053 34 -3019
rect -34 -3161 34 -3127
rect -34 -4289 34 -4255
<< locali >>
rect -210 4357 -114 4391
rect 114 4357 210 4391
rect -210 4295 -176 4357
rect 176 4295 210 4357
rect -50 4255 -34 4289
rect 34 4255 50 4289
rect -96 4196 -62 4212
rect -96 3204 -62 3220
rect 62 4196 96 4212
rect 62 3204 96 3220
rect -50 3127 -34 3161
rect 34 3127 50 3161
rect -50 3019 -34 3053
rect 34 3019 50 3053
rect -96 2960 -62 2976
rect -96 1968 -62 1984
rect 62 2960 96 2976
rect 62 1968 96 1984
rect -50 1891 -34 1925
rect 34 1891 50 1925
rect -50 1783 -34 1817
rect 34 1783 50 1817
rect -96 1724 -62 1740
rect -96 732 -62 748
rect 62 1724 96 1740
rect 62 732 96 748
rect -50 655 -34 689
rect 34 655 50 689
rect -50 547 -34 581
rect 34 547 50 581
rect -96 488 -62 504
rect -96 -504 -62 -488
rect 62 488 96 504
rect 62 -504 96 -488
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -50 -689 -34 -655
rect 34 -689 50 -655
rect -96 -748 -62 -732
rect -96 -1740 -62 -1724
rect 62 -748 96 -732
rect 62 -1740 96 -1724
rect -50 -1817 -34 -1783
rect 34 -1817 50 -1783
rect -50 -1925 -34 -1891
rect 34 -1925 50 -1891
rect -96 -1984 -62 -1968
rect -96 -2976 -62 -2960
rect 62 -1984 96 -1968
rect 62 -2976 96 -2960
rect -50 -3053 -34 -3019
rect 34 -3053 50 -3019
rect -50 -3161 -34 -3127
rect 34 -3161 50 -3127
rect -96 -3220 -62 -3204
rect -96 -4212 -62 -4196
rect 62 -3220 96 -3204
rect 62 -4212 96 -4196
rect -50 -4289 -34 -4255
rect 34 -4289 50 -4255
rect -210 -4357 -176 -4295
rect 176 -4357 210 -4295
rect -210 -4391 -114 -4357
rect 114 -4391 210 -4357
<< viali >>
rect -34 4255 34 4289
rect -96 3220 -62 4196
rect 62 3220 96 4196
rect -34 3127 34 3161
rect -34 3019 34 3053
rect -96 1984 -62 2960
rect 62 1984 96 2960
rect -34 1891 34 1925
rect -34 1783 34 1817
rect -96 748 -62 1724
rect 62 748 96 1724
rect -34 655 34 689
rect -34 547 34 581
rect -96 -488 -62 488
rect 62 -488 96 488
rect -34 -581 34 -547
rect -34 -689 34 -655
rect -96 -1724 -62 -748
rect 62 -1724 96 -748
rect -34 -1817 34 -1783
rect -34 -1925 34 -1891
rect -96 -2960 -62 -1984
rect 62 -2960 96 -1984
rect -34 -3053 34 -3019
rect -34 -3161 34 -3127
rect -96 -4196 -62 -3220
rect 62 -4196 96 -3220
rect -34 -4289 34 -4255
<< metal1 >>
rect -46 4289 46 4295
rect -46 4255 -34 4289
rect 34 4255 46 4289
rect -46 4249 46 4255
rect -102 4196 -56 4208
rect -102 3220 -96 4196
rect -62 3220 -56 4196
rect -102 3208 -56 3220
rect 56 4196 102 4208
rect 56 3220 62 4196
rect 96 3220 102 4196
rect 56 3208 102 3220
rect -46 3161 46 3167
rect -46 3127 -34 3161
rect 34 3127 46 3161
rect -46 3121 46 3127
rect -46 3053 46 3059
rect -46 3019 -34 3053
rect 34 3019 46 3053
rect -46 3013 46 3019
rect -102 2960 -56 2972
rect -102 1984 -96 2960
rect -62 1984 -56 2960
rect -102 1972 -56 1984
rect 56 2960 102 2972
rect 56 1984 62 2960
rect 96 1984 102 2960
rect 56 1972 102 1984
rect -46 1925 46 1931
rect -46 1891 -34 1925
rect 34 1891 46 1925
rect -46 1885 46 1891
rect -46 1817 46 1823
rect -46 1783 -34 1817
rect 34 1783 46 1817
rect -46 1777 46 1783
rect -102 1724 -56 1736
rect -102 748 -96 1724
rect -62 748 -56 1724
rect -102 736 -56 748
rect 56 1724 102 1736
rect 56 748 62 1724
rect 96 748 102 1724
rect 56 736 102 748
rect -46 689 46 695
rect -46 655 -34 689
rect 34 655 46 689
rect -46 649 46 655
rect -46 581 46 587
rect -46 547 -34 581
rect 34 547 46 581
rect -46 541 46 547
rect -102 488 -56 500
rect -102 -488 -96 488
rect -62 -488 -56 488
rect -102 -500 -56 -488
rect 56 488 102 500
rect 56 -488 62 488
rect 96 -488 102 488
rect 56 -500 102 -488
rect -46 -547 46 -541
rect -46 -581 -34 -547
rect 34 -581 46 -547
rect -46 -587 46 -581
rect -46 -655 46 -649
rect -46 -689 -34 -655
rect 34 -689 46 -655
rect -46 -695 46 -689
rect -102 -748 -56 -736
rect -102 -1724 -96 -748
rect -62 -1724 -56 -748
rect -102 -1736 -56 -1724
rect 56 -748 102 -736
rect 56 -1724 62 -748
rect 96 -1724 102 -748
rect 56 -1736 102 -1724
rect -46 -1783 46 -1777
rect -46 -1817 -34 -1783
rect 34 -1817 46 -1783
rect -46 -1823 46 -1817
rect -46 -1891 46 -1885
rect -46 -1925 -34 -1891
rect 34 -1925 46 -1891
rect -46 -1931 46 -1925
rect -102 -1984 -56 -1972
rect -102 -2960 -96 -1984
rect -62 -2960 -56 -1984
rect -102 -2972 -56 -2960
rect 56 -1984 102 -1972
rect 56 -2960 62 -1984
rect 96 -2960 102 -1984
rect 56 -2972 102 -2960
rect -46 -3019 46 -3013
rect -46 -3053 -34 -3019
rect 34 -3053 46 -3019
rect -46 -3059 46 -3053
rect -46 -3127 46 -3121
rect -46 -3161 -34 -3127
rect 34 -3161 46 -3127
rect -46 -3167 46 -3161
rect -102 -3220 -56 -3208
rect -102 -4196 -96 -3220
rect -62 -4196 -56 -3220
rect -102 -4208 -56 -4196
rect 56 -3220 102 -3208
rect 56 -4196 62 -3220
rect 96 -4196 102 -3220
rect 56 -4208 102 -4196
rect -46 -4255 46 -4249
rect -46 -4289 -34 -4255
rect 34 -4289 46 -4255
rect -46 -4295 46 -4289
<< properties >>
string FIXED_BBOX -193 -4374 193 4374
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l .5 m 7 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
