magic
tech sky130A
magscale 1 2
timestamp 1682004071
<< xpolycontact >>
rect -573 6900 573 7332
rect -573 -7332 573 -6900
<< ppolyres >>
rect -573 -6900 573 6900
<< viali >>
rect -557 6917 557 7314
rect -557 -7314 557 -6917
<< metal1 >>
rect -569 7314 569 7320
rect -569 6917 -557 7314
rect 557 6917 569 7314
rect -569 6911 569 6917
rect -569 -6917 569 -6911
rect -569 -7314 -557 -6917
rect 557 -7314 569 -6917
rect -569 -7320 569 -7314
<< res5p73 >>
rect -575 -6902 575 6902
<< properties >>
string gencell sky130_fd_pr__res_high_po_5p73
string library sky130
string parameters w 5.730 l 69 m 1 nx 1 wmin 5.730 lmin 0.50 rho 319.8 val 3.918k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 5.730 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
