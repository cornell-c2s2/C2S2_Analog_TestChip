magic
tech sky130A
magscale 1 2
timestamp 1683899510
<< metal4 >>
rect -200 200 200 257
rect -200 -257 200 -200
<< rmetal4 >>
rect -200 -200 200 200
<< properties >>
string gencell sky130_fd_pr__res_generic_m4
string library sky130
string parameters w 2 l 2 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 47.0m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
