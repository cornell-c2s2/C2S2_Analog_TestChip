magic
tech sky130A
magscale 1 2
timestamp 1679153697
<< error_p >>
rect -1750 3550 1749 3690
rect -1750 3310 1749 3450
rect -1750 50 1749 190
rect -1750 -190 1749 -50
rect -1750 -3450 1749 -3310
rect -1750 -3690 1749 -3550
<< metal3 >>
rect -1750 6922 1749 6950
rect -1750 3578 1665 6922
rect 1729 3578 1749 6922
rect -1750 3550 1749 3578
rect -1750 3422 1749 3450
rect -1750 78 1665 3422
rect 1729 78 1749 3422
rect -1750 50 1749 78
rect -1750 -78 1749 -50
rect -1750 -3422 1665 -78
rect 1729 -3422 1749 -78
rect -1750 -3450 1749 -3422
rect -1750 -3578 1749 -3550
rect -1750 -6922 1665 -3578
rect 1729 -6922 1749 -3578
rect -1750 -6950 1749 -6922
<< via3 >>
rect 1665 3578 1729 6922
rect 1665 78 1729 3422
rect 1665 -3422 1729 -78
rect 1665 -6922 1729 -3578
<< mimcap >>
rect -1650 6810 1550 6850
rect -1650 3690 -1610 6810
rect 1510 3690 1550 6810
rect -1650 3650 1550 3690
rect -1650 3310 1550 3350
rect -1650 190 -1610 3310
rect 1510 190 1550 3310
rect -1650 150 1550 190
rect -1650 -190 1550 -150
rect -1650 -3310 -1610 -190
rect 1510 -3310 1550 -190
rect -1650 -3350 1550 -3310
rect -1650 -3690 1550 -3650
rect -1650 -6810 -1610 -3690
rect 1510 -6810 1550 -3690
rect -1650 -6850 1550 -6810
<< mimcapcontact >>
rect -1610 3690 1510 6810
rect -1610 190 1510 3310
rect -1610 -3310 1510 -190
rect -1610 -6810 1510 -3690
<< metal4 >>
rect -102 6811 2 7000
rect 1618 6938 1722 7000
rect 1618 6922 1745 6938
rect -1611 6810 1511 6811
rect -1611 3690 -1610 6810
rect 1510 3690 1511 6810
rect -1611 3689 1511 3690
rect -102 3311 2 3689
rect 1618 3578 1665 6922
rect 1729 3578 1745 6922
rect 1618 3562 1745 3578
rect 1618 3438 1722 3562
rect 1618 3422 1745 3438
rect -1611 3310 1511 3311
rect -1611 190 -1610 3310
rect 1510 190 1511 3310
rect -1611 189 1511 190
rect -102 -189 2 189
rect 1618 78 1665 3422
rect 1729 78 1745 3422
rect 1618 62 1745 78
rect 1618 -62 1722 62
rect 1618 -78 1745 -62
rect -1611 -190 1511 -189
rect -1611 -3310 -1610 -190
rect 1510 -3310 1511 -190
rect -1611 -3311 1511 -3310
rect -102 -3689 2 -3311
rect 1618 -3422 1665 -78
rect 1729 -3422 1745 -78
rect 1618 -3438 1745 -3422
rect 1618 -3562 1722 -3438
rect 1618 -3578 1745 -3562
rect -1611 -3690 1511 -3689
rect -1611 -6810 -1610 -3690
rect 1510 -6810 1511 -3690
rect -1611 -6811 1511 -6810
rect -102 -7000 2 -6811
rect 1618 -6922 1665 -3578
rect 1729 -6922 1745 -3578
rect 1618 -6938 1745 -6922
rect 1618 -7000 1722 -6938
<< properties >>
string FIXED_BBOX -1750 3550 1650 6950
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 16 l 16 val 524.159 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
