magic
tech sky130A
magscale 1 2
timestamp 1683391037
<< nwell >>
rect -1410 6040 5250 10790
<< pwell >>
rect 7180 8770 7840 8780
<< locali >>
rect -4070 10060 -3410 10180
rect 7180 10060 7840 10180
<< viali >>
rect -4040 8650 -3860 8750
rect -3620 8650 -3440 8750
rect 7210 8650 7390 8750
rect 7630 8650 7810 8750
rect 900 7430 1470 7670
rect 2370 7430 2940 7670
<< metal1 >>
rect -5050 10230 -4610 11420
rect -5940 10210 -4610 10230
rect -5940 10140 -5810 10210
rect -5740 10140 -4610 10210
rect -5940 10100 -4610 10140
rect -5940 10030 -5920 10100
rect -5850 10030 -4610 10100
rect -5940 10010 -4610 10030
rect -5050 8810 -4610 10010
rect -2620 10150 -2180 11430
rect 1240 10930 2620 10980
rect 1240 10660 1270 10930
rect 1540 10660 2320 10930
rect 2590 10660 2620 10930
rect 1240 10640 2620 10660
rect -1410 10530 5250 10580
rect -1410 10150 -1330 10530
rect -1290 10380 -1280 10450
rect -1210 10380 -1200 10450
rect -970 10380 -960 10450
rect -890 10380 -880 10450
rect -660 10380 -650 10450
rect -580 10380 -570 10450
rect -340 10380 -330 10450
rect -260 10380 -250 10450
rect -30 10380 -20 10450
rect 50 10380 60 10450
rect 290 10380 300 10450
rect 370 10380 380 10450
rect 610 10380 620 10450
rect 690 10380 700 10450
rect 920 10380 930 10450
rect 1000 10380 1010 10450
rect 1240 10380 1250 10450
rect 1320 10380 1330 10450
rect 1560 10380 1570 10450
rect 1640 10380 1650 10450
rect 1870 10380 1880 10450
rect 1950 10380 1960 10450
rect 2190 10380 2200 10450
rect 2270 10380 2280 10450
rect 2500 10380 2510 10450
rect 2580 10380 2590 10450
rect 2820 10380 2830 10450
rect 2900 10380 2910 10450
rect 3140 10380 3150 10450
rect 3220 10380 3230 10450
rect 3450 10380 3460 10450
rect 3530 10380 3540 10450
rect 3770 10380 3780 10450
rect 3850 10380 3860 10450
rect 4080 10380 4090 10450
rect 4160 10380 4170 10450
rect 4400 10380 4410 10450
rect 4480 10380 4490 10450
rect 4720 10380 4730 10450
rect 4800 10380 4810 10450
rect 5030 10380 5040 10450
rect 5110 10380 5120 10450
rect -2620 9860 -1330 10150
rect -1290 10140 -1280 10210
rect -1210 10140 -1200 10210
rect -970 10140 -960 10210
rect -890 10140 -880 10210
rect -660 10140 -650 10210
rect -580 10140 -570 10210
rect -340 10140 -330 10210
rect -260 10140 -250 10210
rect -30 10140 -20 10210
rect 50 10140 60 10210
rect 290 10140 300 10210
rect 370 10140 380 10210
rect 610 10140 620 10210
rect 690 10140 700 10210
rect 920 10140 930 10210
rect 1000 10140 1010 10210
rect 1240 10140 1250 10210
rect 1320 10140 1330 10210
rect 1560 10140 1570 10210
rect 1640 10140 1650 10210
rect 1870 10140 1880 10210
rect 1950 10140 1960 10210
rect 2190 10140 2200 10210
rect 2270 10140 2280 10210
rect 2500 10140 2510 10210
rect 2580 10140 2590 10210
rect 2820 10140 2830 10210
rect 2900 10140 2910 10210
rect 3140 10140 3150 10210
rect 3220 10140 3230 10210
rect 3450 10140 3460 10210
rect 3530 10140 3540 10210
rect 3770 10140 3780 10210
rect 3850 10140 3860 10210
rect 4080 10140 4090 10210
rect 4160 10140 4170 10210
rect 4400 10140 4410 10210
rect 4480 10140 4490 10210
rect 4720 10140 4730 10210
rect 4800 10140 4810 10210
rect 5030 10140 5040 10210
rect 5110 10140 5120 10210
rect 5170 10150 5250 10530
rect 6020 10150 6450 11420
rect -2620 8810 -2180 9860
rect -1410 9450 -1330 9860
rect 5170 9860 6450 10150
rect -1130 9770 -1120 9840
rect -1050 9770 -1040 9840
rect -820 9770 -810 9840
rect -740 9770 -730 9840
rect -500 9770 -490 9840
rect -420 9770 -410 9840
rect -180 9770 -170 9840
rect -100 9770 -90 9840
rect 130 9770 140 9840
rect 210 9770 220 9840
rect 450 9770 460 9840
rect 530 9770 540 9840
rect 760 9770 770 9840
rect 840 9770 850 9840
rect 1080 9770 1090 9840
rect 1160 9770 1170 9840
rect 1400 9770 1410 9840
rect 1480 9770 1490 9840
rect 1710 9770 1720 9840
rect 1790 9770 1800 9840
rect 2030 9770 2040 9840
rect 2110 9770 2120 9840
rect 2350 9770 2360 9840
rect 2430 9770 2440 9840
rect 2660 9770 2670 9840
rect 2740 9770 2750 9840
rect 2980 9770 2990 9840
rect 3060 9770 3070 9840
rect 3290 9770 3300 9840
rect 3370 9770 3380 9840
rect 3610 9770 3620 9840
rect 3690 9770 3700 9840
rect 3930 9770 3940 9840
rect 4010 9770 4020 9840
rect 4240 9770 4250 9840
rect 4320 9770 4330 9840
rect 4560 9770 4570 9840
rect 4640 9770 4650 9840
rect 4880 9770 4890 9840
rect 4960 9770 4970 9840
rect -1130 9530 -1120 9600
rect -1050 9530 -1040 9600
rect -820 9530 -810 9600
rect -740 9530 -730 9600
rect -500 9530 -490 9600
rect -420 9530 -410 9600
rect -180 9530 -170 9600
rect -100 9530 -90 9600
rect 130 9530 140 9600
rect 210 9530 220 9600
rect 450 9530 460 9600
rect 530 9530 540 9600
rect 760 9530 770 9600
rect 840 9530 850 9600
rect 1080 9530 1090 9600
rect 1160 9530 1170 9600
rect 1400 9530 1410 9600
rect 1480 9530 1490 9600
rect 1710 9530 1720 9600
rect 1790 9530 1800 9600
rect 2030 9530 2040 9600
rect 2110 9530 2120 9600
rect 2350 9530 2360 9600
rect 2430 9530 2440 9600
rect 2660 9530 2670 9600
rect 2740 9530 2750 9600
rect 2980 9530 2990 9600
rect 3060 9530 3070 9600
rect 3290 9530 3300 9600
rect 3370 9530 3380 9600
rect 3610 9530 3620 9600
rect 3690 9530 3700 9600
rect 3930 9530 3940 9600
rect 4010 9530 4020 9600
rect 4240 9530 4250 9600
rect 4320 9530 4330 9600
rect 4560 9530 4570 9600
rect 4640 9530 4650 9600
rect 4880 9530 4890 9600
rect 4960 9530 4970 9600
rect 5170 9450 5250 9860
rect -1410 9430 5250 9450
rect -1410 9400 -160 9430
rect -200 9350 -160 9400
rect -80 9400 3900 9430
rect -80 9350 -40 9400
rect 3860 9350 3900 9400
rect 3980 9400 5250 9430
rect 3980 9350 4020 9400
rect -200 9340 -40 9350
rect 1020 9290 2810 9350
rect 3860 9340 4020 9350
rect 1020 9020 1270 9290
rect 1540 9020 2320 9290
rect 2590 9020 2810 9290
rect 1020 8960 2810 9020
rect 90 8860 3740 8910
rect -4052 8750 -3848 8756
rect -4052 8650 -4040 8750
rect -3860 8650 -3848 8750
rect -4052 8644 -3848 8650
rect -3632 8750 -3428 8756
rect -3632 8650 -3620 8750
rect -3440 8650 -3428 8750
rect -3632 8644 -3428 8650
rect 90 7780 170 8860
rect 210 8710 220 8780
rect 290 8710 300 8780
rect 530 8710 540 8780
rect 610 8710 620 8780
rect 840 8710 850 8780
rect 920 8710 930 8780
rect 1160 8710 1170 8780
rect 1240 8710 1250 8780
rect 1480 8710 1490 8780
rect 1560 8710 1570 8780
rect 1790 8710 1800 8780
rect 1870 8710 1880 8780
rect 2110 8710 2120 8780
rect 2190 8710 2200 8780
rect 2430 8710 2440 8780
rect 2510 8710 2520 8780
rect 2740 8710 2750 8780
rect 2820 8710 2830 8780
rect 3060 8710 3070 8780
rect 3140 8710 3150 8780
rect 3370 8710 3380 8780
rect 3450 8710 3460 8780
rect 210 8500 220 8570
rect 290 8500 300 8570
rect 530 8500 540 8570
rect 610 8500 620 8570
rect 840 8500 850 8570
rect 920 8500 930 8570
rect 1160 8500 1170 8570
rect 1240 8500 1250 8570
rect 1480 8500 1490 8570
rect 1560 8500 1570 8570
rect 1790 8500 1800 8570
rect 1870 8500 1880 8570
rect 2110 8500 2120 8570
rect 2190 8500 2200 8570
rect 2430 8500 2440 8570
rect 2510 8500 2520 8570
rect 2740 8500 2750 8570
rect 2820 8500 2830 8570
rect 3060 8500 3070 8570
rect 3140 8500 3150 8570
rect 3370 8500 3380 8570
rect 3450 8500 3460 8570
rect 370 8070 380 8140
rect 450 8070 460 8140
rect 690 8070 700 8140
rect 770 8070 780 8140
rect 1000 8070 1010 8140
rect 1080 8070 1090 8140
rect 1320 8070 1330 8140
rect 1400 8070 1410 8140
rect 1640 8070 1650 8140
rect 1720 8070 1730 8140
rect 1950 8070 1960 8140
rect 2030 8070 2040 8140
rect 2270 8070 2280 8140
rect 2350 8070 2360 8140
rect 2580 8070 2590 8140
rect 2660 8070 2670 8140
rect 2900 8070 2910 8140
rect 2980 8070 2990 8140
rect 3220 8070 3230 8140
rect 3300 8070 3310 8140
rect 3530 8070 3540 8140
rect 3610 8070 3620 8140
rect 370 7860 380 7930
rect 450 7860 460 7930
rect 690 7860 700 7930
rect 770 7860 780 7930
rect 1000 7860 1010 7930
rect 1080 7860 1090 7930
rect 1320 7860 1330 7930
rect 1400 7860 1410 7930
rect 1640 7860 1650 7930
rect 1720 7860 1730 7930
rect 1950 7860 1960 7930
rect 2030 7860 2040 7930
rect 2270 7860 2280 7930
rect 2350 7860 2360 7930
rect 2580 7860 2590 7930
rect 2660 7860 2670 7930
rect 2900 7860 2910 7930
rect 2980 7860 2990 7930
rect 3220 7860 3230 7930
rect 3300 7860 3310 7930
rect 3530 7860 3540 7930
rect 3610 7860 3620 7930
rect 3660 7780 3740 8860
rect 6020 8810 6450 9860
rect 8450 10230 8890 11420
rect 8450 10210 9780 10230
rect 8450 10140 9580 10210
rect 9650 10140 9780 10210
rect 8450 10100 9780 10140
rect 8450 10030 9690 10100
rect 9760 10030 9780 10100
rect 8450 10010 9780 10030
rect 8450 8810 8890 10010
rect 7198 8750 7402 8756
rect 7198 8650 7210 8750
rect 7390 8650 7402 8750
rect 7198 8644 7402 8650
rect 7618 8750 7822 8756
rect 7618 8650 7630 8750
rect 7810 8650 7822 8750
rect 7618 8644 7822 8650
rect 90 7730 3740 7780
rect 280 7370 550 7730
rect 1030 7676 1040 7680
rect 888 7670 1040 7676
rect 1300 7676 1310 7680
rect 1300 7670 1482 7676
rect 888 7430 900 7670
rect 1470 7430 1482 7670
rect 888 7424 1040 7430
rect 1030 7420 1040 7424
rect 1300 7424 1482 7430
rect 1300 7420 1310 7424
rect 1780 7370 2050 7730
rect 2530 7676 2540 7680
rect 2358 7670 2540 7676
rect 2800 7676 2810 7680
rect 2800 7670 2952 7676
rect 2358 7430 2370 7670
rect 2940 7430 2952 7670
rect 2358 7424 2540 7430
rect 2530 7420 2540 7424
rect 2800 7424 2952 7430
rect 2800 7420 2810 7424
rect 3280 7370 3550 7730
rect 280 7320 3550 7370
rect 210 7160 220 7230
rect 290 7160 300 7230
rect 530 7160 540 7230
rect 610 7160 620 7230
rect 210 6950 220 7020
rect 290 6950 300 7020
rect 530 6950 540 7020
rect 610 6950 620 7020
rect 700 6600 760 7320
rect 840 7160 850 7230
rect 920 7160 930 7230
rect 840 6950 850 7020
rect 920 6950 930 7020
rect 1020 6600 1080 7320
rect 1160 7160 1170 7230
rect 1240 7160 1250 7230
rect 1480 7160 1490 7230
rect 1560 7160 1570 7230
rect 1790 7160 1800 7230
rect 1870 7160 1880 7230
rect 2110 7160 2120 7230
rect 2190 7160 2200 7230
rect 2420 7160 2430 7230
rect 2500 7160 2510 7230
rect 2740 7160 2750 7230
rect 2820 7160 2830 7230
rect 1160 6950 1170 7020
rect 1240 6950 1250 7020
rect 1480 6950 1490 7020
rect 1560 6950 1570 7020
rect 1790 6950 1800 7020
rect 1870 6950 1880 7020
rect 2110 6950 2120 7020
rect 2190 6950 2200 7020
rect 2420 6950 2430 7020
rect 2500 6950 2510 7020
rect 2740 6950 2750 7020
rect 2820 6950 2830 7020
rect 2910 6600 2970 7320
rect 3060 7160 3070 7230
rect 3140 7160 3150 7230
rect 3060 6950 3070 7020
rect 3140 6950 3150 7020
rect 3230 6600 3290 7320
rect 3370 7160 3380 7230
rect 3450 7160 3460 7230
rect 3370 6950 3380 7020
rect 3450 6950 3460 7020
rect 370 6530 380 6600
rect 450 6530 460 6600
rect 690 6530 700 6600
rect 770 6530 780 6600
rect 1000 6530 1010 6600
rect 1080 6530 1090 6600
rect 1320 6530 1330 6600
rect 1400 6530 1410 6600
rect 1630 6530 1640 6600
rect 1710 6530 1720 6600
rect 1950 6530 1960 6600
rect 2030 6530 2040 6600
rect 2270 6530 2280 6600
rect 2350 6530 2360 6600
rect 2580 6530 2590 6600
rect 2660 6530 2670 6600
rect 2900 6530 2910 6600
rect 2980 6530 2990 6600
rect 3210 6530 3220 6600
rect 3290 6530 3300 6600
rect 3530 6530 3540 6600
rect 3610 6530 3620 6600
rect 700 6390 760 6530
rect 1020 6390 1080 6530
rect 2910 6390 2970 6530
rect 3230 6390 3290 6530
rect 370 6320 380 6390
rect 450 6320 460 6390
rect 690 6320 700 6390
rect 770 6320 780 6390
rect 1000 6320 1010 6390
rect 1080 6320 1090 6390
rect 1320 6320 1330 6390
rect 1400 6320 1410 6390
rect 1630 6320 1640 6390
rect 1710 6320 1720 6390
rect 1950 6320 1960 6390
rect 2030 6320 2040 6390
rect 2270 6320 2280 6390
rect 2350 6320 2360 6390
rect 2580 6320 2590 6390
rect 2660 6320 2670 6390
rect 2900 6320 2910 6390
rect 2980 6320 2990 6390
rect 3210 6320 3220 6390
rect 3290 6320 3300 6390
rect 3530 6320 3540 6390
rect 3610 6320 3620 6390
rect 700 6240 760 6320
rect 1020 6240 1080 6320
rect 2910 6240 2970 6320
rect 3230 6240 3290 6320
rect 280 6190 3550 6240
rect 1130 5740 2690 5790
rect 1130 4680 1210 5740
rect 1310 5600 1320 5670
rect 1390 5600 1400 5670
rect 1630 5600 1640 5670
rect 1710 5600 1720 5670
rect 1940 5600 1950 5670
rect 2020 5600 2030 5670
rect 2260 5600 2270 5670
rect 2340 5600 2350 5670
rect 1310 5310 1320 5380
rect 1390 5310 1400 5380
rect 1630 5310 1640 5380
rect 1710 5310 1720 5380
rect 1940 5310 1950 5380
rect 2020 5310 2030 5380
rect 2260 5310 2270 5380
rect 2340 5310 2350 5380
rect 1470 5040 1480 5110
rect 1550 5040 1560 5110
rect 1780 5040 1790 5110
rect 1860 5040 1870 5110
rect 2100 5040 2110 5110
rect 2180 5040 2190 5110
rect 2420 5040 2430 5110
rect 2500 5040 2510 5110
rect 1470 4750 1480 4820
rect 1550 4750 1560 4820
rect 1780 4750 1790 4820
rect 1860 4750 1870 4820
rect 2100 4750 2110 4820
rect 2180 4750 2190 4820
rect 2420 4750 2430 4820
rect 2500 4750 2510 4820
rect 2610 4680 2690 5740
rect 1130 4630 2690 4680
rect 1770 4320 1780 4580
rect 2040 4320 2050 4580
rect 1130 4220 2690 4270
rect 1130 3160 1210 4220
rect 1310 4080 1320 4150
rect 1390 4080 1400 4150
rect 1630 4080 1640 4150
rect 1710 4080 1720 4150
rect 1940 4080 1950 4150
rect 2020 4080 2030 4150
rect 2260 4080 2270 4150
rect 2340 4080 2350 4150
rect 1310 3790 1320 3860
rect 1390 3790 1400 3860
rect 1630 3790 1640 3860
rect 1710 3790 1720 3860
rect 1940 3790 1950 3860
rect 2020 3790 2030 3860
rect 2260 3790 2270 3860
rect 2340 3790 2350 3860
rect 1470 3520 1480 3590
rect 1550 3520 1560 3590
rect 1780 3520 1790 3590
rect 1860 3520 1870 3590
rect 2100 3520 2110 3590
rect 2180 3520 2190 3590
rect 2420 3520 2430 3590
rect 2500 3520 2510 3590
rect 1470 3230 1480 3300
rect 1550 3230 1560 3300
rect 1780 3230 1790 3300
rect 1860 3230 1870 3300
rect 2100 3230 2110 3300
rect 2180 3230 2190 3300
rect 2420 3230 2430 3300
rect 2500 3230 2510 3300
rect 2610 3160 2690 4220
rect 1130 3110 2690 3160
rect 1770 2800 1780 3060
rect 2040 2800 2050 3060
rect -490 2750 -480 2780
rect -500 2700 -480 2750
rect -490 2670 -480 2700
rect -370 2750 -360 2780
rect -240 2750 -230 2780
rect -370 2700 -230 2750
rect -370 2670 -360 2700
rect -240 2670 -230 2700
rect -120 2750 -110 2780
rect 3910 2750 3920 2780
rect -120 2700 3920 2750
rect -120 2670 -110 2700
rect 3910 2670 3920 2700
rect 4030 2750 4040 2780
rect 4160 2750 4170 2780
rect 4030 2700 4170 2750
rect 4030 2670 4040 2700
rect 4160 2670 4170 2700
rect 4280 2750 4290 2780
rect 4280 2700 4300 2750
rect 4280 2670 4290 2700
rect 320 2560 330 2630
rect 400 2560 410 2630
rect 840 2560 850 2630
rect 920 2560 930 2630
rect 1350 2560 1360 2630
rect 1430 2560 1440 2630
rect 1870 2560 1880 2630
rect 1950 2560 1960 2630
rect 2380 2560 2390 2630
rect 2460 2560 2470 2630
rect 2900 2560 2910 2630
rect 2980 2560 2990 2630
rect 3420 2560 3430 2630
rect 3500 2560 3510 2630
rect 320 2380 330 2450
rect 400 2380 410 2450
rect 840 2380 850 2450
rect 920 2380 930 2450
rect 1350 2380 1360 2450
rect 1430 2380 1440 2450
rect 1870 2380 1880 2450
rect 1950 2380 1960 2450
rect 2380 2380 2390 2450
rect 2460 2380 2470 2450
rect 2900 2380 2910 2450
rect 2980 2380 2990 2450
rect 3420 2380 3430 2450
rect 3500 2380 3510 2450
rect 580 1890 590 1960
rect 660 1890 670 1960
rect 1090 1890 1100 1960
rect 1170 1890 1180 1960
rect 1610 1890 1620 1960
rect 1690 1890 1700 1960
rect 2130 1890 2140 1960
rect 2210 1890 2220 1960
rect 2640 1890 2650 1960
rect 2720 1890 2730 1960
rect 3160 1890 3170 1960
rect 3240 1890 3250 1960
rect 580 1710 590 1780
rect 660 1710 670 1780
rect 1090 1710 1100 1780
rect 1170 1710 1180 1780
rect 1610 1710 1620 1780
rect 1690 1710 1700 1780
rect 2130 1710 2140 1780
rect 2210 1710 2220 1780
rect 2640 1710 2650 1780
rect 2720 1710 2730 1780
rect 3160 1710 3170 1780
rect 3240 1710 3250 1780
rect -490 1640 -480 1670
rect -500 1590 -480 1640
rect -490 1560 -480 1590
rect -370 1640 -360 1670
rect -240 1640 -230 1670
rect -370 1590 -230 1640
rect -370 1560 -360 1590
rect -240 1560 -230 1590
rect -120 1640 -110 1670
rect 3910 1640 3920 1670
rect -120 1590 3920 1640
rect -120 1560 -110 1590
rect 3910 1560 3920 1590
rect 4030 1640 4040 1670
rect 4160 1640 4170 1670
rect 4030 1590 4170 1640
rect 4030 1560 4040 1590
rect 4160 1560 4170 1590
rect 4280 1640 4290 1670
rect 4280 1590 4300 1640
rect 4280 1560 4290 1590
rect 1780 1290 1790 1540
rect 2040 1290 2050 1540
rect 1780 1280 2050 1290
rect -490 1230 -480 1260
rect -500 1180 -480 1230
rect -490 1150 -480 1180
rect -370 1230 -360 1260
rect -240 1230 -230 1260
rect -370 1180 -230 1230
rect -370 1150 -360 1180
rect -240 1150 -230 1180
rect -120 1230 -110 1260
rect 3910 1230 3920 1260
rect -120 1180 3920 1230
rect -120 1150 -110 1180
rect 3910 1150 3920 1180
rect 4030 1230 4040 1260
rect 4160 1230 4170 1260
rect 4030 1180 4170 1230
rect 4030 1150 4040 1180
rect 4160 1150 4170 1180
rect 4280 1230 4290 1260
rect 4280 1180 4300 1230
rect 4280 1150 4290 1180
rect 60 1040 70 1110
rect 140 1040 150 1110
rect 580 1040 590 1110
rect 660 1040 670 1110
rect 1090 1040 1100 1110
rect 1170 1040 1180 1110
rect 1610 1040 1620 1110
rect 1690 1040 1700 1110
rect 2120 1040 2130 1110
rect 2200 1040 2210 1110
rect 2640 1040 2650 1110
rect 2720 1040 2730 1110
rect 3160 1040 3170 1110
rect 3240 1040 3250 1110
rect 3670 1040 3680 1110
rect 3750 1040 3760 1110
rect 60 860 70 930
rect 140 860 150 930
rect 580 860 590 930
rect 660 860 670 930
rect 1090 860 1100 930
rect 1170 860 1180 930
rect 1610 860 1620 930
rect 1690 860 1700 930
rect 2120 860 2130 930
rect 2200 860 2210 930
rect 2640 860 2650 930
rect 2720 860 2730 930
rect 3160 860 3170 930
rect 3240 860 3250 930
rect 3670 860 3680 930
rect 3750 860 3760 930
rect 320 370 330 440
rect 400 370 410 440
rect 830 370 840 440
rect 910 370 920 440
rect 1350 370 1360 440
rect 1430 370 1440 440
rect 1870 370 1880 440
rect 1950 370 1960 440
rect 2380 370 2390 440
rect 2460 370 2470 440
rect 2900 370 2910 440
rect 2980 370 2990 440
rect 3410 370 3420 440
rect 3490 370 3500 440
rect 320 190 330 260
rect 400 190 410 260
rect 830 190 840 260
rect 910 190 920 260
rect 1350 190 1360 260
rect 1430 190 1440 260
rect 1870 190 1880 260
rect 1950 190 1960 260
rect 2380 190 2390 260
rect 2460 190 2470 260
rect 2900 190 2910 260
rect 2980 190 2990 260
rect 3410 190 3420 260
rect 3490 190 3500 260
rect -490 120 -480 150
rect -500 70 -480 120
rect -490 40 -480 70
rect -370 120 -360 150
rect -240 120 -230 150
rect -370 70 -230 120
rect -370 40 -360 70
rect -240 40 -230 70
rect -120 120 -110 150
rect 3910 120 3920 150
rect -120 70 3920 120
rect -120 40 -110 70
rect 3910 40 3920 70
rect 4030 120 4040 150
rect 4160 120 4170 150
rect 4030 70 4170 120
rect 4030 40 4040 70
rect 4160 40 4170 70
rect 4280 120 4290 150
rect 4280 70 4300 120
rect 4280 40 4290 70
rect 1780 -240 1790 10
rect 2040 -240 2050 10
<< via1 >>
rect -5810 10140 -5740 10210
rect -5920 10030 -5850 10100
rect 1270 10660 1540 10930
rect 2320 10660 2590 10930
rect -1280 10380 -1210 10450
rect -960 10380 -890 10450
rect -650 10380 -580 10450
rect -330 10380 -260 10450
rect -20 10380 50 10450
rect 300 10380 370 10450
rect 620 10380 690 10450
rect 930 10380 1000 10450
rect 1250 10380 1320 10450
rect 1570 10380 1640 10450
rect 1880 10380 1950 10450
rect 2200 10380 2270 10450
rect 2510 10380 2580 10450
rect 2830 10380 2900 10450
rect 3150 10380 3220 10450
rect 3460 10380 3530 10450
rect 3780 10380 3850 10450
rect 4090 10380 4160 10450
rect 4410 10380 4480 10450
rect 4730 10380 4800 10450
rect 5040 10380 5110 10450
rect -1280 10140 -1210 10210
rect -960 10140 -890 10210
rect -650 10140 -580 10210
rect -330 10140 -260 10210
rect -20 10140 50 10210
rect 300 10140 370 10210
rect 620 10140 690 10210
rect 930 10140 1000 10210
rect 1250 10140 1320 10210
rect 1570 10140 1640 10210
rect 1880 10140 1950 10210
rect 2200 10140 2270 10210
rect 2510 10140 2580 10210
rect 2830 10140 2900 10210
rect 3150 10140 3220 10210
rect 3460 10140 3530 10210
rect 3780 10140 3850 10210
rect 4090 10140 4160 10210
rect 4410 10140 4480 10210
rect 4730 10140 4800 10210
rect 5040 10140 5110 10210
rect -1120 9770 -1050 9840
rect -810 9770 -740 9840
rect -490 9770 -420 9840
rect -170 9770 -100 9840
rect 140 9770 210 9840
rect 460 9770 530 9840
rect 770 9770 840 9840
rect 1090 9770 1160 9840
rect 1410 9770 1480 9840
rect 1720 9770 1790 9840
rect 2040 9770 2110 9840
rect 2360 9770 2430 9840
rect 2670 9770 2740 9840
rect 2990 9770 3060 9840
rect 3300 9770 3370 9840
rect 3620 9770 3690 9840
rect 3940 9770 4010 9840
rect 4250 9770 4320 9840
rect 4570 9770 4640 9840
rect 4890 9770 4960 9840
rect -1120 9530 -1050 9600
rect -810 9530 -740 9600
rect -490 9530 -420 9600
rect -170 9530 -100 9600
rect 140 9530 210 9600
rect 460 9530 530 9600
rect 770 9530 840 9600
rect 1090 9530 1160 9600
rect 1410 9530 1480 9600
rect 1720 9530 1790 9600
rect 2040 9530 2110 9600
rect 2360 9530 2430 9600
rect 2670 9530 2740 9600
rect 2990 9530 3060 9600
rect 3300 9530 3370 9600
rect 3620 9530 3690 9600
rect 3940 9530 4010 9600
rect 4250 9530 4320 9600
rect 4570 9530 4640 9600
rect 4890 9530 4960 9600
rect -160 9350 -80 9430
rect 3900 9350 3980 9430
rect 1270 9020 1540 9290
rect 2320 9020 2590 9290
rect -4040 8650 -3860 8750
rect -3620 8650 -3440 8750
rect 220 8710 290 8780
rect 540 8710 610 8780
rect 850 8710 920 8780
rect 1170 8710 1240 8780
rect 1490 8710 1560 8780
rect 1800 8710 1870 8780
rect 2120 8710 2190 8780
rect 2440 8710 2510 8780
rect 2750 8710 2820 8780
rect 3070 8710 3140 8780
rect 3380 8710 3450 8780
rect 220 8500 290 8570
rect 540 8500 610 8570
rect 850 8500 920 8570
rect 1170 8500 1240 8570
rect 1490 8500 1560 8570
rect 1800 8500 1870 8570
rect 2120 8500 2190 8570
rect 2440 8500 2510 8570
rect 2750 8500 2820 8570
rect 3070 8500 3140 8570
rect 3380 8500 3450 8570
rect 380 8070 450 8140
rect 700 8070 770 8140
rect 1010 8070 1080 8140
rect 1330 8070 1400 8140
rect 1650 8070 1720 8140
rect 1960 8070 2030 8140
rect 2280 8070 2350 8140
rect 2590 8070 2660 8140
rect 2910 8070 2980 8140
rect 3230 8070 3300 8140
rect 3540 8070 3610 8140
rect 380 7860 450 7930
rect 700 7860 770 7930
rect 1010 7860 1080 7930
rect 1330 7860 1400 7930
rect 1650 7860 1720 7930
rect 1960 7860 2030 7930
rect 2280 7860 2350 7930
rect 2590 7860 2660 7930
rect 2910 7860 2980 7930
rect 3230 7860 3300 7930
rect 3540 7860 3610 7930
rect 9580 10140 9650 10210
rect 9690 10030 9760 10100
rect 7210 8650 7390 8750
rect 7630 8650 7810 8750
rect 1040 7670 1300 7680
rect 1040 7430 1300 7670
rect 1040 7420 1300 7430
rect 2540 7670 2800 7680
rect 2540 7430 2800 7670
rect 2540 7420 2800 7430
rect 220 7160 290 7230
rect 540 7160 610 7230
rect 220 6950 290 7020
rect 540 6950 610 7020
rect 850 7160 920 7230
rect 850 6950 920 7020
rect 1170 7160 1240 7230
rect 1490 7160 1560 7230
rect 1800 7160 1870 7230
rect 2120 7160 2190 7230
rect 2430 7160 2500 7230
rect 2750 7160 2820 7230
rect 1170 6950 1240 7020
rect 1490 6950 1560 7020
rect 1800 6950 1870 7020
rect 2120 6950 2190 7020
rect 2430 6950 2500 7020
rect 2750 6950 2820 7020
rect 3070 7160 3140 7230
rect 3070 6950 3140 7020
rect 3380 7160 3450 7230
rect 3380 6950 3450 7020
rect 380 6530 450 6600
rect 700 6530 770 6600
rect 1010 6530 1080 6600
rect 1330 6530 1400 6600
rect 1640 6530 1710 6600
rect 1960 6530 2030 6600
rect 2280 6530 2350 6600
rect 2590 6530 2660 6600
rect 2910 6530 2980 6600
rect 3220 6530 3290 6600
rect 3540 6530 3610 6600
rect 380 6320 450 6390
rect 700 6320 770 6390
rect 1010 6320 1080 6390
rect 1330 6320 1400 6390
rect 1640 6320 1710 6390
rect 1960 6320 2030 6390
rect 2280 6320 2350 6390
rect 2590 6320 2660 6390
rect 2910 6320 2980 6390
rect 3220 6320 3290 6390
rect 3540 6320 3610 6390
rect 1320 5600 1390 5670
rect 1640 5600 1710 5670
rect 1950 5600 2020 5670
rect 2270 5600 2340 5670
rect 1320 5310 1390 5380
rect 1640 5310 1710 5380
rect 1950 5310 2020 5380
rect 2270 5310 2340 5380
rect 1480 5040 1550 5110
rect 1790 5040 1860 5110
rect 2110 5040 2180 5110
rect 2430 5040 2500 5110
rect 1480 4750 1550 4820
rect 1790 4750 1860 4820
rect 2110 4750 2180 4820
rect 2430 4750 2500 4820
rect 1780 4320 2040 4580
rect 1320 4080 1390 4150
rect 1640 4080 1710 4150
rect 1950 4080 2020 4150
rect 2270 4080 2340 4150
rect 1320 3790 1390 3860
rect 1640 3790 1710 3860
rect 1950 3790 2020 3860
rect 2270 3790 2340 3860
rect 1480 3520 1550 3590
rect 1790 3520 1860 3590
rect 2110 3520 2180 3590
rect 2430 3520 2500 3590
rect 1480 3230 1550 3300
rect 1790 3230 1860 3300
rect 2110 3230 2180 3300
rect 2430 3230 2500 3300
rect 1780 2800 2040 3060
rect -480 2670 -370 2780
rect -230 2670 -120 2780
rect 3920 2670 4030 2780
rect 4170 2670 4280 2780
rect 330 2560 400 2630
rect 850 2560 920 2630
rect 1360 2560 1430 2630
rect 1880 2560 1950 2630
rect 2390 2560 2460 2630
rect 2910 2560 2980 2630
rect 3430 2560 3500 2630
rect 330 2380 400 2450
rect 850 2380 920 2450
rect 1360 2380 1430 2450
rect 1880 2380 1950 2450
rect 2390 2380 2460 2450
rect 2910 2380 2980 2450
rect 3430 2380 3500 2450
rect 590 1890 660 1960
rect 1100 1890 1170 1960
rect 1620 1890 1690 1960
rect 2140 1890 2210 1960
rect 2650 1890 2720 1960
rect 3170 1890 3240 1960
rect 590 1710 660 1780
rect 1100 1710 1170 1780
rect 1620 1710 1690 1780
rect 2140 1710 2210 1780
rect 2650 1710 2720 1780
rect 3170 1710 3240 1780
rect -480 1560 -370 1670
rect -230 1560 -120 1670
rect 3920 1560 4030 1670
rect 4170 1560 4280 1670
rect 1790 1290 2040 1540
rect -480 1150 -370 1260
rect -230 1150 -120 1260
rect 3920 1150 4030 1260
rect 4170 1150 4280 1260
rect 70 1040 140 1110
rect 590 1040 660 1110
rect 1100 1040 1170 1110
rect 1620 1040 1690 1110
rect 2130 1040 2200 1110
rect 2650 1040 2720 1110
rect 3170 1040 3240 1110
rect 3680 1040 3750 1110
rect 70 860 140 930
rect 590 860 660 930
rect 1100 860 1170 930
rect 1620 860 1690 930
rect 2130 860 2200 930
rect 2650 860 2720 930
rect 3170 860 3240 930
rect 3680 860 3750 930
rect 330 370 400 440
rect 840 370 910 440
rect 1360 370 1430 440
rect 1880 370 1950 440
rect 2390 370 2460 440
rect 2910 370 2980 440
rect 3420 370 3490 440
rect 330 190 400 260
rect 840 190 910 260
rect 1360 190 1430 260
rect 1880 190 1950 260
rect 2390 190 2460 260
rect 2910 190 2980 260
rect 3420 190 3490 260
rect -480 40 -370 150
rect -230 40 -120 150
rect 3920 40 4030 150
rect 4170 40 4280 150
rect 1790 -240 2040 10
<< metal2 >>
rect 1270 10930 1540 10940
rect 1270 10650 1540 10660
rect 2320 10930 2590 10940
rect 2320 10650 2590 10660
rect -1280 10450 -1210 10460
rect -1280 10370 -1210 10380
rect -960 10450 -890 10460
rect -960 10370 -890 10380
rect -650 10450 -580 10460
rect -650 10370 -580 10380
rect -330 10450 -260 10460
rect -330 10370 -260 10380
rect -20 10450 50 10460
rect -20 10370 50 10380
rect 300 10450 370 10460
rect 300 10370 370 10380
rect 620 10450 690 10460
rect 620 10370 690 10380
rect 930 10450 1000 10460
rect 930 10370 1000 10380
rect 1250 10450 1320 10460
rect 1250 10370 1320 10380
rect 1570 10450 1640 10460
rect 1570 10370 1640 10380
rect 1880 10450 1950 10460
rect 1880 10370 1950 10380
rect 2200 10450 2270 10460
rect 2200 10370 2270 10380
rect 2510 10450 2580 10460
rect 2510 10370 2580 10380
rect 2830 10450 2900 10460
rect 2830 10370 2900 10380
rect 3150 10450 3220 10460
rect 3150 10370 3220 10380
rect 3460 10450 3530 10460
rect 3460 10370 3530 10380
rect 3780 10450 3850 10460
rect 3780 10370 3850 10380
rect 4090 10450 4160 10460
rect 4090 10370 4160 10380
rect 4410 10450 4480 10460
rect 4410 10370 4480 10380
rect 4730 10450 4800 10460
rect 4730 10370 4800 10380
rect 5040 10450 5110 10460
rect 5040 10370 5110 10380
rect -5940 10210 -5720 10230
rect -5940 10140 -5810 10210
rect -5740 10140 -5720 10210
rect -5940 10100 -5720 10140
rect -1280 10210 -1210 10220
rect -1280 10130 -1210 10140
rect -960 10210 -890 10220
rect -960 10130 -890 10140
rect -650 10210 -580 10220
rect -650 10130 -580 10140
rect -330 10210 -260 10220
rect -330 10130 -260 10140
rect -20 10210 50 10220
rect -20 10130 50 10140
rect 300 10210 370 10220
rect 300 10130 370 10140
rect 620 10210 690 10220
rect 620 10130 690 10140
rect 930 10210 1000 10220
rect 930 10130 1000 10140
rect 1250 10210 1320 10220
rect 1250 10130 1320 10140
rect 1570 10210 1640 10220
rect 1570 10130 1640 10140
rect 1880 10210 1950 10220
rect 1880 10130 1950 10140
rect 2200 10210 2270 10220
rect 2200 10130 2270 10140
rect 2510 10210 2580 10220
rect 2510 10130 2580 10140
rect 2830 10210 2900 10220
rect 2830 10130 2900 10140
rect 3150 10210 3220 10220
rect 3150 10130 3220 10140
rect 3460 10210 3530 10220
rect 3460 10130 3530 10140
rect 3780 10210 3850 10220
rect 3780 10130 3850 10140
rect 4090 10210 4160 10220
rect 4090 10130 4160 10140
rect 4410 10210 4480 10220
rect 4410 10130 4480 10140
rect 4730 10210 4800 10220
rect 4730 10130 4800 10140
rect 5040 10210 5110 10220
rect 5040 10130 5110 10140
rect 9560 10210 9780 10230
rect 9560 10140 9580 10210
rect 9650 10140 9780 10210
rect -5940 10030 -5920 10100
rect -5850 10030 -5720 10100
rect -5940 10010 -5720 10030
rect 9560 10100 9780 10140
rect 9560 10030 9690 10100
rect 9760 10030 9780 10100
rect 9560 10010 9780 10030
rect -1150 9840 -1020 9850
rect -1150 9770 -1120 9840
rect -1050 9770 -1020 9840
rect -1150 9600 -1020 9770
rect -810 9840 -740 9850
rect -810 9760 -740 9770
rect -490 9840 -420 9850
rect -490 9760 -420 9770
rect -170 9840 -100 9850
rect -170 9760 -100 9770
rect 140 9840 210 9850
rect 140 9760 210 9770
rect 460 9840 530 9850
rect 460 9760 530 9770
rect 770 9840 840 9850
rect 770 9760 840 9770
rect 1090 9840 1160 9850
rect 1090 9760 1160 9770
rect 1410 9840 1480 9850
rect 1410 9760 1480 9770
rect 1720 9840 1790 9850
rect 1720 9760 1790 9770
rect 2040 9840 2110 9850
rect 2040 9760 2110 9770
rect 2360 9840 2430 9850
rect 2360 9760 2430 9770
rect 2670 9840 2740 9850
rect 2670 9760 2740 9770
rect 2990 9840 3060 9850
rect 2990 9760 3060 9770
rect 3300 9840 3370 9850
rect 3300 9760 3370 9770
rect 3620 9840 3690 9850
rect 3620 9760 3690 9770
rect 3940 9840 4010 9850
rect 3940 9760 4010 9770
rect 4250 9840 4320 9850
rect 4250 9760 4320 9770
rect 4570 9840 4640 9850
rect 4570 9760 4640 9770
rect 4860 9840 4990 9850
rect 4860 9770 4890 9840
rect 4960 9770 4990 9840
rect -1150 9530 -1120 9600
rect -1050 9530 -1020 9600
rect -1150 9230 -1020 9530
rect -810 9600 -740 9610
rect -810 9520 -740 9530
rect -490 9600 -420 9610
rect -490 9520 -420 9530
rect -170 9600 -100 9610
rect -170 9520 -100 9530
rect 140 9600 210 9610
rect 140 9520 210 9530
rect 460 9600 530 9610
rect 460 9520 530 9530
rect 770 9600 840 9610
rect 770 9520 840 9530
rect 1090 9600 1160 9610
rect 1090 9520 1160 9530
rect 1410 9600 1480 9610
rect 1410 9520 1480 9530
rect 1720 9600 1790 9610
rect 1720 9520 1790 9530
rect 2040 9600 2110 9610
rect 2040 9520 2110 9530
rect 2360 9600 2430 9610
rect 2360 9520 2430 9530
rect 2670 9600 2740 9610
rect 2670 9520 2740 9530
rect 2990 9600 3060 9610
rect 2990 9520 3060 9530
rect 3300 9600 3370 9610
rect 3300 9520 3370 9530
rect 3620 9600 3690 9610
rect 3620 9520 3690 9530
rect 3940 9600 4010 9610
rect 3940 9520 4010 9530
rect 4250 9600 4320 9610
rect 4250 9520 4320 9530
rect 4570 9600 4640 9610
rect 4570 9520 4640 9530
rect 4860 9600 4990 9770
rect 4860 9530 4890 9600
rect 4960 9530 4990 9600
rect -1150 9160 -1120 9230
rect -1050 9160 -1020 9230
rect -4040 8750 -3860 8760
rect -4040 8640 -3860 8650
rect -3620 8750 -3440 8760
rect -3620 8640 -3440 8650
rect -1150 2620 -1020 9160
rect -200 9430 -40 9450
rect -200 9350 -160 9430
rect -80 9350 -40 9430
rect -200 8130 -40 9350
rect 3860 9430 4020 9450
rect 3860 9350 3900 9430
rect 3980 9350 4020 9430
rect 1270 9290 1540 9300
rect 1270 9010 1540 9020
rect 2320 9290 2590 9300
rect 2320 9010 2590 9020
rect 220 8780 290 8790
rect 220 8700 290 8710
rect 540 8780 610 8790
rect 540 8700 610 8710
rect 850 8780 920 8790
rect 850 8700 920 8710
rect 1170 8780 1240 8790
rect 1170 8700 1240 8710
rect 1490 8780 1560 8790
rect 1490 8700 1560 8710
rect 1800 8780 1870 8790
rect 1800 8700 1870 8710
rect 2120 8780 2190 8790
rect 2120 8700 2190 8710
rect 2440 8780 2510 8790
rect 2440 8700 2510 8710
rect 2750 8780 2820 8790
rect 2750 8700 2820 8710
rect 3070 8780 3140 8790
rect 3070 8700 3140 8710
rect 3380 8780 3450 8790
rect 3380 8700 3450 8710
rect 220 8570 290 8580
rect 220 8490 290 8500
rect 540 8570 610 8580
rect 540 8490 610 8500
rect 850 8570 920 8580
rect 850 8490 920 8500
rect 1170 8570 1240 8580
rect 1170 8490 1240 8500
rect 1490 8570 1560 8580
rect 1490 8490 1560 8500
rect 1800 8570 1870 8580
rect 1800 8490 1870 8500
rect 2120 8570 2190 8580
rect 2120 8490 2190 8500
rect 2440 8570 2510 8580
rect 2440 8490 2510 8500
rect 2750 8570 2820 8580
rect 2750 8490 2820 8500
rect 3070 8570 3140 8580
rect 3070 8490 3140 8500
rect 3380 8570 3450 8580
rect 3380 8490 3450 8500
rect -200 8050 -160 8130
rect -80 8050 -40 8130
rect 380 8140 450 8150
rect 380 8060 450 8070
rect 700 8140 770 8150
rect 700 8060 770 8070
rect 1010 8140 1080 8150
rect 1010 8060 1080 8070
rect 1330 8140 1400 8150
rect 1330 8060 1400 8070
rect 1650 8140 1720 8150
rect 1650 8060 1720 8070
rect 1960 8140 2030 8150
rect 1960 8060 2030 8070
rect 2280 8140 2350 8150
rect 2280 8060 2350 8070
rect 2590 8140 2660 8150
rect 2590 8060 2660 8070
rect 2910 8140 2980 8150
rect 2910 8060 2980 8070
rect 3230 8140 3300 8150
rect 3230 8060 3300 8070
rect 3540 8140 3610 8150
rect 3540 8060 3610 8070
rect 3860 8130 4020 9350
rect -200 7950 -40 8050
rect -200 7870 -160 7950
rect -80 7870 -40 7950
rect 3860 8050 3900 8130
rect 3980 8050 4020 8130
rect 3860 7950 4020 8050
rect -200 5660 -40 7870
rect 380 7930 450 7940
rect 380 7850 450 7860
rect 700 7930 770 7940
rect 700 7850 770 7860
rect 1010 7930 1080 7940
rect 1010 7850 1080 7860
rect 1330 7930 1400 7940
rect 1330 7850 1400 7860
rect 1650 7930 1720 7940
rect 1650 7850 1720 7860
rect 1960 7930 2030 7940
rect 1960 7850 2030 7860
rect 2280 7930 2350 7940
rect 2280 7850 2350 7860
rect 2590 7930 2660 7940
rect 2590 7850 2660 7860
rect 2910 7930 2980 7940
rect 2910 7850 2980 7860
rect 3230 7930 3300 7940
rect 3230 7850 3300 7860
rect 3540 7930 3610 7940
rect 3540 7850 3610 7860
rect 3860 7870 3900 7950
rect 3980 7870 4020 7950
rect 1040 7680 1300 7690
rect 1040 7410 1300 7420
rect 2540 7680 2800 7690
rect 2540 7410 2800 7420
rect 220 7230 290 7240
rect 220 7150 290 7160
rect 540 7230 610 7240
rect 540 7150 610 7160
rect 850 7230 920 7240
rect 850 7150 920 7160
rect 1170 7230 1240 7240
rect 1170 7150 1240 7160
rect 1490 7230 1560 7240
rect 1490 7150 1560 7160
rect 1800 7230 1870 7240
rect 1800 7150 1870 7160
rect 2120 7230 2190 7240
rect 2120 7150 2190 7160
rect 2430 7230 2500 7240
rect 2430 7150 2500 7160
rect 2750 7230 2820 7240
rect 2750 7150 2820 7160
rect 3070 7230 3140 7240
rect 3070 7150 3140 7160
rect 3380 7230 3450 7240
rect 3380 7150 3450 7160
rect 220 7020 290 7030
rect 220 6940 290 6950
rect 540 7020 610 7030
rect 540 6940 610 6950
rect 850 7020 920 7030
rect 850 6940 920 6950
rect 1170 7020 1240 7030
rect 1170 6940 1240 6950
rect 1490 7020 1560 7030
rect 1490 6940 1560 6950
rect 1800 7020 1870 7030
rect 1800 6940 1870 6950
rect 2120 7020 2190 7030
rect 2120 6940 2190 6950
rect 2430 7020 2500 7030
rect 2430 6940 2500 6950
rect 2750 7020 2820 7030
rect 2750 6940 2820 6950
rect 3070 7020 3140 7030
rect 3070 6940 3140 6950
rect 3380 7020 3450 7030
rect 3380 6940 3450 6950
rect 380 6600 450 6610
rect 380 6520 450 6530
rect 670 6600 800 6610
rect 670 6530 700 6600
rect 770 6530 800 6600
rect 380 6390 450 6400
rect 380 6310 450 6320
rect 670 6390 800 6530
rect 1010 6600 1080 6610
rect 1010 6520 1080 6530
rect 1330 6600 1400 6610
rect 1330 6520 1400 6530
rect 1640 6600 1710 6610
rect 1640 6520 1710 6530
rect 1960 6600 2030 6610
rect 1960 6520 2030 6530
rect 2280 6600 2350 6610
rect 2280 6520 2350 6530
rect 2590 6600 2660 6610
rect 2590 6520 2660 6530
rect 2910 6600 2980 6610
rect 2910 6520 2980 6530
rect 3190 6600 3320 6610
rect 3190 6530 3220 6600
rect 3290 6530 3320 6600
rect 670 6320 700 6390
rect 770 6320 800 6390
rect -200 5540 -180 5660
rect -60 5540 -40 5660
rect -200 5440 -40 5540
rect -200 5320 -180 5440
rect -60 5320 -40 5440
rect -200 5300 -40 5320
rect 40 5100 200 5120
rect 40 4980 60 5100
rect 180 4980 200 5100
rect 40 4880 200 4980
rect 40 4760 60 4880
rect 180 4760 200 4880
rect 40 4140 200 4760
rect 40 4020 60 4140
rect 180 4020 200 4140
rect 40 3920 200 4020
rect 40 3800 60 3920
rect 180 3800 200 3920
rect -1150 2550 -1120 2620
rect -1050 2550 -1020 2620
rect -1150 2460 -1020 2550
rect -1150 2390 -1120 2460
rect -1050 2390 -1020 2460
rect -1150 2370 -1020 2390
rect -500 2780 -100 2900
rect -500 2670 -480 2780
rect -370 2670 -230 2780
rect -120 2670 -100 2780
rect -500 1670 -100 2670
rect -500 1560 -480 1670
rect -370 1560 -230 1670
rect -120 1560 -100 1670
rect -500 1260 -100 1560
rect -500 1150 -480 1260
rect -370 1150 -230 1260
rect -120 1150 -100 1260
rect -500 150 -100 1150
rect 40 1110 200 3800
rect 670 3570 800 6320
rect 1010 6390 1080 6400
rect 1010 6310 1080 6320
rect 1330 6390 1400 6400
rect 1330 6310 1400 6320
rect 1640 6390 1710 6400
rect 1640 6310 1710 6320
rect 1960 6390 2030 6400
rect 1960 6310 2030 6320
rect 2280 6390 2350 6400
rect 2280 6310 2350 6320
rect 2590 6390 2660 6400
rect 2590 6310 2660 6320
rect 2910 6390 2980 6400
rect 2910 6310 2980 6320
rect 3190 6390 3320 6530
rect 3540 6600 3610 6610
rect 3540 6520 3610 6530
rect 3190 6320 3220 6390
rect 3290 6320 3320 6390
rect 1320 5670 1390 5680
rect 1320 5590 1390 5600
rect 1640 5670 1710 5680
rect 1640 5590 1710 5600
rect 1950 5670 2020 5680
rect 1950 5590 2020 5600
rect 2270 5670 2340 5680
rect 2270 5590 2340 5600
rect 1320 5380 1390 5390
rect 1320 5300 1390 5310
rect 1640 5380 1710 5390
rect 1640 5300 1710 5310
rect 1950 5380 2020 5390
rect 1950 5300 2020 5310
rect 2270 5380 2340 5390
rect 2270 5300 2340 5310
rect 1480 5110 1550 5120
rect 1480 5030 1550 5040
rect 1790 5110 1860 5120
rect 1790 5030 1860 5040
rect 2110 5110 2180 5120
rect 2110 5030 2180 5040
rect 2430 5110 2500 5120
rect 2430 5030 2500 5040
rect 1480 4820 1550 4830
rect 1480 4740 1550 4750
rect 1790 4820 1860 4830
rect 1790 4740 1860 4750
rect 2110 4820 2180 4830
rect 2110 4740 2180 4750
rect 2430 4820 2500 4830
rect 2430 4740 2500 4750
rect 1780 4580 2040 4590
rect 1780 4310 2040 4320
rect 1320 4150 1390 4160
rect 1320 4070 1390 4080
rect 1640 4150 1710 4160
rect 1640 4070 1710 4080
rect 1950 4150 2020 4160
rect 1950 4070 2020 4080
rect 2270 4150 2340 4160
rect 2270 4070 2340 4080
rect 1320 3860 1390 3870
rect 1320 3780 1390 3790
rect 1640 3860 1710 3870
rect 1640 3780 1710 3790
rect 1950 3860 2020 3870
rect 1950 3780 2020 3790
rect 2270 3860 2340 3870
rect 2270 3780 2340 3790
rect 670 3500 700 3570
rect 770 3500 800 3570
rect 1480 3590 1550 3600
rect 1480 3510 1550 3520
rect 1790 3590 1860 3600
rect 1790 3510 1860 3520
rect 2110 3590 2180 3600
rect 2110 3510 2180 3520
rect 2430 3590 2500 3600
rect 2430 3510 2500 3520
rect 3190 3570 3320 6320
rect 3540 6390 3610 6400
rect 3540 6310 3610 6320
rect 3860 5660 4020 7870
rect 3860 5540 3880 5660
rect 4000 5540 4020 5660
rect 3860 5440 4020 5540
rect 3860 5320 3880 5440
rect 4000 5320 4020 5440
rect 3860 5300 4020 5320
rect 4860 9230 4990 9530
rect 4860 9160 4890 9230
rect 4960 9160 4990 9230
rect 670 3320 800 3500
rect 670 3250 700 3320
rect 770 3250 800 3320
rect 3190 3500 3220 3570
rect 3290 3500 3320 3570
rect 3190 3320 3320 3500
rect 670 3220 800 3250
rect 1480 3300 1550 3310
rect 1480 3220 1550 3230
rect 1790 3300 1860 3310
rect 1790 3220 1860 3230
rect 2110 3300 2180 3310
rect 2110 3220 2180 3230
rect 2430 3300 2500 3310
rect 2430 3220 2500 3230
rect 3190 3250 3220 3320
rect 3290 3250 3320 3320
rect 3190 3220 3320 3250
rect 3620 5100 3780 5120
rect 3620 4980 3640 5100
rect 3760 4980 3780 5100
rect 3620 4880 3780 4980
rect 3620 4760 3640 4880
rect 3760 4760 3780 4880
rect 3620 4140 3780 4760
rect 3620 4020 3640 4140
rect 3760 4020 3780 4140
rect 3620 3920 3780 4020
rect 3620 3800 3640 3920
rect 3760 3800 3780 3920
rect 1780 3060 2040 3070
rect 1780 2790 2040 2800
rect 330 2630 400 2640
rect 330 2550 400 2560
rect 850 2630 920 2640
rect 850 2550 920 2560
rect 1360 2630 1430 2640
rect 1360 2550 1430 2560
rect 1880 2630 1950 2640
rect 1880 2550 1950 2560
rect 2390 2630 2460 2640
rect 2390 2550 2460 2560
rect 2910 2630 2980 2640
rect 2910 2550 2980 2560
rect 3430 2630 3500 2640
rect 3430 2550 3500 2560
rect 330 2450 400 2460
rect 330 2370 400 2380
rect 850 2450 920 2460
rect 850 2370 920 2380
rect 1360 2450 1430 2460
rect 1360 2370 1430 2380
rect 1880 2450 1950 2460
rect 1880 2370 1950 2380
rect 2390 2450 2460 2460
rect 2390 2370 2460 2380
rect 2910 2450 2980 2460
rect 2910 2370 2980 2380
rect 3430 2450 3500 2460
rect 3430 2370 3500 2380
rect 590 1960 660 1970
rect 590 1880 660 1890
rect 1100 1960 1170 1970
rect 1100 1880 1170 1890
rect 1620 1960 1690 1970
rect 1620 1880 1690 1890
rect 2140 1960 2210 1970
rect 2140 1880 2210 1890
rect 2650 1960 2720 1970
rect 2650 1880 2720 1890
rect 3170 1960 3240 1970
rect 3170 1880 3240 1890
rect 590 1780 660 1790
rect 590 1700 660 1710
rect 1100 1780 1170 1790
rect 1100 1700 1170 1710
rect 1620 1780 1690 1790
rect 1620 1700 1690 1710
rect 2140 1780 2210 1790
rect 2140 1700 2210 1710
rect 2650 1780 2720 1790
rect 2650 1700 2720 1710
rect 3170 1780 3240 1790
rect 3170 1700 3240 1710
rect 1790 1540 2040 1550
rect 1790 1280 2040 1290
rect 40 1040 70 1110
rect 140 1040 200 1110
rect 40 930 200 1040
rect 590 1110 660 1120
rect 590 1030 660 1040
rect 1100 1110 1170 1120
rect 1100 1030 1170 1040
rect 1620 1110 1690 1120
rect 1620 1030 1690 1040
rect 2130 1110 2200 1120
rect 2130 1030 2200 1040
rect 2650 1110 2720 1120
rect 2650 1030 2720 1040
rect 3170 1110 3240 1120
rect 3170 1030 3240 1040
rect 3620 1110 3780 3800
rect 3620 1040 3680 1110
rect 3750 1040 3780 1110
rect 40 860 70 930
rect 140 860 200 930
rect 40 850 200 860
rect 590 930 660 940
rect 590 850 660 860
rect 1100 930 1170 940
rect 1100 850 1170 860
rect 1620 930 1690 940
rect 1620 850 1690 860
rect 2130 930 2200 940
rect 2130 850 2200 860
rect 2650 930 2720 940
rect 2650 850 2720 860
rect 3170 930 3240 940
rect 3170 850 3240 860
rect 3620 930 3780 1040
rect 3620 860 3680 930
rect 3750 860 3780 930
rect 3620 850 3780 860
rect 3900 2780 4300 2900
rect 3900 2670 3920 2780
rect 4030 2670 4170 2780
rect 4280 2670 4300 2780
rect 3900 1670 4300 2670
rect 4860 2620 4990 9160
rect 7210 8750 7390 8760
rect 7210 8640 7390 8650
rect 7630 8750 7810 8760
rect 7630 8640 7810 8650
rect 4860 2550 4890 2620
rect 4960 2550 4990 2620
rect 4860 2460 4990 2550
rect 4860 2390 4890 2460
rect 4960 2390 4990 2460
rect 4860 2370 4990 2390
rect 3900 1560 3920 1670
rect 4030 1560 4170 1670
rect 4280 1560 4300 1670
rect 3900 1260 4300 1560
rect 3900 1150 3920 1260
rect 4030 1150 4170 1260
rect 4280 1150 4300 1260
rect 330 440 400 450
rect 330 360 400 370
rect 840 440 910 450
rect 840 360 910 370
rect 1360 440 1430 450
rect 1360 360 1430 370
rect 1880 440 1950 450
rect 1880 360 1950 370
rect 2390 440 2460 450
rect 2390 360 2460 370
rect 2910 440 2980 450
rect 2910 360 2980 370
rect 3420 440 3490 450
rect 3420 360 3490 370
rect 330 260 400 270
rect 330 180 400 190
rect 840 260 910 270
rect 840 180 910 190
rect 1360 260 1430 270
rect 1360 180 1430 190
rect 1880 260 1950 270
rect 1880 180 1950 190
rect 2390 260 2460 270
rect 2390 180 2460 190
rect 2910 260 2980 270
rect 2910 180 2980 190
rect 3420 260 3490 270
rect 3420 180 3490 190
rect -500 40 -480 150
rect -370 40 -230 150
rect -120 40 -100 150
rect -500 -100 -100 40
rect 3900 150 4300 1150
rect 3900 40 3920 150
rect 4030 40 4170 150
rect 4280 40 4300 150
rect 1790 10 2040 20
rect 3900 -100 4300 40
rect 1790 -250 2040 -240
<< via2 >>
rect 1270 10660 1540 10930
rect 2320 10660 2590 10930
rect -1280 10380 -1210 10450
rect -960 10380 -890 10450
rect -650 10380 -580 10450
rect -330 10380 -260 10450
rect -20 10380 50 10450
rect 300 10380 370 10450
rect 620 10380 690 10450
rect 930 10380 1000 10450
rect 1250 10380 1320 10450
rect 1570 10380 1640 10450
rect 1880 10380 1950 10450
rect 2200 10380 2270 10450
rect 2510 10380 2580 10450
rect 2830 10380 2900 10450
rect 3150 10380 3220 10450
rect 3460 10380 3530 10450
rect 3780 10380 3850 10450
rect 4090 10380 4160 10450
rect 4410 10380 4480 10450
rect 4730 10380 4800 10450
rect 5040 10380 5110 10450
rect -5810 10140 -5740 10210
rect -1280 10140 -1210 10210
rect -960 10140 -890 10210
rect -650 10140 -580 10210
rect -330 10140 -260 10210
rect -20 10140 50 10210
rect 300 10140 370 10210
rect 620 10140 690 10210
rect 930 10140 1000 10210
rect 1250 10140 1320 10210
rect 1570 10140 1640 10210
rect 1880 10140 1950 10210
rect 2200 10140 2270 10210
rect 2510 10140 2580 10210
rect 2830 10140 2900 10210
rect 3150 10140 3220 10210
rect 3460 10140 3530 10210
rect 3780 10140 3850 10210
rect 4090 10140 4160 10210
rect 4410 10140 4480 10210
rect 4730 10140 4800 10210
rect 5040 10140 5110 10210
rect 9580 10140 9650 10210
rect -5920 10030 -5850 10100
rect 9690 10030 9760 10100
rect -1120 9770 -1050 9840
rect -810 9770 -740 9840
rect -490 9770 -420 9840
rect -170 9770 -100 9840
rect 140 9770 210 9840
rect 460 9770 530 9840
rect 770 9770 840 9840
rect 1090 9770 1160 9840
rect 1410 9770 1480 9840
rect 1720 9770 1790 9840
rect 2040 9770 2110 9840
rect 2360 9770 2430 9840
rect 2670 9770 2740 9840
rect 2990 9770 3060 9840
rect 3300 9770 3370 9840
rect 3620 9770 3690 9840
rect 3940 9770 4010 9840
rect 4250 9770 4320 9840
rect 4570 9770 4640 9840
rect 4890 9770 4960 9840
rect -1120 9530 -1050 9600
rect -810 9530 -740 9600
rect -490 9530 -420 9600
rect -170 9530 -100 9600
rect 140 9530 210 9600
rect 460 9530 530 9600
rect 770 9530 840 9600
rect 1090 9530 1160 9600
rect 1410 9530 1480 9600
rect 1720 9530 1790 9600
rect 2040 9530 2110 9600
rect 2360 9530 2430 9600
rect 2670 9530 2740 9600
rect 2990 9530 3060 9600
rect 3300 9530 3370 9600
rect 3620 9530 3690 9600
rect 3940 9530 4010 9600
rect 4250 9530 4320 9600
rect 4570 9530 4640 9600
rect 4890 9530 4960 9600
rect -1120 9160 -1050 9230
rect -4040 8650 -3860 8750
rect -3620 8650 -3440 8750
rect 1270 9020 1540 9290
rect 2320 9020 2590 9290
rect 220 8710 290 8780
rect 540 8710 610 8780
rect 850 8710 920 8780
rect 1170 8710 1240 8780
rect 1490 8710 1560 8780
rect 1800 8710 1870 8780
rect 2120 8710 2190 8780
rect 2440 8710 2510 8780
rect 2750 8710 2820 8780
rect 3070 8710 3140 8780
rect 3380 8710 3450 8780
rect 220 8500 290 8570
rect 540 8500 610 8570
rect 850 8500 920 8570
rect 1170 8500 1240 8570
rect 1490 8500 1560 8570
rect 1800 8500 1870 8570
rect 2120 8500 2190 8570
rect 2440 8500 2510 8570
rect 2750 8500 2820 8570
rect 3070 8500 3140 8570
rect 3380 8500 3450 8570
rect -160 8050 -80 8130
rect 380 8070 450 8140
rect 700 8070 770 8140
rect 1010 8070 1080 8140
rect 1330 8070 1400 8140
rect 1650 8070 1720 8140
rect 1960 8070 2030 8140
rect 2280 8070 2350 8140
rect 2590 8070 2660 8140
rect 2910 8070 2980 8140
rect 3230 8070 3300 8140
rect 3540 8070 3610 8140
rect -160 7870 -80 7950
rect 3900 8050 3980 8130
rect 380 7860 450 7930
rect 700 7860 770 7930
rect 1010 7860 1080 7930
rect 1330 7860 1400 7930
rect 1650 7860 1720 7930
rect 1960 7860 2030 7930
rect 2280 7860 2350 7930
rect 2590 7860 2660 7930
rect 2910 7860 2980 7930
rect 3230 7860 3300 7930
rect 3540 7860 3610 7930
rect 3900 7870 3980 7950
rect 1040 7420 1300 7680
rect 2540 7420 2800 7680
rect 220 7160 290 7230
rect 540 7160 610 7230
rect 850 7160 920 7230
rect 1170 7160 1240 7230
rect 1490 7160 1560 7230
rect 1800 7160 1870 7230
rect 2120 7160 2190 7230
rect 2430 7160 2500 7230
rect 2750 7160 2820 7230
rect 3070 7160 3140 7230
rect 3380 7160 3450 7230
rect 220 6950 290 7020
rect 540 6950 610 7020
rect 850 6950 920 7020
rect 1170 6950 1240 7020
rect 1490 6950 1560 7020
rect 1800 6950 1870 7020
rect 2120 6950 2190 7020
rect 2430 6950 2500 7020
rect 2750 6950 2820 7020
rect 3070 6950 3140 7020
rect 3380 6950 3450 7020
rect 380 6530 450 6600
rect 700 6530 770 6600
rect 380 6320 450 6390
rect 1010 6530 1080 6600
rect 1330 6530 1400 6600
rect 1640 6530 1710 6600
rect 1960 6530 2030 6600
rect 2280 6530 2350 6600
rect 2590 6530 2660 6600
rect 2910 6530 2980 6600
rect 3220 6530 3290 6600
rect 700 6320 770 6390
rect -180 5540 -60 5660
rect -180 5320 -60 5440
rect 60 4980 180 5100
rect 60 4760 180 4880
rect 60 4020 180 4140
rect 60 3800 180 3920
rect -1120 2550 -1050 2620
rect -1120 2390 -1050 2460
rect 1010 6320 1080 6390
rect 1330 6320 1400 6390
rect 1640 6320 1710 6390
rect 1960 6320 2030 6390
rect 2280 6320 2350 6390
rect 2590 6320 2660 6390
rect 2910 6320 2980 6390
rect 3540 6530 3610 6600
rect 3220 6320 3290 6390
rect 1320 5600 1390 5670
rect 1640 5600 1710 5670
rect 1950 5600 2020 5670
rect 2270 5600 2340 5670
rect 1320 5310 1390 5380
rect 1640 5310 1710 5380
rect 1950 5310 2020 5380
rect 2270 5310 2340 5380
rect 1480 5040 1550 5110
rect 1790 5040 1860 5110
rect 2110 5040 2180 5110
rect 2430 5040 2500 5110
rect 1480 4750 1550 4820
rect 1790 4750 1860 4820
rect 2110 4750 2180 4820
rect 2430 4750 2500 4820
rect 1780 4320 2040 4580
rect 1320 4080 1390 4150
rect 1640 4080 1710 4150
rect 1950 4080 2020 4150
rect 2270 4080 2340 4150
rect 1320 3790 1390 3860
rect 1640 3790 1710 3860
rect 1950 3790 2020 3860
rect 2270 3790 2340 3860
rect 700 3500 770 3570
rect 1480 3520 1550 3590
rect 1790 3520 1860 3590
rect 2110 3520 2180 3590
rect 2430 3520 2500 3590
rect 3540 6320 3610 6390
rect 3880 5540 4000 5660
rect 3880 5320 4000 5440
rect 4890 9160 4960 9230
rect 700 3250 770 3320
rect 3220 3500 3290 3570
rect 1480 3230 1550 3300
rect 1790 3230 1860 3300
rect 2110 3230 2180 3300
rect 2430 3230 2500 3300
rect 3220 3250 3290 3320
rect 3640 4980 3760 5100
rect 3640 4760 3760 4880
rect 3640 4020 3760 4140
rect 3640 3800 3760 3920
rect 1780 2800 2040 3060
rect 330 2560 400 2630
rect 850 2560 920 2630
rect 1360 2560 1430 2630
rect 1880 2560 1950 2630
rect 2390 2560 2460 2630
rect 2910 2560 2980 2630
rect 3430 2560 3500 2630
rect 330 2380 400 2450
rect 850 2380 920 2450
rect 1360 2380 1430 2450
rect 1880 2380 1950 2450
rect 2390 2380 2460 2450
rect 2910 2380 2980 2450
rect 3430 2380 3500 2450
rect 590 1890 660 1960
rect 1100 1890 1170 1960
rect 1620 1890 1690 1960
rect 2140 1890 2210 1960
rect 2650 1890 2720 1960
rect 3170 1890 3240 1960
rect 590 1710 660 1780
rect 1100 1710 1170 1780
rect 1620 1710 1690 1780
rect 2140 1710 2210 1780
rect 2650 1710 2720 1780
rect 3170 1710 3240 1780
rect 1790 1290 2040 1540
rect 70 1040 140 1110
rect 590 1040 660 1110
rect 1100 1040 1170 1110
rect 1620 1040 1690 1110
rect 2130 1040 2200 1110
rect 2650 1040 2720 1110
rect 3170 1040 3240 1110
rect 3680 1040 3750 1110
rect 70 860 140 930
rect 590 860 660 930
rect 1100 860 1170 930
rect 1620 860 1690 930
rect 2130 860 2200 930
rect 2650 860 2720 930
rect 3170 860 3240 930
rect 3680 860 3750 930
rect 7210 8650 7390 8750
rect 7630 8650 7810 8750
rect 4890 2550 4960 2620
rect 4890 2390 4960 2460
rect 330 370 400 440
rect 840 370 910 440
rect 1360 370 1430 440
rect 1880 370 1950 440
rect 2390 370 2460 440
rect 2910 370 2980 440
rect 3420 370 3490 440
rect 330 190 400 260
rect 840 190 910 260
rect 1360 190 1430 260
rect 1880 190 1950 260
rect 2390 190 2460 260
rect 2910 190 2980 260
rect 3420 190 3490 260
rect 1790 -240 2040 10
<< metal3 >>
rect 1260 10930 1550 10935
rect 1260 10660 1270 10930
rect 1540 10660 1550 10930
rect 1260 10655 1550 10660
rect 2310 10930 2600 10935
rect 2310 10660 2320 10930
rect 2590 10660 2600 10930
rect 2310 10655 2600 10660
rect -1280 10455 5110 10460
rect -1290 10450 5120 10455
rect -1290 10380 -1280 10450
rect -1210 10380 -960 10450
rect -890 10430 -650 10450
rect -580 10380 -330 10450
rect -260 10380 -20 10450
rect 50 10380 300 10450
rect 370 10380 620 10450
rect 690 10380 930 10450
rect 1000 10420 1250 10450
rect -1290 10375 -900 10380
rect -5940 10210 -5720 10230
rect -1280 10215 -900 10375
rect -5940 10140 -5810 10210
rect -5740 10140 -5720 10210
rect -5940 10100 -5720 10140
rect -1290 10210 -900 10215
rect -650 10210 1000 10380
rect -1290 10140 -1280 10210
rect -1210 10140 -960 10210
rect -890 10140 -650 10180
rect -580 10140 -330 10210
rect -260 10140 -20 10210
rect 50 10140 300 10210
rect 370 10140 620 10210
rect 690 10140 930 10210
rect 1320 10380 1570 10450
rect 1640 10380 1880 10450
rect 1950 10380 2200 10450
rect 2270 10380 2510 10450
rect 2580 10420 2830 10450
rect 1250 10210 2580 10380
rect 1000 10140 1250 10170
rect 1320 10140 1570 10210
rect 1640 10140 1880 10210
rect 1950 10140 2200 10210
rect 2270 10140 2510 10210
rect 2900 10380 3150 10450
rect 3220 10380 3460 10450
rect 3530 10380 3780 10450
rect 3850 10380 4090 10450
rect 4160 10380 4410 10450
rect 4480 10420 4730 10450
rect 2830 10210 4480 10380
rect 2580 10140 2830 10170
rect 2900 10140 3150 10210
rect 3220 10140 3460 10210
rect 3530 10140 3780 10210
rect 3850 10140 4090 10210
rect 4160 10140 4410 10210
rect 4800 10380 5040 10450
rect 5110 10380 5120 10450
rect 4730 10375 5120 10380
rect 4730 10215 5110 10375
rect 4730 10210 5120 10215
rect 4480 10140 4730 10170
rect 4800 10140 5040 10210
rect 5110 10140 5120 10210
rect -1290 10135 5120 10140
rect 9560 10210 9780 10230
rect 9560 10140 9580 10210
rect 9650 10140 9780 10210
rect -1280 10130 5110 10135
rect -5940 10030 -5920 10100
rect -5850 10030 -5720 10100
rect -5940 10010 -5720 10030
rect 9560 10100 9780 10140
rect 9560 10030 9690 10100
rect 9760 10030 9780 10100
rect 9560 10010 9780 10030
rect -1280 9840 5110 9850
rect -1280 9770 -1120 9840
rect -1050 9770 -810 9840
rect -740 9770 -490 9840
rect -420 9770 -170 9840
rect -100 9770 140 9840
rect 210 9770 460 9840
rect 530 9770 770 9840
rect 840 9770 1090 9840
rect 1160 9770 1410 9840
rect 1480 9770 1720 9840
rect 1790 9770 2040 9840
rect 2110 9770 2360 9840
rect 2430 9770 2670 9840
rect 2740 9770 2990 9840
rect 3060 9770 3300 9840
rect 3370 9770 3620 9840
rect 3690 9770 3940 9840
rect 4010 9770 4250 9840
rect 4320 9770 4570 9840
rect 4640 9770 4890 9840
rect 4960 9770 5110 9840
rect -1280 9600 5110 9770
rect -1280 9530 -1120 9600
rect -1050 9530 -810 9600
rect -740 9530 -490 9600
rect -420 9530 -170 9600
rect -100 9530 140 9600
rect 210 9530 460 9600
rect 530 9530 770 9600
rect 840 9530 1090 9600
rect 1160 9530 1410 9600
rect 1480 9530 1720 9600
rect 1790 9530 2040 9600
rect 2110 9530 2360 9600
rect 2430 9530 2670 9600
rect 2740 9530 2990 9600
rect 3060 9530 3300 9600
rect 3370 9530 3620 9600
rect 3690 9530 3940 9600
rect 4010 9530 4250 9600
rect 4320 9530 4570 9600
rect 4640 9530 4890 9600
rect 4960 9530 5110 9600
rect -1280 9520 5110 9530
rect 1260 9290 1550 9295
rect -2050 9250 -1020 9270
rect -2050 9150 -2030 9250
rect -1940 9150 -1840 9250
rect -1750 9230 -1020 9250
rect -1750 9160 -1120 9230
rect -1050 9160 -1020 9230
rect -1750 9150 -1020 9160
rect -2050 9130 -1020 9150
rect 1260 9020 1270 9290
rect 1540 9020 1550 9290
rect 1260 9015 1550 9020
rect 2310 9290 2600 9295
rect 2310 9020 2320 9290
rect 2590 9020 2600 9290
rect 4860 9250 5880 9270
rect 4860 9230 5580 9250
rect 4860 9160 4890 9230
rect 4960 9160 5580 9230
rect 4860 9150 5580 9160
rect 5670 9150 5770 9250
rect 5860 9150 5880 9250
rect 4860 9130 5880 9150
rect 2310 9015 2600 9020
rect 220 8785 3610 8790
rect 210 8780 3610 8785
rect -4050 8750 -3850 8755
rect -4050 8650 -4040 8750
rect -3860 8650 -3850 8750
rect -4050 8645 -3850 8650
rect -3630 8750 -3430 8755
rect -3630 8650 -3620 8750
rect -3440 8650 -3430 8750
rect 210 8710 220 8780
rect 290 8710 540 8780
rect 610 8770 850 8780
rect 920 8710 1170 8780
rect 1240 8710 1490 8780
rect 1560 8710 1800 8780
rect 1870 8770 2120 8780
rect 2190 8710 2440 8780
rect 2510 8710 2750 8780
rect 2820 8710 3070 8780
rect 3140 8770 3380 8780
rect 3450 8710 3610 8780
rect 210 8705 600 8710
rect -3630 8645 -3430 8650
rect 220 8575 600 8705
rect 210 8570 600 8575
rect 860 8570 1870 8710
rect 2130 8570 3130 8710
rect 3390 8570 3610 8710
rect 7200 8750 7400 8755
rect 7200 8650 7210 8750
rect 7390 8650 7400 8750
rect 7200 8645 7400 8650
rect 7620 8750 7820 8755
rect 7620 8650 7630 8750
rect 7810 8650 7820 8750
rect 7620 8645 7820 8650
rect 210 8500 220 8570
rect 290 8500 540 8570
rect 610 8500 850 8510
rect 920 8500 1170 8570
rect 1240 8500 1490 8570
rect 1560 8500 1800 8570
rect 1870 8500 2120 8510
rect 2190 8500 2440 8570
rect 2510 8500 2750 8570
rect 2820 8500 3070 8570
rect 3140 8500 3380 8510
rect 3450 8500 3610 8570
rect 210 8495 3610 8500
rect 220 8490 3610 8495
rect -200 8140 4020 8150
rect -200 8130 380 8140
rect -200 8050 -160 8130
rect -80 8070 380 8130
rect 450 8070 700 8140
rect 770 8070 1010 8140
rect 1080 8070 1330 8140
rect 1400 8070 1650 8140
rect 1720 8070 1960 8140
rect 2030 8070 2280 8140
rect 2350 8070 2590 8140
rect 2660 8070 2910 8140
rect 2980 8070 3230 8140
rect 3300 8070 3540 8140
rect 3610 8130 4020 8140
rect 3610 8070 3900 8130
rect -80 8050 3900 8070
rect 3980 8050 4020 8130
rect -200 7950 4020 8050
rect -200 7870 -160 7950
rect -80 7930 3900 7950
rect -80 7870 380 7930
rect -200 7860 380 7870
rect 450 7860 700 7930
rect 770 7860 1010 7930
rect 1080 7860 1330 7930
rect 1400 7860 1650 7930
rect 1720 7860 1960 7930
rect 2030 7860 2280 7930
rect 2350 7860 2590 7930
rect 2660 7860 2910 7930
rect 2980 7860 3230 7930
rect 3300 7860 3540 7930
rect 3610 7870 3900 7930
rect 3980 7870 4020 7950
rect 3610 7860 4020 7870
rect -200 7850 4020 7860
rect 1030 7680 1310 7685
rect 1030 7420 1040 7680
rect 1300 7420 1310 7680
rect 1030 7415 1310 7420
rect 2530 7680 2810 7685
rect 2530 7420 2540 7680
rect 2800 7420 2810 7680
rect 2530 7415 2810 7420
rect 220 7235 3610 7240
rect 210 7230 3610 7235
rect 210 7160 220 7230
rect 290 7160 540 7230
rect 610 7220 850 7230
rect 920 7160 1170 7230
rect 1240 7160 1490 7230
rect 1560 7160 1800 7230
rect 1870 7220 2120 7230
rect 2190 7160 2430 7230
rect 2500 7160 2750 7230
rect 2820 7160 3070 7230
rect 3140 7220 3380 7230
rect 3450 7160 3610 7230
rect 210 7155 600 7160
rect 220 7025 600 7155
rect 210 7020 600 7025
rect 860 7020 1870 7160
rect 2130 7020 3130 7160
rect 3390 7020 3610 7160
rect 210 6950 220 7020
rect 290 6950 540 7020
rect 610 6950 850 6960
rect 920 6950 1170 7020
rect 1240 6950 1490 7020
rect 1560 6950 1800 7020
rect 1870 6950 2120 6960
rect 2190 6950 2430 7020
rect 2500 6950 2750 7020
rect 2820 6950 3070 7020
rect 3140 6950 3380 6960
rect 3450 6950 3610 7020
rect 210 6945 3610 6950
rect 220 6940 3610 6945
rect 220 6605 3610 6610
rect 220 6600 3620 6605
rect 220 6530 380 6600
rect 450 6530 700 6600
rect 770 6530 1010 6600
rect 1080 6530 1330 6600
rect 1400 6530 1640 6600
rect 1710 6530 1960 6600
rect 2030 6530 2280 6600
rect 2350 6530 2590 6600
rect 2660 6530 2910 6600
rect 2980 6530 3220 6600
rect 3290 6530 3540 6600
rect 3610 6530 3620 6600
rect 220 6525 3620 6530
rect 220 6395 3610 6525
rect 220 6390 3620 6395
rect 220 6320 380 6390
rect 450 6320 700 6390
rect 770 6320 1010 6390
rect 1080 6320 1330 6390
rect 1400 6320 1640 6390
rect 1710 6320 1960 6390
rect 2030 6320 2280 6390
rect 2350 6320 2590 6390
rect 2660 6320 2910 6390
rect 2980 6320 3220 6390
rect 3290 6320 3540 6390
rect 3610 6320 3620 6390
rect 220 6315 3620 6320
rect 220 6310 3610 6315
rect -200 5670 4020 5680
rect -200 5660 1320 5670
rect -200 5540 -180 5660
rect -60 5600 1320 5660
rect 1390 5600 1640 5670
rect 1710 5600 1950 5670
rect 2020 5600 2270 5670
rect 2340 5660 4020 5670
rect 2340 5600 3880 5660
rect -60 5540 3880 5600
rect 4000 5540 4020 5660
rect -200 5440 4020 5540
rect -200 5320 -180 5440
rect -60 5380 3880 5440
rect -60 5320 1320 5380
rect -200 5310 1320 5320
rect 1390 5310 1640 5380
rect 1710 5310 1950 5380
rect 2020 5310 2270 5380
rect 2340 5320 3880 5380
rect 4000 5320 4020 5440
rect 2340 5310 4020 5320
rect -200 5300 4020 5310
rect 40 5110 3780 5120
rect 40 5100 1480 5110
rect 40 4980 60 5100
rect 180 5040 1480 5100
rect 1550 5040 1790 5110
rect 1860 5040 2110 5110
rect 2180 5040 2430 5110
rect 2500 5100 3780 5110
rect 2500 5040 3640 5100
rect 180 4980 3640 5040
rect 3760 4980 3780 5100
rect 40 4880 3780 4980
rect 40 4760 60 4880
rect 180 4820 3640 4880
rect 180 4760 1480 4820
rect 40 4750 1480 4760
rect 1550 4750 1790 4820
rect 1860 4750 2110 4820
rect 2180 4750 2430 4820
rect 2500 4760 3640 4820
rect 3760 4760 3780 4880
rect 2500 4750 3780 4760
rect 40 4740 3780 4750
rect 1770 4580 2050 4585
rect 1770 4320 1780 4580
rect 2040 4320 2050 4580
rect 1770 4315 2050 4320
rect 40 4150 3780 4160
rect 40 4140 1320 4150
rect 40 4020 60 4140
rect 180 4080 1320 4140
rect 1390 4080 1640 4150
rect 1710 4080 1950 4150
rect 2020 4080 2270 4150
rect 2340 4140 3780 4150
rect 2340 4080 3640 4140
rect 180 4020 3640 4080
rect 3760 4020 3780 4140
rect 40 3920 3780 4020
rect 40 3800 60 3920
rect 180 3860 3640 3920
rect 180 3800 1320 3860
rect 40 3790 1320 3800
rect 1390 3790 1640 3860
rect 1710 3790 1950 3860
rect 2020 3790 2270 3860
rect 2340 3800 3640 3860
rect 3760 3800 3780 3920
rect 2340 3790 3780 3800
rect 40 3780 3780 3790
rect 670 3590 3320 3600
rect 670 3570 1480 3590
rect 670 3500 700 3570
rect 770 3520 1480 3570
rect 1550 3520 1790 3590
rect 1860 3520 2110 3590
rect 2180 3520 2430 3590
rect 2500 3570 3320 3590
rect 2500 3520 3220 3570
rect 770 3500 3220 3520
rect 3290 3500 3320 3570
rect 670 3320 3320 3500
rect 670 3250 700 3320
rect 770 3300 3220 3320
rect 770 3250 1480 3300
rect 670 3230 1480 3250
rect 1550 3230 1790 3300
rect 1860 3230 2110 3300
rect 2180 3230 2430 3300
rect 2500 3250 3220 3300
rect 3290 3250 3320 3320
rect 2500 3230 3320 3250
rect 670 3220 3320 3230
rect 1770 3060 2050 3065
rect 1770 2800 1780 3060
rect 2040 2800 2050 3060
rect 1770 2795 2050 2800
rect -1150 2630 4990 2640
rect -1150 2620 330 2630
rect -1150 2550 -1120 2620
rect -1050 2560 330 2620
rect 400 2560 850 2630
rect 920 2560 1360 2630
rect 1430 2560 1880 2630
rect 1950 2560 2390 2630
rect 2460 2560 2910 2630
rect 2980 2560 3430 2630
rect 3500 2620 4990 2630
rect 3500 2560 4890 2620
rect -1050 2550 4890 2560
rect 4960 2550 4990 2620
rect -1150 2460 4990 2550
rect -1150 2390 -1120 2460
rect -1050 2450 4890 2460
rect -1050 2390 330 2450
rect -1150 2380 330 2390
rect 400 2380 850 2450
rect 920 2380 1360 2450
rect 1430 2380 1880 2450
rect 1950 2380 2390 2450
rect 2460 2380 2910 2450
rect 2980 2380 3430 2450
rect 3500 2390 4890 2450
rect 4960 2390 4990 2460
rect 3500 2380 4990 2390
rect -1150 2370 4990 2380
rect 330 1960 3500 1970
rect 330 1890 590 1960
rect 660 1890 760 1960
rect 330 1780 760 1890
rect 330 1710 590 1780
rect 660 1710 760 1780
rect 1010 1890 1100 1960
rect 1170 1890 1620 1960
rect 1690 1890 2140 1960
rect 2210 1890 2650 1960
rect 2720 1890 2820 1960
rect 1010 1780 2820 1890
rect 1010 1710 1100 1780
rect 1170 1710 1620 1780
rect 1690 1710 2140 1780
rect 2210 1710 2650 1780
rect 2720 1710 2820 1780
rect 3070 1890 3170 1960
rect 3240 1890 3500 1960
rect 3070 1780 3500 1890
rect 3070 1710 3170 1780
rect 3240 1710 3500 1780
rect 330 1700 3500 1710
rect 1780 1540 2050 1545
rect 1780 1290 1790 1540
rect 2040 1290 2050 1540
rect 1780 1285 2050 1290
rect 70 1115 3750 1120
rect 60 1110 3760 1115
rect 60 1040 70 1110
rect 140 1040 590 1110
rect 660 1040 1100 1110
rect 1170 1040 1620 1110
rect 1690 1040 2130 1110
rect 2200 1040 2650 1110
rect 2720 1040 3170 1110
rect 3240 1040 3680 1110
rect 3750 1040 3760 1110
rect 60 1035 3760 1040
rect 70 935 3750 1035
rect 60 930 3760 935
rect 60 860 70 930
rect 140 860 590 930
rect 660 860 1100 930
rect 1170 860 1620 930
rect 1690 860 2130 930
rect 2200 860 2650 930
rect 2720 860 3170 930
rect 3240 860 3680 930
rect 3750 860 3760 930
rect 60 855 3760 860
rect 70 850 3750 855
rect 70 440 3750 450
rect 70 370 330 440
rect 400 370 500 440
rect 70 260 500 370
rect 70 190 330 260
rect 400 190 500 260
rect 750 370 840 440
rect 910 370 1360 440
rect 1430 370 1880 440
rect 1950 370 2390 440
rect 2460 370 2910 440
rect 2980 370 3080 440
rect 750 260 3080 370
rect 750 190 840 260
rect 910 190 1360 260
rect 1430 190 1880 260
rect 1950 190 2390 260
rect 2460 190 2910 260
rect 2980 190 3080 260
rect 3330 370 3420 440
rect 3490 370 3750 440
rect 3330 260 3750 370
rect 3330 190 3420 260
rect 3490 190 3750 260
rect 70 180 3750 190
rect 1780 10 2050 15
rect 1780 -240 1790 10
rect 2040 -240 2050 10
rect 1780 -245 2050 -240
<< via3 >>
rect 1270 10660 1540 10930
rect 2320 10660 2590 10930
rect -900 10380 -890 10430
rect -890 10380 -650 10430
rect -5810 10140 -5740 10210
rect -900 10210 -650 10380
rect -900 10180 -890 10210
rect -890 10180 -650 10210
rect 1000 10170 1250 10420
rect 2580 10170 2830 10420
rect 4480 10170 4730 10420
rect 9580 10140 9650 10210
rect -5920 10030 -5850 10100
rect 9690 10030 9760 10100
rect -2030 9150 -1940 9250
rect -1840 9150 -1750 9250
rect 1270 9020 1540 9290
rect 2320 9020 2590 9290
rect 5580 9150 5670 9250
rect 5770 9150 5860 9250
rect -4040 8650 -3860 8750
rect -3620 8650 -3440 8750
rect 600 8710 610 8770
rect 610 8710 850 8770
rect 850 8710 860 8770
rect 1870 8710 2120 8770
rect 2120 8710 2130 8770
rect 3130 8710 3140 8770
rect 3140 8710 3380 8770
rect 3380 8710 3390 8770
rect 600 8570 860 8710
rect 1870 8570 2130 8710
rect 3130 8570 3390 8710
rect 7210 8650 7390 8750
rect 7630 8650 7810 8750
rect 600 8510 610 8570
rect 610 8510 850 8570
rect 850 8510 860 8570
rect 1870 8510 2120 8570
rect 2120 8510 2130 8570
rect 3130 8510 3140 8570
rect 3140 8510 3380 8570
rect 3380 8510 3390 8570
rect 1040 7420 1300 7680
rect 2540 7420 2800 7680
rect 600 7160 610 7220
rect 610 7160 850 7220
rect 850 7160 860 7220
rect 1870 7160 2120 7220
rect 2120 7160 2130 7220
rect 3130 7160 3140 7220
rect 3140 7160 3380 7220
rect 3380 7160 3390 7220
rect 600 7020 860 7160
rect 1870 7020 2130 7160
rect 3130 7020 3390 7160
rect 600 6960 610 7020
rect 610 6960 850 7020
rect 850 6960 860 7020
rect 1870 6960 2120 7020
rect 2120 6960 2130 7020
rect 3130 6960 3140 7020
rect 3140 6960 3380 7020
rect 3380 6960 3390 7020
rect 1780 4320 2040 4580
rect 1780 2800 2040 3060
rect 760 1710 1010 1960
rect 2820 1710 3070 1960
rect 1790 1290 2040 1540
rect 500 190 750 440
rect 3080 190 3330 440
rect 1790 -240 2040 10
<< metal4 >>
rect -5940 16310 9780 16550
rect -5940 10210 -5720 16310
rect -2350 14480 9150 14840
rect -5940 10140 -5810 10210
rect -5740 10140 -5720 10210
rect -5940 10100 -5720 10140
rect -5940 10030 -5920 10100
rect -5850 10030 -5720 10100
rect -5940 10010 -5720 10030
rect -2050 9250 -1730 14480
rect 1269 10930 1541 10931
rect 1269 10660 1270 10930
rect 1540 10660 1541 10930
rect 1269 10659 1541 10660
rect 2319 10930 2591 10931
rect 2319 10660 2320 10930
rect 2590 10660 2591 10930
rect 2319 10659 2591 10660
rect -901 10430 -649 10431
rect -901 10180 -900 10430
rect -650 10180 -649 10430
rect -901 10179 -649 10180
rect 999 10420 1251 10421
rect 999 10170 1000 10420
rect 1250 10170 1251 10420
rect 999 10169 1251 10170
rect 2579 10420 2831 10421
rect 2579 10170 2580 10420
rect 2830 10170 2831 10420
rect 2579 10169 2831 10170
rect 4479 10420 4731 10421
rect 4479 10170 4480 10420
rect 4730 10170 4731 10420
rect 4479 10169 4731 10170
rect -2050 9150 -2030 9250
rect -1940 9150 -1840 9250
rect -1750 9150 -1730 9250
rect -2050 9130 -1730 9150
rect 1269 9290 1541 9291
rect 1269 9020 1270 9290
rect 1540 9020 1541 9290
rect 1269 9019 1541 9020
rect 2319 9290 2591 9291
rect 2319 9020 2320 9290
rect 2590 9020 2591 9290
rect 5560 9250 5880 14480
rect 9560 10210 9780 16310
rect 9560 10140 9580 10210
rect 9650 10140 9780 10210
rect 9560 10100 9780 10140
rect 9560 10030 9690 10100
rect 9760 10030 9780 10100
rect 9560 10010 9780 10030
rect 5560 9150 5580 9250
rect 5670 9150 5770 9250
rect 5860 9150 5880 9250
rect 5560 9130 5880 9150
rect 2319 9019 2591 9020
rect -4070 8750 -3410 8780
rect -4070 8650 -4040 8750
rect -3860 8650 -3620 8750
rect -3440 8650 -3410 8750
rect -4070 1310 -3410 8650
rect 599 8770 861 8771
rect 599 8510 600 8770
rect 860 8510 861 8770
rect 599 8509 861 8510
rect 1869 8770 2131 8771
rect 1869 8510 1870 8770
rect 2130 8510 2131 8770
rect 1869 8509 2131 8510
rect 3129 8770 3391 8771
rect 3129 8510 3130 8770
rect 3390 8510 3391 8770
rect 3129 8509 3391 8510
rect 7180 8750 7840 8780
rect 7180 8650 7210 8750
rect 7390 8650 7630 8750
rect 7810 8650 7840 8750
rect 1039 7680 1301 7681
rect 1039 7420 1040 7680
rect 1300 7420 1301 7680
rect 1039 7419 1301 7420
rect 2539 7680 2801 7681
rect 2539 7420 2540 7680
rect 2800 7420 2801 7680
rect 2539 7419 2801 7420
rect 599 7220 861 7221
rect 599 6960 600 7220
rect 860 6960 861 7220
rect 599 6959 861 6960
rect 1869 7220 2131 7221
rect 1869 6960 1870 7220
rect 2130 6960 2131 7220
rect 1869 6959 2131 6960
rect 3129 7220 3391 7221
rect 3129 6960 3130 7220
rect 3390 6960 3391 7220
rect 3129 6959 3391 6960
rect 1779 4580 2041 4581
rect 1779 4320 1780 4580
rect 2040 4320 2041 4580
rect 1779 4319 2041 4320
rect 1779 3060 2041 3061
rect 1779 2800 1780 3060
rect 2040 2800 2041 3060
rect 1779 2799 2041 2800
rect 759 1960 1011 1961
rect 759 1710 760 1960
rect 1010 1710 1011 1960
rect 759 1709 1011 1710
rect 2819 1960 3071 1961
rect 2819 1710 2820 1960
rect 3070 1710 3071 1960
rect 2819 1709 3071 1710
rect -4070 1070 -4040 1310
rect -3800 1070 -3680 1310
rect -3440 1070 -3410 1310
rect 1789 1540 2041 1541
rect 1789 1290 1790 1540
rect 2040 1290 2041 1540
rect 1789 1289 2041 1290
rect 7180 1310 7840 8650
rect -4070 970 -3410 1070
rect -4070 730 -4040 970
rect -3800 730 -3680 970
rect -3440 730 -3410 970
rect -4070 700 -3410 730
rect 7180 1070 7210 1310
rect 7450 1070 7570 1310
rect 7810 1070 7840 1310
rect 7180 970 7840 1070
rect 7180 730 7210 970
rect 7450 730 7570 970
rect 7810 730 7840 970
rect 7180 700 7840 730
rect 499 440 751 441
rect 499 190 500 440
rect 750 190 751 440
rect 499 189 751 190
rect 3079 440 3331 441
rect 3079 190 3080 440
rect 3330 190 3331 440
rect 3079 189 3331 190
rect 1789 10 2041 11
rect 1789 -240 1790 10
rect 2040 -240 2041 10
rect 1789 -241 2041 -240
<< via4 >>
rect 1270 10660 1540 10930
rect 2320 10660 2590 10930
rect -900 10180 -650 10430
rect 1000 10170 1250 10420
rect 2580 10170 2830 10420
rect 4480 10170 4730 10420
rect 1270 9020 1540 9290
rect 2320 9020 2590 9290
rect 600 8510 860 8770
rect 1870 8510 2130 8770
rect 3130 8510 3390 8770
rect 1040 7420 1300 7680
rect 2540 7420 2800 7680
rect 600 6960 860 7220
rect 1870 6960 2130 7220
rect 3130 6960 3390 7220
rect 1780 4320 2040 4580
rect 1780 2800 2040 3060
rect 760 1710 1010 1960
rect 2820 1710 3070 1960
rect -4040 1070 -3800 1310
rect -3680 1070 -3440 1310
rect 1790 1290 2040 1540
rect -4040 730 -3800 970
rect -3680 730 -3440 970
rect 7210 1070 7450 1310
rect 7570 1070 7810 1310
rect 7210 730 7450 970
rect 7570 730 7810 970
rect 500 190 750 440
rect 3080 190 3330 440
rect 1790 -240 2040 10
<< metal5 >>
rect 1240 10930 2620 10980
rect 1240 10660 1270 10930
rect 1540 10660 2320 10930
rect 2590 10660 2620 10930
rect 1240 10460 2620 10660
rect -930 10430 4770 10460
rect -930 10180 -900 10430
rect -650 10420 4770 10430
rect -650 10180 1000 10420
rect -930 10170 1000 10180
rect 1250 10170 2580 10420
rect 2830 10170 4480 10420
rect 4730 10170 4770 10420
rect -930 10130 4770 10170
rect 1240 9290 2620 10130
rect 1240 9020 1270 9290
rect 1540 9020 2320 9290
rect 2590 9020 2620 9290
rect 1240 8800 2620 9020
rect 450 8770 3430 8800
rect 450 8510 600 8770
rect 860 8510 1870 8770
rect 2130 8510 3130 8770
rect 3390 8510 3430 8770
rect 450 8480 3430 8510
rect 1240 7710 2620 8480
rect 1010 7680 2830 7710
rect 1010 7420 1040 7680
rect 1300 7420 2540 7680
rect 2800 7420 2830 7680
rect 1010 7250 2830 7420
rect 560 7220 3430 7250
rect 560 6960 600 7220
rect 860 6960 1870 7220
rect 2130 6960 3130 7220
rect 3390 6960 3430 7220
rect 560 6930 3430 6960
rect 1690 4580 2130 4620
rect 1690 4320 1780 4580
rect 2040 4320 2130 4580
rect 1690 3060 2130 4320
rect 1690 2800 1780 3060
rect 2040 2800 2130 3060
rect 1690 2000 2130 2800
rect -920 1960 4720 2000
rect -920 1710 760 1960
rect 1010 1710 2820 1960
rect 3070 1710 4720 1960
rect -920 1540 4720 1710
rect -920 1340 1790 1540
rect -4070 1310 1790 1340
rect -4070 1070 -4040 1310
rect -3800 1070 -3680 1310
rect -3440 1290 1790 1310
rect 2040 1340 4720 1540
rect 2040 1310 7840 1340
rect 2040 1290 7210 1310
rect -3440 1070 7210 1290
rect 7450 1070 7570 1310
rect 7810 1070 7840 1310
rect -4070 970 7840 1070
rect -4070 730 -4040 970
rect -3800 730 -3680 970
rect -3440 730 7210 970
rect 7450 730 7570 970
rect 7810 730 7840 970
rect -4070 700 7840 730
rect -920 440 4720 700
rect -920 190 500 440
rect 750 190 3080 440
rect 3330 190 4720 440
rect -920 150 4720 190
rect 1700 10 2140 150
rect 1700 -240 1790 10
rect 2040 -240 2140 10
rect 1700 -310 2140 -240
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_0
timestamp 1683391037
transform 0 -1 7610 1 0 14670
box -1750 -1700 1749 1700
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_1
timestamp 1683391037
transform 0 -1 3810 1 0 14670
box -1750 -1700 1749 1700
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_2
timestamp 1683391037
transform 0 -1 10 1 0 14670
box -1750 -1700 1749 1700
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_3
timestamp 1683391037
transform 0 -1 -3790 1 0 14670
box -1750 -1700 1749 1700
use sky130_fd_pr__nfet_01v8_EJ3ASN  sky130_fd_pr__nfet_01v8_EJ3ASN_0
timestamp 1683391037
transform 1 0 1911 0 1 5211
box -720 -710 720 710
use sky130_fd_pr__nfet_01v8_EJ3ASN  sky130_fd_pr__nfet_01v8_EJ3ASN_1
timestamp 1683391037
transform 1 0 1911 0 1 3691
box -720 -710 720 710
use sky130_fd_pr__nfet_01v8_JEXVB9  sky130_fd_pr__nfet_01v8_JEXVB9_0
timestamp 1683391037
transform 1 0 1915 0 1 2170
box -1715 -710 1715 710
use sky130_fd_pr__nfet_01v8_JT3SH9  sky130_fd_pr__nfet_01v8_JT3SH9_0
timestamp 1683391037
transform 1 0 1913 0 1 650
box -1973 -710 1973 710
use sky130_fd_pr__pfet_01v8_9F67JW  sky130_fd_pr__pfet_01v8_9F67JW_0
timestamp 1683391037
transform 1 0 1917 0 1 9989
box -3327 -719 3327 719
use sky130_fd_pr__pfet_01v8_49C6SK  sky130_fd_pr__pfet_01v8_49C6SK_0
timestamp 1683391037
transform 1 0 1916 0 1 8319
box -1826 -719 1826 719
use sky130_fd_pr__pfet_01v8_GNAJ57  sky130_fd_pr__pfet_01v8_GNAJ57_0
timestamp 1683391037
transform 1 0 1916 0 1 6779
box -1826 -719 1826 719
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_0
timestamp 1683391037
transform 0 1 -3615 -1 0 10846
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_1
timestamp 1683391037
transform 0 1 -3615 -1 0 9386
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_2
timestamp 1683391037
transform 0 1 7455 -1 0 9386
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_3
timestamp 1683391037
transform 0 1 7455 -1 0 10846
box -739 -1598 739 1598
<< end >>
