magic
tech sky130A
magscale 1 2
timestamp 1676503286
<< nwell >>
rect -296 -7517 296 7517
<< pmos >>
rect -100 6298 100 7298
rect -100 5062 100 6062
rect -100 3826 100 4826
rect -100 2590 100 3590
rect -100 1354 100 2354
rect -100 118 100 1118
rect -100 -1118 100 -118
rect -100 -2354 100 -1354
rect -100 -3590 100 -2590
rect -100 -4826 100 -3826
rect -100 -6062 100 -5062
rect -100 -7298 100 -6298
<< pdiff >>
rect -158 7286 -100 7298
rect -158 6310 -146 7286
rect -112 6310 -100 7286
rect -158 6298 -100 6310
rect 100 7286 158 7298
rect 100 6310 112 7286
rect 146 6310 158 7286
rect 100 6298 158 6310
rect -158 6050 -100 6062
rect -158 5074 -146 6050
rect -112 5074 -100 6050
rect -158 5062 -100 5074
rect 100 6050 158 6062
rect 100 5074 112 6050
rect 146 5074 158 6050
rect 100 5062 158 5074
rect -158 4814 -100 4826
rect -158 3838 -146 4814
rect -112 3838 -100 4814
rect -158 3826 -100 3838
rect 100 4814 158 4826
rect 100 3838 112 4814
rect 146 3838 158 4814
rect 100 3826 158 3838
rect -158 3578 -100 3590
rect -158 2602 -146 3578
rect -112 2602 -100 3578
rect -158 2590 -100 2602
rect 100 3578 158 3590
rect 100 2602 112 3578
rect 146 2602 158 3578
rect 100 2590 158 2602
rect -158 2342 -100 2354
rect -158 1366 -146 2342
rect -112 1366 -100 2342
rect -158 1354 -100 1366
rect 100 2342 158 2354
rect 100 1366 112 2342
rect 146 1366 158 2342
rect 100 1354 158 1366
rect -158 1106 -100 1118
rect -158 130 -146 1106
rect -112 130 -100 1106
rect -158 118 -100 130
rect 100 1106 158 1118
rect 100 130 112 1106
rect 146 130 158 1106
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -1106 -146 -130
rect -112 -1106 -100 -130
rect -158 -1118 -100 -1106
rect 100 -130 158 -118
rect 100 -1106 112 -130
rect 146 -1106 158 -130
rect 100 -1118 158 -1106
rect -158 -1366 -100 -1354
rect -158 -2342 -146 -1366
rect -112 -2342 -100 -1366
rect -158 -2354 -100 -2342
rect 100 -1366 158 -1354
rect 100 -2342 112 -1366
rect 146 -2342 158 -1366
rect 100 -2354 158 -2342
rect -158 -2602 -100 -2590
rect -158 -3578 -146 -2602
rect -112 -3578 -100 -2602
rect -158 -3590 -100 -3578
rect 100 -2602 158 -2590
rect 100 -3578 112 -2602
rect 146 -3578 158 -2602
rect 100 -3590 158 -3578
rect -158 -3838 -100 -3826
rect -158 -4814 -146 -3838
rect -112 -4814 -100 -3838
rect -158 -4826 -100 -4814
rect 100 -3838 158 -3826
rect 100 -4814 112 -3838
rect 146 -4814 158 -3838
rect 100 -4826 158 -4814
rect -158 -5074 -100 -5062
rect -158 -6050 -146 -5074
rect -112 -6050 -100 -5074
rect -158 -6062 -100 -6050
rect 100 -5074 158 -5062
rect 100 -6050 112 -5074
rect 146 -6050 158 -5074
rect 100 -6062 158 -6050
rect -158 -6310 -100 -6298
rect -158 -7286 -146 -6310
rect -112 -7286 -100 -6310
rect -158 -7298 -100 -7286
rect 100 -6310 158 -6298
rect 100 -7286 112 -6310
rect 146 -7286 158 -6310
rect 100 -7298 158 -7286
<< pdiffc >>
rect -146 6310 -112 7286
rect 112 6310 146 7286
rect -146 5074 -112 6050
rect 112 5074 146 6050
rect -146 3838 -112 4814
rect 112 3838 146 4814
rect -146 2602 -112 3578
rect 112 2602 146 3578
rect -146 1366 -112 2342
rect 112 1366 146 2342
rect -146 130 -112 1106
rect 112 130 146 1106
rect -146 -1106 -112 -130
rect 112 -1106 146 -130
rect -146 -2342 -112 -1366
rect 112 -2342 146 -1366
rect -146 -3578 -112 -2602
rect 112 -3578 146 -2602
rect -146 -4814 -112 -3838
rect 112 -4814 146 -3838
rect -146 -6050 -112 -5074
rect 112 -6050 146 -5074
rect -146 -7286 -112 -6310
rect 112 -7286 146 -6310
<< nsubdiff >>
rect -260 7447 -164 7481
rect 164 7447 260 7481
rect -260 7385 -226 7447
rect 226 7385 260 7447
rect -260 -7447 -226 -7385
rect 226 -7447 260 -7385
rect -260 -7481 -164 -7447
rect 164 -7481 260 -7447
<< nsubdiffcont >>
rect -164 7447 164 7481
rect -260 -7385 -226 7385
rect 226 -7385 260 7385
rect -164 -7481 164 -7447
<< poly >>
rect -100 7379 100 7395
rect -100 7345 -84 7379
rect 84 7345 100 7379
rect -100 7298 100 7345
rect -100 6251 100 6298
rect -100 6217 -84 6251
rect 84 6217 100 6251
rect -100 6201 100 6217
rect -100 6143 100 6159
rect -100 6109 -84 6143
rect 84 6109 100 6143
rect -100 6062 100 6109
rect -100 5015 100 5062
rect -100 4981 -84 5015
rect 84 4981 100 5015
rect -100 4965 100 4981
rect -100 4907 100 4923
rect -100 4873 -84 4907
rect 84 4873 100 4907
rect -100 4826 100 4873
rect -100 3779 100 3826
rect -100 3745 -84 3779
rect 84 3745 100 3779
rect -100 3729 100 3745
rect -100 3671 100 3687
rect -100 3637 -84 3671
rect 84 3637 100 3671
rect -100 3590 100 3637
rect -100 2543 100 2590
rect -100 2509 -84 2543
rect 84 2509 100 2543
rect -100 2493 100 2509
rect -100 2435 100 2451
rect -100 2401 -84 2435
rect 84 2401 100 2435
rect -100 2354 100 2401
rect -100 1307 100 1354
rect -100 1273 -84 1307
rect 84 1273 100 1307
rect -100 1257 100 1273
rect -100 1199 100 1215
rect -100 1165 -84 1199
rect 84 1165 100 1199
rect -100 1118 100 1165
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -1165 100 -1118
rect -100 -1199 -84 -1165
rect 84 -1199 100 -1165
rect -100 -1215 100 -1199
rect -100 -1273 100 -1257
rect -100 -1307 -84 -1273
rect 84 -1307 100 -1273
rect -100 -1354 100 -1307
rect -100 -2401 100 -2354
rect -100 -2435 -84 -2401
rect 84 -2435 100 -2401
rect -100 -2451 100 -2435
rect -100 -2509 100 -2493
rect -100 -2543 -84 -2509
rect 84 -2543 100 -2509
rect -100 -2590 100 -2543
rect -100 -3637 100 -3590
rect -100 -3671 -84 -3637
rect 84 -3671 100 -3637
rect -100 -3687 100 -3671
rect -100 -3745 100 -3729
rect -100 -3779 -84 -3745
rect 84 -3779 100 -3745
rect -100 -3826 100 -3779
rect -100 -4873 100 -4826
rect -100 -4907 -84 -4873
rect 84 -4907 100 -4873
rect -100 -4923 100 -4907
rect -100 -4981 100 -4965
rect -100 -5015 -84 -4981
rect 84 -5015 100 -4981
rect -100 -5062 100 -5015
rect -100 -6109 100 -6062
rect -100 -6143 -84 -6109
rect 84 -6143 100 -6109
rect -100 -6159 100 -6143
rect -100 -6217 100 -6201
rect -100 -6251 -84 -6217
rect 84 -6251 100 -6217
rect -100 -6298 100 -6251
rect -100 -7345 100 -7298
rect -100 -7379 -84 -7345
rect 84 -7379 100 -7345
rect -100 -7395 100 -7379
<< polycont >>
rect -84 7345 84 7379
rect -84 6217 84 6251
rect -84 6109 84 6143
rect -84 4981 84 5015
rect -84 4873 84 4907
rect -84 3745 84 3779
rect -84 3637 84 3671
rect -84 2509 84 2543
rect -84 2401 84 2435
rect -84 1273 84 1307
rect -84 1165 84 1199
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1199 84 -1165
rect -84 -1307 84 -1273
rect -84 -2435 84 -2401
rect -84 -2543 84 -2509
rect -84 -3671 84 -3637
rect -84 -3779 84 -3745
rect -84 -4907 84 -4873
rect -84 -5015 84 -4981
rect -84 -6143 84 -6109
rect -84 -6251 84 -6217
rect -84 -7379 84 -7345
<< locali >>
rect -260 7447 -164 7481
rect 164 7447 260 7481
rect -260 7385 -226 7447
rect 226 7385 260 7447
rect -100 7345 -84 7379
rect 84 7345 100 7379
rect -146 7286 -112 7302
rect -146 6294 -112 6310
rect 112 7286 146 7302
rect 112 6294 146 6310
rect -100 6217 -84 6251
rect 84 6217 100 6251
rect -100 6109 -84 6143
rect 84 6109 100 6143
rect -146 6050 -112 6066
rect -146 5058 -112 5074
rect 112 6050 146 6066
rect 112 5058 146 5074
rect -100 4981 -84 5015
rect 84 4981 100 5015
rect -100 4873 -84 4907
rect 84 4873 100 4907
rect -146 4814 -112 4830
rect -146 3822 -112 3838
rect 112 4814 146 4830
rect 112 3822 146 3838
rect -100 3745 -84 3779
rect 84 3745 100 3779
rect -100 3637 -84 3671
rect 84 3637 100 3671
rect -146 3578 -112 3594
rect -146 2586 -112 2602
rect 112 3578 146 3594
rect 112 2586 146 2602
rect -100 2509 -84 2543
rect 84 2509 100 2543
rect -100 2401 -84 2435
rect 84 2401 100 2435
rect -146 2342 -112 2358
rect -146 1350 -112 1366
rect 112 2342 146 2358
rect 112 1350 146 1366
rect -100 1273 -84 1307
rect 84 1273 100 1307
rect -100 1165 -84 1199
rect 84 1165 100 1199
rect -146 1106 -112 1122
rect -146 114 -112 130
rect 112 1106 146 1122
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -1122 -112 -1106
rect 112 -130 146 -114
rect 112 -1122 146 -1106
rect -100 -1199 -84 -1165
rect 84 -1199 100 -1165
rect -100 -1307 -84 -1273
rect 84 -1307 100 -1273
rect -146 -1366 -112 -1350
rect -146 -2358 -112 -2342
rect 112 -1366 146 -1350
rect 112 -2358 146 -2342
rect -100 -2435 -84 -2401
rect 84 -2435 100 -2401
rect -100 -2543 -84 -2509
rect 84 -2543 100 -2509
rect -146 -2602 -112 -2586
rect -146 -3594 -112 -3578
rect 112 -2602 146 -2586
rect 112 -3594 146 -3578
rect -100 -3671 -84 -3637
rect 84 -3671 100 -3637
rect -100 -3779 -84 -3745
rect 84 -3779 100 -3745
rect -146 -3838 -112 -3822
rect -146 -4830 -112 -4814
rect 112 -3838 146 -3822
rect 112 -4830 146 -4814
rect -100 -4907 -84 -4873
rect 84 -4907 100 -4873
rect -100 -5015 -84 -4981
rect 84 -5015 100 -4981
rect -146 -5074 -112 -5058
rect -146 -6066 -112 -6050
rect 112 -5074 146 -5058
rect 112 -6066 146 -6050
rect -100 -6143 -84 -6109
rect 84 -6143 100 -6109
rect -100 -6251 -84 -6217
rect 84 -6251 100 -6217
rect -146 -6310 -112 -6294
rect -146 -7302 -112 -7286
rect 112 -6310 146 -6294
rect 112 -7302 146 -7286
rect -100 -7379 -84 -7345
rect 84 -7379 100 -7345
rect -260 -7447 -226 -7385
rect 226 -7447 260 -7385
rect -260 -7481 -164 -7447
rect 164 -7481 260 -7447
<< viali >>
rect -84 7345 84 7379
rect -146 6310 -112 7286
rect 112 6310 146 7286
rect -84 6217 84 6251
rect -84 6109 84 6143
rect -146 5074 -112 6050
rect 112 5074 146 6050
rect -84 4981 84 5015
rect -84 4873 84 4907
rect -146 3838 -112 4814
rect 112 3838 146 4814
rect -84 3745 84 3779
rect -84 3637 84 3671
rect -146 2602 -112 3578
rect 112 2602 146 3578
rect -84 2509 84 2543
rect -84 2401 84 2435
rect -146 1366 -112 2342
rect 112 1366 146 2342
rect -84 1273 84 1307
rect -84 1165 84 1199
rect -146 130 -112 1106
rect 112 130 146 1106
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1106 -112 -130
rect 112 -1106 146 -130
rect -84 -1199 84 -1165
rect -84 -1307 84 -1273
rect -146 -2342 -112 -1366
rect 112 -2342 146 -1366
rect -84 -2435 84 -2401
rect -84 -2543 84 -2509
rect -146 -3578 -112 -2602
rect 112 -3578 146 -2602
rect -84 -3671 84 -3637
rect -84 -3779 84 -3745
rect -146 -4814 -112 -3838
rect 112 -4814 146 -3838
rect -84 -4907 84 -4873
rect -84 -5015 84 -4981
rect -146 -6050 -112 -5074
rect 112 -6050 146 -5074
rect -84 -6143 84 -6109
rect -84 -6251 84 -6217
rect -146 -7286 -112 -6310
rect 112 -7286 146 -6310
rect -84 -7379 84 -7345
<< metal1 >>
rect -96 7379 96 7385
rect -96 7345 -84 7379
rect 84 7345 96 7379
rect -96 7339 96 7345
rect -152 7286 -106 7298
rect -152 6310 -146 7286
rect -112 6310 -106 7286
rect -152 6298 -106 6310
rect 106 7286 152 7298
rect 106 6310 112 7286
rect 146 6310 152 7286
rect 106 6298 152 6310
rect -96 6251 96 6257
rect -96 6217 -84 6251
rect 84 6217 96 6251
rect -96 6211 96 6217
rect -96 6143 96 6149
rect -96 6109 -84 6143
rect 84 6109 96 6143
rect -96 6103 96 6109
rect -152 6050 -106 6062
rect -152 5074 -146 6050
rect -112 5074 -106 6050
rect -152 5062 -106 5074
rect 106 6050 152 6062
rect 106 5074 112 6050
rect 146 5074 152 6050
rect 106 5062 152 5074
rect -96 5015 96 5021
rect -96 4981 -84 5015
rect 84 4981 96 5015
rect -96 4975 96 4981
rect -96 4907 96 4913
rect -96 4873 -84 4907
rect 84 4873 96 4907
rect -96 4867 96 4873
rect -152 4814 -106 4826
rect -152 3838 -146 4814
rect -112 3838 -106 4814
rect -152 3826 -106 3838
rect 106 4814 152 4826
rect 106 3838 112 4814
rect 146 3838 152 4814
rect 106 3826 152 3838
rect -96 3779 96 3785
rect -96 3745 -84 3779
rect 84 3745 96 3779
rect -96 3739 96 3745
rect -96 3671 96 3677
rect -96 3637 -84 3671
rect 84 3637 96 3671
rect -96 3631 96 3637
rect -152 3578 -106 3590
rect -152 2602 -146 3578
rect -112 2602 -106 3578
rect -152 2590 -106 2602
rect 106 3578 152 3590
rect 106 2602 112 3578
rect 146 2602 152 3578
rect 106 2590 152 2602
rect -96 2543 96 2549
rect -96 2509 -84 2543
rect 84 2509 96 2543
rect -96 2503 96 2509
rect -96 2435 96 2441
rect -96 2401 -84 2435
rect 84 2401 96 2435
rect -96 2395 96 2401
rect -152 2342 -106 2354
rect -152 1366 -146 2342
rect -112 1366 -106 2342
rect -152 1354 -106 1366
rect 106 2342 152 2354
rect 106 1366 112 2342
rect 146 1366 152 2342
rect 106 1354 152 1366
rect -96 1307 96 1313
rect -96 1273 -84 1307
rect 84 1273 96 1307
rect -96 1267 96 1273
rect -96 1199 96 1205
rect -96 1165 -84 1199
rect 84 1165 96 1199
rect -96 1159 96 1165
rect -152 1106 -106 1118
rect -152 130 -146 1106
rect -112 130 -106 1106
rect -152 118 -106 130
rect 106 1106 152 1118
rect 106 130 112 1106
rect 146 130 152 1106
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -1106 -146 -130
rect -112 -1106 -106 -130
rect -152 -1118 -106 -1106
rect 106 -130 152 -118
rect 106 -1106 112 -130
rect 146 -1106 152 -130
rect 106 -1118 152 -1106
rect -96 -1165 96 -1159
rect -96 -1199 -84 -1165
rect 84 -1199 96 -1165
rect -96 -1205 96 -1199
rect -96 -1273 96 -1267
rect -96 -1307 -84 -1273
rect 84 -1307 96 -1273
rect -96 -1313 96 -1307
rect -152 -1366 -106 -1354
rect -152 -2342 -146 -1366
rect -112 -2342 -106 -1366
rect -152 -2354 -106 -2342
rect 106 -1366 152 -1354
rect 106 -2342 112 -1366
rect 146 -2342 152 -1366
rect 106 -2354 152 -2342
rect -96 -2401 96 -2395
rect -96 -2435 -84 -2401
rect 84 -2435 96 -2401
rect -96 -2441 96 -2435
rect -96 -2509 96 -2503
rect -96 -2543 -84 -2509
rect 84 -2543 96 -2509
rect -96 -2549 96 -2543
rect -152 -2602 -106 -2590
rect -152 -3578 -146 -2602
rect -112 -3578 -106 -2602
rect -152 -3590 -106 -3578
rect 106 -2602 152 -2590
rect 106 -3578 112 -2602
rect 146 -3578 152 -2602
rect 106 -3590 152 -3578
rect -96 -3637 96 -3631
rect -96 -3671 -84 -3637
rect 84 -3671 96 -3637
rect -96 -3677 96 -3671
rect -96 -3745 96 -3739
rect -96 -3779 -84 -3745
rect 84 -3779 96 -3745
rect -96 -3785 96 -3779
rect -152 -3838 -106 -3826
rect -152 -4814 -146 -3838
rect -112 -4814 -106 -3838
rect -152 -4826 -106 -4814
rect 106 -3838 152 -3826
rect 106 -4814 112 -3838
rect 146 -4814 152 -3838
rect 106 -4826 152 -4814
rect -96 -4873 96 -4867
rect -96 -4907 -84 -4873
rect 84 -4907 96 -4873
rect -96 -4913 96 -4907
rect -96 -4981 96 -4975
rect -96 -5015 -84 -4981
rect 84 -5015 96 -4981
rect -96 -5021 96 -5015
rect -152 -5074 -106 -5062
rect -152 -6050 -146 -5074
rect -112 -6050 -106 -5074
rect -152 -6062 -106 -6050
rect 106 -5074 152 -5062
rect 106 -6050 112 -5074
rect 146 -6050 152 -5074
rect 106 -6062 152 -6050
rect -96 -6109 96 -6103
rect -96 -6143 -84 -6109
rect 84 -6143 96 -6109
rect -96 -6149 96 -6143
rect -96 -6217 96 -6211
rect -96 -6251 -84 -6217
rect 84 -6251 96 -6217
rect -96 -6257 96 -6251
rect -152 -6310 -106 -6298
rect -152 -7286 -146 -6310
rect -112 -7286 -106 -6310
rect -152 -7298 -106 -7286
rect 106 -6310 152 -6298
rect 106 -7286 112 -6310
rect 146 -7286 152 -6310
rect 106 -7298 152 -7286
rect -96 -7345 96 -7339
rect -96 -7379 -84 -7345
rect 84 -7379 96 -7345
rect -96 -7385 96 -7379
<< properties >>
string FIXED_BBOX -243 -7464 243 7464
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 1 m 12 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
