magic
tech sky130A
magscale 1 2
timestamp 1676748949
<< xpolycontact >>
rect -573 8470 573 8902
rect -573 -8902 573 -8470
<< xpolyres >>
rect -573 -8470 573 8470
<< viali >>
rect -557 8487 557 8884
rect -557 -8884 557 -8487
<< metal1 >>
rect -569 8884 569 8890
rect -569 8487 -557 8884
rect 557 8487 569 8884
rect -569 8481 569 8487
rect -569 -8487 569 -8481
rect -569 -8884 -557 -8487
rect 557 -8884 569 -8487
rect -569 -8890 569 -8884
<< res5p73 >>
rect -575 -8472 575 8472
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 84.7 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 29.629k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
