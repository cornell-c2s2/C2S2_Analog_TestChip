magic
tech sky130A
magscale 1 2
timestamp 1682004261
<< pwell >>
rect -739 -7498 739 7498
<< psubdiff >>
rect -703 7428 -607 7462
rect 607 7428 703 7462
rect -703 7366 -669 7428
rect 669 7366 703 7428
rect -703 -7428 -669 -7366
rect 669 -7428 703 -7366
rect -703 -7462 -607 -7428
rect 607 -7462 703 -7428
<< psubdiffcont >>
rect -607 7428 607 7462
rect -703 -7366 -669 7366
rect 669 -7366 703 7366
rect -607 -7462 607 -7428
<< xpolycontact >>
rect -573 6900 573 7332
rect -573 -7332 573 -6900
<< xpolyres >>
rect -573 -6900 573 6900
<< locali >>
rect -703 7428 -607 7462
rect 607 7428 703 7462
rect -703 7366 -669 7428
rect 669 7366 703 7428
rect -703 -7428 -669 -7366
rect 669 -7428 703 -7366
rect -703 -7462 -607 -7428
rect 607 -7462 703 -7428
<< viali >>
rect -557 6917 557 7314
rect -557 -7314 557 -6917
<< metal1 >>
rect -569 7314 569 7320
rect -569 6917 -557 7314
rect 557 6917 569 7314
rect -569 6911 569 6917
rect -569 -6917 569 -6911
rect -569 -7314 -557 -6917
rect 557 -7314 569 -6917
rect -569 -7320 569 -7314
<< res5p73 >>
rect -575 -6902 575 6902
<< properties >>
string FIXED_BBOX -686 -7445 686 7445
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 69 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 24.149k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
