magic
tech sky130A
timestamp 1683391037
<< pwell >>
rect -123 -2182 123 2182
<< nmos >>
rect -25 1577 25 2077
rect -25 968 25 1468
rect -25 359 25 859
rect -25 -250 25 250
rect -25 -859 25 -359
rect -25 -1468 25 -968
rect -25 -2077 25 -1577
<< ndiff >>
rect -54 2071 -25 2077
rect -54 1583 -48 2071
rect -31 1583 -25 2071
rect -54 1577 -25 1583
rect 25 2071 54 2077
rect 25 1583 31 2071
rect 48 1583 54 2071
rect 25 1577 54 1583
rect -54 1462 -25 1468
rect -54 974 -48 1462
rect -31 974 -25 1462
rect -54 968 -25 974
rect 25 1462 54 1468
rect 25 974 31 1462
rect 48 974 54 1462
rect 25 968 54 974
rect -54 853 -25 859
rect -54 365 -48 853
rect -31 365 -25 853
rect -54 359 -25 365
rect 25 853 54 859
rect 25 365 31 853
rect 48 365 54 853
rect 25 359 54 365
rect -54 244 -25 250
rect -54 -244 -48 244
rect -31 -244 -25 244
rect -54 -250 -25 -244
rect 25 244 54 250
rect 25 -244 31 244
rect 48 -244 54 244
rect 25 -250 54 -244
rect -54 -365 -25 -359
rect -54 -853 -48 -365
rect -31 -853 -25 -365
rect -54 -859 -25 -853
rect 25 -365 54 -359
rect 25 -853 31 -365
rect 48 -853 54 -365
rect 25 -859 54 -853
rect -54 -974 -25 -968
rect -54 -1462 -48 -974
rect -31 -1462 -25 -974
rect -54 -1468 -25 -1462
rect 25 -974 54 -968
rect 25 -1462 31 -974
rect 48 -1462 54 -974
rect 25 -1468 54 -1462
rect -54 -1583 -25 -1577
rect -54 -2071 -48 -1583
rect -31 -2071 -25 -1583
rect -54 -2077 -25 -2071
rect 25 -1583 54 -1577
rect 25 -2071 31 -1583
rect 48 -2071 54 -1583
rect 25 -2077 54 -2071
<< ndiffc >>
rect -48 1583 -31 2071
rect 31 1583 48 2071
rect -48 974 -31 1462
rect 31 974 48 1462
rect -48 365 -31 853
rect 31 365 48 853
rect -48 -244 -31 244
rect 31 -244 48 244
rect -48 -853 -31 -365
rect 31 -853 48 -365
rect -48 -1462 -31 -974
rect 31 -1462 48 -974
rect -48 -2071 -31 -1583
rect 31 -2071 48 -1583
<< psubdiff >>
rect -105 2147 -57 2164
rect 57 2147 105 2164
rect -105 2116 -88 2147
rect 88 2116 105 2147
rect -105 -2147 -88 -2116
rect 88 -2147 105 -2116
rect -105 -2164 -57 -2147
rect 57 -2164 105 -2147
<< psubdiffcont >>
rect -57 2147 57 2164
rect -105 -2116 -88 2116
rect 88 -2116 105 2116
rect -57 -2164 57 -2147
<< poly >>
rect -25 2113 25 2121
rect -25 2096 -17 2113
rect 17 2096 25 2113
rect -25 2077 25 2096
rect -25 1558 25 1577
rect -25 1541 -17 1558
rect 17 1541 25 1558
rect -25 1533 25 1541
rect -25 1504 25 1512
rect -25 1487 -17 1504
rect 17 1487 25 1504
rect -25 1468 25 1487
rect -25 949 25 968
rect -25 932 -17 949
rect 17 932 25 949
rect -25 924 25 932
rect -25 895 25 903
rect -25 878 -17 895
rect 17 878 25 895
rect -25 859 25 878
rect -25 340 25 359
rect -25 323 -17 340
rect 17 323 25 340
rect -25 315 25 323
rect -25 286 25 294
rect -25 269 -17 286
rect 17 269 25 286
rect -25 250 25 269
rect -25 -269 25 -250
rect -25 -286 -17 -269
rect 17 -286 25 -269
rect -25 -294 25 -286
rect -25 -323 25 -315
rect -25 -340 -17 -323
rect 17 -340 25 -323
rect -25 -359 25 -340
rect -25 -878 25 -859
rect -25 -895 -17 -878
rect 17 -895 25 -878
rect -25 -903 25 -895
rect -25 -932 25 -924
rect -25 -949 -17 -932
rect 17 -949 25 -932
rect -25 -968 25 -949
rect -25 -1487 25 -1468
rect -25 -1504 -17 -1487
rect 17 -1504 25 -1487
rect -25 -1512 25 -1504
rect -25 -1541 25 -1533
rect -25 -1558 -17 -1541
rect 17 -1558 25 -1541
rect -25 -1577 25 -1558
rect -25 -2096 25 -2077
rect -25 -2113 -17 -2096
rect 17 -2113 25 -2096
rect -25 -2121 25 -2113
<< polycont >>
rect -17 2096 17 2113
rect -17 1541 17 1558
rect -17 1487 17 1504
rect -17 932 17 949
rect -17 878 17 895
rect -17 323 17 340
rect -17 269 17 286
rect -17 -286 17 -269
rect -17 -340 17 -323
rect -17 -895 17 -878
rect -17 -949 17 -932
rect -17 -1504 17 -1487
rect -17 -1558 17 -1541
rect -17 -2113 17 -2096
<< locali >>
rect -105 2147 -57 2164
rect 57 2147 105 2164
rect -105 2116 -88 2147
rect 88 2116 105 2147
rect -25 2096 -17 2113
rect 17 2096 25 2113
rect -48 2071 -31 2079
rect -48 1575 -31 1583
rect 31 2071 48 2079
rect 31 1575 48 1583
rect -25 1541 -17 1558
rect 17 1541 25 1558
rect -25 1487 -17 1504
rect 17 1487 25 1504
rect -48 1462 -31 1470
rect -48 966 -31 974
rect 31 1462 48 1470
rect 31 966 48 974
rect -25 932 -17 949
rect 17 932 25 949
rect -25 878 -17 895
rect 17 878 25 895
rect -48 853 -31 861
rect -48 357 -31 365
rect 31 853 48 861
rect 31 357 48 365
rect -25 323 -17 340
rect 17 323 25 340
rect -25 269 -17 286
rect 17 269 25 286
rect -48 244 -31 252
rect -48 -252 -31 -244
rect 31 244 48 252
rect 31 -252 48 -244
rect -25 -286 -17 -269
rect 17 -286 25 -269
rect -25 -340 -17 -323
rect 17 -340 25 -323
rect -48 -365 -31 -357
rect -48 -861 -31 -853
rect 31 -365 48 -357
rect 31 -861 48 -853
rect -25 -895 -17 -878
rect 17 -895 25 -878
rect -25 -949 -17 -932
rect 17 -949 25 -932
rect -48 -974 -31 -966
rect -48 -1470 -31 -1462
rect 31 -974 48 -966
rect 31 -1470 48 -1462
rect -25 -1504 -17 -1487
rect 17 -1504 25 -1487
rect -25 -1558 -17 -1541
rect 17 -1558 25 -1541
rect -48 -1583 -31 -1575
rect -48 -2079 -31 -2071
rect 31 -1583 48 -1575
rect 31 -2079 48 -2071
rect -25 -2113 -17 -2096
rect 17 -2113 25 -2096
rect -105 -2147 -88 -2116
rect 88 -2147 105 -2116
rect -105 -2164 -57 -2147
rect 57 -2164 105 -2147
<< viali >>
rect -17 2096 17 2113
rect -48 1583 -31 2071
rect 31 1583 48 2071
rect -17 1541 17 1558
rect -17 1487 17 1504
rect -48 974 -31 1462
rect 31 974 48 1462
rect -17 932 17 949
rect -17 878 17 895
rect -48 365 -31 853
rect 31 365 48 853
rect -17 323 17 340
rect -17 269 17 286
rect -48 -244 -31 244
rect 31 -244 48 244
rect -17 -286 17 -269
rect -17 -340 17 -323
rect -48 -853 -31 -365
rect 31 -853 48 -365
rect -17 -895 17 -878
rect -17 -949 17 -932
rect -48 -1462 -31 -974
rect 31 -1462 48 -974
rect -17 -1504 17 -1487
rect -17 -1558 17 -1541
rect -48 -2071 -31 -1583
rect 31 -2071 48 -1583
rect -17 -2113 17 -2096
<< metal1 >>
rect -23 2113 23 2116
rect -23 2096 -17 2113
rect 17 2096 23 2113
rect -23 2093 23 2096
rect -51 2071 -28 2077
rect -51 1583 -48 2071
rect -31 1583 -28 2071
rect -51 1577 -28 1583
rect 28 2071 51 2077
rect 28 1583 31 2071
rect 48 1583 51 2071
rect 28 1577 51 1583
rect -23 1558 23 1561
rect -23 1541 -17 1558
rect 17 1541 23 1558
rect -23 1538 23 1541
rect -23 1504 23 1507
rect -23 1487 -17 1504
rect 17 1487 23 1504
rect -23 1484 23 1487
rect -51 1462 -28 1468
rect -51 974 -48 1462
rect -31 974 -28 1462
rect -51 968 -28 974
rect 28 1462 51 1468
rect 28 974 31 1462
rect 48 974 51 1462
rect 28 968 51 974
rect -23 949 23 952
rect -23 932 -17 949
rect 17 932 23 949
rect -23 929 23 932
rect -23 895 23 898
rect -23 878 -17 895
rect 17 878 23 895
rect -23 875 23 878
rect -51 853 -28 859
rect -51 365 -48 853
rect -31 365 -28 853
rect -51 359 -28 365
rect 28 853 51 859
rect 28 365 31 853
rect 48 365 51 853
rect 28 359 51 365
rect -23 340 23 343
rect -23 323 -17 340
rect 17 323 23 340
rect -23 320 23 323
rect -23 286 23 289
rect -23 269 -17 286
rect 17 269 23 286
rect -23 266 23 269
rect -51 244 -28 250
rect -51 -244 -48 244
rect -31 -244 -28 244
rect -51 -250 -28 -244
rect 28 244 51 250
rect 28 -244 31 244
rect 48 -244 51 244
rect 28 -250 51 -244
rect -23 -269 23 -266
rect -23 -286 -17 -269
rect 17 -286 23 -269
rect -23 -289 23 -286
rect -23 -323 23 -320
rect -23 -340 -17 -323
rect 17 -340 23 -323
rect -23 -343 23 -340
rect -51 -365 -28 -359
rect -51 -853 -48 -365
rect -31 -853 -28 -365
rect -51 -859 -28 -853
rect 28 -365 51 -359
rect 28 -853 31 -365
rect 48 -853 51 -365
rect 28 -859 51 -853
rect -23 -878 23 -875
rect -23 -895 -17 -878
rect 17 -895 23 -878
rect -23 -898 23 -895
rect -23 -932 23 -929
rect -23 -949 -17 -932
rect 17 -949 23 -932
rect -23 -952 23 -949
rect -51 -974 -28 -968
rect -51 -1462 -48 -974
rect -31 -1462 -28 -974
rect -51 -1468 -28 -1462
rect 28 -974 51 -968
rect 28 -1462 31 -974
rect 48 -1462 51 -974
rect 28 -1468 51 -1462
rect -23 -1487 23 -1484
rect -23 -1504 -17 -1487
rect 17 -1504 23 -1487
rect -23 -1507 23 -1504
rect -23 -1541 23 -1538
rect -23 -1558 -17 -1541
rect 17 -1558 23 -1541
rect -23 -1561 23 -1558
rect -51 -1583 -28 -1577
rect -51 -2071 -48 -1583
rect -31 -2071 -28 -1583
rect -51 -2077 -28 -2071
rect 28 -1583 51 -1577
rect 28 -2071 31 -1583
rect 48 -2071 51 -1583
rect 28 -2077 51 -2071
rect -23 -2096 23 -2093
rect -23 -2113 -17 -2096
rect 17 -2113 23 -2096
rect -23 -2116 23 -2113
<< properties >>
string FIXED_BBOX -96 -2155 96 2155
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.5 m 7 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
