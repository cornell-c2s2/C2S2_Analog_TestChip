magic
tech sky130A
magscale 1 2
timestamp 1679690840
<< pwell >>
rect -739 -1598 739 1598
<< psubdiff >>
rect -703 1528 -607 1562
rect 607 1528 703 1562
rect -703 1466 -669 1528
rect 669 1466 703 1528
rect -703 -1528 -669 -1466
rect 669 -1528 703 -1466
rect -703 -1562 -607 -1528
rect 607 -1562 703 -1528
<< psubdiffcont >>
rect -607 1528 607 1562
rect -703 -1466 -669 1466
rect 669 -1466 703 1466
rect -607 -1562 607 -1528
<< xpolycontact >>
rect -573 1000 573 1432
rect -573 -1432 573 -1000
<< xpolyres >>
rect -573 -1000 573 1000
<< locali >>
rect -703 1528 -607 1562
rect 607 1528 703 1562
rect -703 1466 -669 1528
rect 669 1466 703 1528
rect -703 -1528 -669 -1466
rect 669 -1528 703 -1466
rect -703 -1562 -607 -1528
rect 607 -1562 703 -1528
<< viali >>
rect -557 1017 557 1414
rect -557 -1414 557 -1017
<< metal1 >>
rect -569 1414 569 1420
rect -569 1017 -557 1414
rect 557 1017 569 1414
rect -569 1011 569 1017
rect -569 -1017 569 -1011
rect -569 -1414 -557 -1017
rect 557 -1414 569 -1017
rect -569 -1420 569 -1414
<< res5p73 >>
rect -575 -1002 575 1002
<< properties >>
string FIXED_BBOX -686 -1545 686 1545
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 10 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 3.556k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
