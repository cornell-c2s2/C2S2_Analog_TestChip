magic
tech sky130A
timestamp 1676134575
<< pwell >>
rect -148 -2182 148 2182
<< nmos >>
rect -50 1577 50 2077
rect -50 968 50 1468
rect -50 359 50 859
rect -50 -250 50 250
rect -50 -859 50 -359
rect -50 -1468 50 -968
rect -50 -2077 50 -1577
<< ndiff >>
rect -79 2071 -50 2077
rect -79 1583 -73 2071
rect -56 1583 -50 2071
rect -79 1577 -50 1583
rect 50 2071 79 2077
rect 50 1583 56 2071
rect 73 1583 79 2071
rect 50 1577 79 1583
rect -79 1462 -50 1468
rect -79 974 -73 1462
rect -56 974 -50 1462
rect -79 968 -50 974
rect 50 1462 79 1468
rect 50 974 56 1462
rect 73 974 79 1462
rect 50 968 79 974
rect -79 853 -50 859
rect -79 365 -73 853
rect -56 365 -50 853
rect -79 359 -50 365
rect 50 853 79 859
rect 50 365 56 853
rect 73 365 79 853
rect 50 359 79 365
rect -79 244 -50 250
rect -79 -244 -73 244
rect -56 -244 -50 244
rect -79 -250 -50 -244
rect 50 244 79 250
rect 50 -244 56 244
rect 73 -244 79 244
rect 50 -250 79 -244
rect -79 -365 -50 -359
rect -79 -853 -73 -365
rect -56 -853 -50 -365
rect -79 -859 -50 -853
rect 50 -365 79 -359
rect 50 -853 56 -365
rect 73 -853 79 -365
rect 50 -859 79 -853
rect -79 -974 -50 -968
rect -79 -1462 -73 -974
rect -56 -1462 -50 -974
rect -79 -1468 -50 -1462
rect 50 -974 79 -968
rect 50 -1462 56 -974
rect 73 -1462 79 -974
rect 50 -1468 79 -1462
rect -79 -1583 -50 -1577
rect -79 -2071 -73 -1583
rect -56 -2071 -50 -1583
rect -79 -2077 -50 -2071
rect 50 -1583 79 -1577
rect 50 -2071 56 -1583
rect 73 -2071 79 -1583
rect 50 -2077 79 -2071
<< ndiffc >>
rect -73 1583 -56 2071
rect 56 1583 73 2071
rect -73 974 -56 1462
rect 56 974 73 1462
rect -73 365 -56 853
rect 56 365 73 853
rect -73 -244 -56 244
rect 56 -244 73 244
rect -73 -853 -56 -365
rect 56 -853 73 -365
rect -73 -1462 -56 -974
rect 56 -1462 73 -974
rect -73 -2071 -56 -1583
rect 56 -2071 73 -1583
<< psubdiff >>
rect -130 2147 -82 2164
rect 82 2147 130 2164
rect -130 2116 -113 2147
rect 113 2116 130 2147
rect -130 -2147 -113 -2116
rect 113 -2147 130 -2116
rect -130 -2164 -82 -2147
rect 82 -2164 130 -2147
<< psubdiffcont >>
rect -82 2147 82 2164
rect -130 -2116 -113 2116
rect 113 -2116 130 2116
rect -82 -2164 82 -2147
<< poly >>
rect -50 2113 50 2121
rect -50 2096 -42 2113
rect 42 2096 50 2113
rect -50 2077 50 2096
rect -50 1558 50 1577
rect -50 1541 -42 1558
rect 42 1541 50 1558
rect -50 1533 50 1541
rect -50 1504 50 1512
rect -50 1487 -42 1504
rect 42 1487 50 1504
rect -50 1468 50 1487
rect -50 949 50 968
rect -50 932 -42 949
rect 42 932 50 949
rect -50 924 50 932
rect -50 895 50 903
rect -50 878 -42 895
rect 42 878 50 895
rect -50 859 50 878
rect -50 340 50 359
rect -50 323 -42 340
rect 42 323 50 340
rect -50 315 50 323
rect -50 286 50 294
rect -50 269 -42 286
rect 42 269 50 286
rect -50 250 50 269
rect -50 -269 50 -250
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -50 -294 50 -286
rect -50 -323 50 -315
rect -50 -340 -42 -323
rect 42 -340 50 -323
rect -50 -359 50 -340
rect -50 -878 50 -859
rect -50 -895 -42 -878
rect 42 -895 50 -878
rect -50 -903 50 -895
rect -50 -932 50 -924
rect -50 -949 -42 -932
rect 42 -949 50 -932
rect -50 -968 50 -949
rect -50 -1487 50 -1468
rect -50 -1504 -42 -1487
rect 42 -1504 50 -1487
rect -50 -1512 50 -1504
rect -50 -1541 50 -1533
rect -50 -1558 -42 -1541
rect 42 -1558 50 -1541
rect -50 -1577 50 -1558
rect -50 -2096 50 -2077
rect -50 -2113 -42 -2096
rect 42 -2113 50 -2096
rect -50 -2121 50 -2113
<< polycont >>
rect -42 2096 42 2113
rect -42 1541 42 1558
rect -42 1487 42 1504
rect -42 932 42 949
rect -42 878 42 895
rect -42 323 42 340
rect -42 269 42 286
rect -42 -286 42 -269
rect -42 -340 42 -323
rect -42 -895 42 -878
rect -42 -949 42 -932
rect -42 -1504 42 -1487
rect -42 -1558 42 -1541
rect -42 -2113 42 -2096
<< locali >>
rect -130 2147 -82 2164
rect 82 2147 130 2164
rect -130 2116 -113 2147
rect 113 2116 130 2147
rect -50 2096 -42 2113
rect 42 2096 50 2113
rect -73 2071 -56 2079
rect -73 1575 -56 1583
rect 56 2071 73 2079
rect 56 1575 73 1583
rect -50 1541 -42 1558
rect 42 1541 50 1558
rect -50 1487 -42 1504
rect 42 1487 50 1504
rect -73 1462 -56 1470
rect -73 966 -56 974
rect 56 1462 73 1470
rect 56 966 73 974
rect -50 932 -42 949
rect 42 932 50 949
rect -50 878 -42 895
rect 42 878 50 895
rect -73 853 -56 861
rect -73 357 -56 365
rect 56 853 73 861
rect 56 357 73 365
rect -50 323 -42 340
rect 42 323 50 340
rect -50 269 -42 286
rect 42 269 50 286
rect -73 244 -56 252
rect -73 -252 -56 -244
rect 56 244 73 252
rect 56 -252 73 -244
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -50 -340 -42 -323
rect 42 -340 50 -323
rect -73 -365 -56 -357
rect -73 -861 -56 -853
rect 56 -365 73 -357
rect 56 -861 73 -853
rect -50 -895 -42 -878
rect 42 -895 50 -878
rect -50 -949 -42 -932
rect 42 -949 50 -932
rect -73 -974 -56 -966
rect -73 -1470 -56 -1462
rect 56 -974 73 -966
rect 56 -1470 73 -1462
rect -50 -1504 -42 -1487
rect 42 -1504 50 -1487
rect -50 -1558 -42 -1541
rect 42 -1558 50 -1541
rect -73 -1583 -56 -1575
rect -73 -2079 -56 -2071
rect 56 -1583 73 -1575
rect 56 -2079 73 -2071
rect -50 -2113 -42 -2096
rect 42 -2113 50 -2096
rect -130 -2147 -113 -2116
rect 113 -2147 130 -2116
rect -130 -2164 -82 -2147
rect 82 -2164 130 -2147
<< viali >>
rect -42 2096 42 2113
rect -73 1583 -56 2071
rect 56 1583 73 2071
rect -42 1541 42 1558
rect -42 1487 42 1504
rect -73 974 -56 1462
rect 56 974 73 1462
rect -42 932 42 949
rect -42 878 42 895
rect -73 365 -56 853
rect 56 365 73 853
rect -42 323 42 340
rect -42 269 42 286
rect -73 -244 -56 244
rect 56 -244 73 244
rect -42 -286 42 -269
rect -42 -340 42 -323
rect -73 -853 -56 -365
rect 56 -853 73 -365
rect -42 -895 42 -878
rect -42 -949 42 -932
rect -73 -1462 -56 -974
rect 56 -1462 73 -974
rect -42 -1504 42 -1487
rect -42 -1558 42 -1541
rect -73 -2071 -56 -1583
rect 56 -2071 73 -1583
rect -42 -2113 42 -2096
<< metal1 >>
rect -48 2113 48 2116
rect -48 2096 -42 2113
rect 42 2096 48 2113
rect -48 2093 48 2096
rect -76 2071 -53 2077
rect -76 1583 -73 2071
rect -56 1583 -53 2071
rect -76 1577 -53 1583
rect 53 2071 76 2077
rect 53 1583 56 2071
rect 73 1583 76 2071
rect 53 1577 76 1583
rect -48 1558 48 1561
rect -48 1541 -42 1558
rect 42 1541 48 1558
rect -48 1538 48 1541
rect -48 1504 48 1507
rect -48 1487 -42 1504
rect 42 1487 48 1504
rect -48 1484 48 1487
rect -76 1462 -53 1468
rect -76 974 -73 1462
rect -56 974 -53 1462
rect -76 968 -53 974
rect 53 1462 76 1468
rect 53 974 56 1462
rect 73 974 76 1462
rect 53 968 76 974
rect -48 949 48 952
rect -48 932 -42 949
rect 42 932 48 949
rect -48 929 48 932
rect -48 895 48 898
rect -48 878 -42 895
rect 42 878 48 895
rect -48 875 48 878
rect -76 853 -53 859
rect -76 365 -73 853
rect -56 365 -53 853
rect -76 359 -53 365
rect 53 853 76 859
rect 53 365 56 853
rect 73 365 76 853
rect 53 359 76 365
rect -48 340 48 343
rect -48 323 -42 340
rect 42 323 48 340
rect -48 320 48 323
rect -48 286 48 289
rect -48 269 -42 286
rect 42 269 48 286
rect -48 266 48 269
rect -76 244 -53 250
rect -76 -244 -73 244
rect -56 -244 -53 244
rect -76 -250 -53 -244
rect 53 244 76 250
rect 53 -244 56 244
rect 73 -244 76 244
rect 53 -250 76 -244
rect -48 -269 48 -266
rect -48 -286 -42 -269
rect 42 -286 48 -269
rect -48 -289 48 -286
rect -48 -323 48 -320
rect -48 -340 -42 -323
rect 42 -340 48 -323
rect -48 -343 48 -340
rect -76 -365 -53 -359
rect -76 -853 -73 -365
rect -56 -853 -53 -365
rect -76 -859 -53 -853
rect 53 -365 76 -359
rect 53 -853 56 -365
rect 73 -853 76 -365
rect 53 -859 76 -853
rect -48 -878 48 -875
rect -48 -895 -42 -878
rect 42 -895 48 -878
rect -48 -898 48 -895
rect -48 -932 48 -929
rect -48 -949 -42 -932
rect 42 -949 48 -932
rect -48 -952 48 -949
rect -76 -974 -53 -968
rect -76 -1462 -73 -974
rect -56 -1462 -53 -974
rect -76 -1468 -53 -1462
rect 53 -974 76 -968
rect 53 -1462 56 -974
rect 73 -1462 76 -974
rect 53 -1468 76 -1462
rect -48 -1487 48 -1484
rect -48 -1504 -42 -1487
rect 42 -1504 48 -1487
rect -48 -1507 48 -1504
rect -48 -1541 48 -1538
rect -48 -1558 -42 -1541
rect 42 -1558 48 -1541
rect -48 -1561 48 -1558
rect -76 -1583 -53 -1577
rect -76 -2071 -73 -1583
rect -56 -2071 -53 -1583
rect -76 -2077 -53 -2071
rect 53 -1583 76 -1577
rect 53 -2071 56 -1583
rect 73 -2071 76 -1583
rect 53 -2077 76 -2071
rect -48 -2096 48 -2093
rect -48 -2113 -42 -2096
rect 42 -2113 48 -2096
rect -48 -2116 48 -2113
<< properties >>
string FIXED_BBOX -121 -2155 121 2155
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 1 m 7 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
