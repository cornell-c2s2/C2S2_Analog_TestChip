magic
tech sky130A
magscale 1 2
timestamp 1678919179
<< error_p >>
rect -3589 -1700 -3529 1700
rect -3509 -1700 -3449 1700
rect -70 -1700 -10 1700
rect 10 -1700 70 1700
rect 3449 -1700 3509 1700
rect 3529 -1700 3589 1700
<< metal3 >>
rect -7028 1672 -3529 1700
rect -7028 -1672 -3613 1672
rect -3549 -1672 -3529 1672
rect -7028 -1700 -3529 -1672
rect -3509 1672 -10 1700
rect -3509 -1672 -94 1672
rect -30 -1672 -10 1672
rect -3509 -1700 -10 -1672
rect 10 1672 3509 1700
rect 10 -1672 3425 1672
rect 3489 -1672 3509 1672
rect 10 -1700 3509 -1672
rect 3529 1672 7028 1700
rect 3529 -1672 6944 1672
rect 7008 -1672 7028 1672
rect 3529 -1700 7028 -1672
<< via3 >>
rect -3613 -1672 -3549 1672
rect -94 -1672 -30 1672
rect 3425 -1672 3489 1672
rect 6944 -1672 7008 1672
<< mimcap >>
rect -6928 1560 -3728 1600
rect -6928 -1560 -6888 1560
rect -3768 -1560 -3728 1560
rect -6928 -1600 -3728 -1560
rect -3409 1560 -209 1600
rect -3409 -1560 -3369 1560
rect -249 -1560 -209 1560
rect -3409 -1600 -209 -1560
rect 110 1560 3310 1600
rect 110 -1560 150 1560
rect 3270 -1560 3310 1560
rect 110 -1600 3310 -1560
rect 3629 1560 6829 1600
rect 3629 -1560 3669 1560
rect 6789 -1560 6829 1560
rect 3629 -1600 6829 -1560
<< mimcapcontact >>
rect -6888 -1560 -3768 1560
rect -3369 -1560 -249 1560
rect 150 -1560 3270 1560
rect 3669 -1560 6789 1560
<< metal4 >>
rect -3629 1672 -3533 1688
rect -6889 1560 -3767 1561
rect -6889 -1560 -6888 1560
rect -3768 -1560 -3767 1560
rect -6889 -1561 -3767 -1560
rect -3629 -1672 -3613 1672
rect -3549 -1672 -3533 1672
rect -110 1672 -14 1688
rect -3370 1560 -248 1561
rect -3370 -1560 -3369 1560
rect -249 -1560 -248 1560
rect -3370 -1561 -248 -1560
rect -3629 -1688 -3533 -1672
rect -110 -1672 -94 1672
rect -30 -1672 -14 1672
rect 3409 1672 3505 1688
rect 149 1560 3271 1561
rect 149 -1560 150 1560
rect 3270 -1560 3271 1560
rect 149 -1561 3271 -1560
rect -110 -1688 -14 -1672
rect 3409 -1672 3425 1672
rect 3489 -1672 3505 1672
rect 6928 1672 7024 1688
rect 3668 1560 6790 1561
rect 3668 -1560 3669 1560
rect 6789 -1560 6790 1560
rect 3668 -1561 6790 -1560
rect 3409 -1688 3505 -1672
rect 6928 -1672 6944 1672
rect 7008 -1672 7024 1672
rect 6928 -1688 7024 -1672
<< properties >>
string FIXED_BBOX 3529 -1700 6929 1700
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 16 l 16 val 524.159 carea 2.00 cperi 0.19 nx 4 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
