magic
tech sky130A
magscale 1 2
timestamp 1683391037
<< pwell >>
rect -683 -335 683 335
<< nmos >>
rect -487 -125 -287 125
rect -229 -125 -29 125
rect 29 -125 229 125
rect 287 -125 487 125
<< ndiff >>
rect -545 113 -487 125
rect -545 -113 -533 113
rect -499 -113 -487 113
rect -545 -125 -487 -113
rect -287 113 -229 125
rect -287 -113 -275 113
rect -241 -113 -229 113
rect -287 -125 -229 -113
rect -29 113 29 125
rect -29 -113 -17 113
rect 17 -113 29 113
rect -29 -125 29 -113
rect 229 113 287 125
rect 229 -113 241 113
rect 275 -113 287 113
rect 229 -125 287 -113
rect 487 113 545 125
rect 487 -113 499 113
rect 533 -113 545 113
rect 487 -125 545 -113
<< ndiffc >>
rect -533 -113 -499 113
rect -275 -113 -241 113
rect -17 -113 17 113
rect 241 -113 275 113
rect 499 -113 533 113
<< psubdiff >>
rect -647 265 -551 299
rect 551 265 647 299
rect -647 203 -613 265
rect 613 203 647 265
rect -647 -265 -613 -203
rect 613 -265 647 -203
rect -647 -299 -551 -265
rect 551 -299 647 -265
<< psubdiffcont >>
rect -551 265 551 299
rect -647 -203 -613 203
rect 613 -203 647 203
rect -551 -299 551 -265
<< poly >>
rect -487 197 -287 213
rect -487 163 -471 197
rect -303 163 -287 197
rect -487 125 -287 163
rect -229 197 -29 213
rect -229 163 -213 197
rect -45 163 -29 197
rect -229 125 -29 163
rect 29 197 229 213
rect 29 163 45 197
rect 213 163 229 197
rect 29 125 229 163
rect 287 197 487 213
rect 287 163 303 197
rect 471 163 487 197
rect 287 125 487 163
rect -487 -163 -287 -125
rect -487 -197 -471 -163
rect -303 -197 -287 -163
rect -487 -213 -287 -197
rect -229 -163 -29 -125
rect -229 -197 -213 -163
rect -45 -197 -29 -163
rect -229 -213 -29 -197
rect 29 -163 229 -125
rect 29 -197 45 -163
rect 213 -197 229 -163
rect 29 -213 229 -197
rect 287 -163 487 -125
rect 287 -197 303 -163
rect 471 -197 487 -163
rect 287 -213 487 -197
<< polycont >>
rect -471 163 -303 197
rect -213 163 -45 197
rect 45 163 213 197
rect 303 163 471 197
rect -471 -197 -303 -163
rect -213 -197 -45 -163
rect 45 -197 213 -163
rect 303 -197 471 -163
<< locali >>
rect -647 265 -551 299
rect 551 265 647 299
rect -647 203 -613 265
rect 613 203 647 265
rect -487 163 -471 197
rect -303 163 -287 197
rect -229 163 -213 197
rect -45 163 -29 197
rect 29 163 45 197
rect 213 163 229 197
rect 287 163 303 197
rect 471 163 487 197
rect -533 113 -499 129
rect -533 -129 -499 -113
rect -275 113 -241 129
rect -275 -129 -241 -113
rect -17 113 17 129
rect -17 -129 17 -113
rect 241 113 275 129
rect 241 -129 275 -113
rect 499 113 533 129
rect 499 -129 533 -113
rect -487 -197 -471 -163
rect -303 -197 -287 -163
rect -229 -197 -213 -163
rect -45 -197 -29 -163
rect 29 -197 45 -163
rect 213 -197 229 -163
rect 287 -197 303 -163
rect 471 -197 487 -163
rect -647 -265 -613 -203
rect 613 -265 647 -203
rect -647 -299 -551 -265
rect 551 -299 647 -265
<< viali >>
rect -471 163 -303 197
rect -213 163 -45 197
rect 45 163 213 197
rect 303 163 471 197
rect -533 -113 -499 113
rect -275 -113 -241 113
rect -17 -113 17 113
rect 241 -113 275 113
rect 499 -113 533 113
rect -471 -197 -303 -163
rect -213 -197 -45 -163
rect 45 -197 213 -163
rect 303 -197 471 -163
<< metal1 >>
rect -483 197 -291 203
rect -483 163 -471 197
rect -303 163 -291 197
rect -483 157 -291 163
rect -225 197 -33 203
rect -225 163 -213 197
rect -45 163 -33 197
rect -225 157 -33 163
rect 33 197 225 203
rect 33 163 45 197
rect 213 163 225 197
rect 33 157 225 163
rect 291 197 483 203
rect 291 163 303 197
rect 471 163 483 197
rect 291 157 483 163
rect -539 113 -493 125
rect -539 -113 -533 113
rect -499 -113 -493 113
rect -539 -125 -493 -113
rect -281 113 -235 125
rect -281 -113 -275 113
rect -241 -113 -235 113
rect -281 -125 -235 -113
rect -23 113 23 125
rect -23 -113 -17 113
rect 17 -113 23 113
rect -23 -125 23 -113
rect 235 113 281 125
rect 235 -113 241 113
rect 275 -113 281 113
rect 235 -125 281 -113
rect 493 113 539 125
rect 493 -113 499 113
rect 533 -113 539 113
rect 493 -125 539 -113
rect -483 -163 -291 -157
rect -483 -197 -471 -163
rect -303 -197 -291 -163
rect -483 -203 -291 -197
rect -225 -163 -33 -157
rect -225 -197 -213 -163
rect -45 -197 -33 -163
rect -225 -203 -33 -197
rect 33 -163 225 -157
rect 33 -197 45 -163
rect 213 -197 225 -163
rect 33 -203 225 -197
rect 291 -163 483 -157
rect 291 -197 303 -163
rect 471 -197 483 -163
rect 291 -203 483 -197
<< properties >>
string FIXED_BBOX -630 -282 630 282
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.25 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
