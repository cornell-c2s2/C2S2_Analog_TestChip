magic
tech sky130A
timestamp 1676129039
<< pwell >>
rect -148 -964 148 964
<< nmos >>
rect -50 359 50 859
rect -50 -250 50 250
rect -50 -859 50 -359
<< ndiff >>
rect -79 853 -50 859
rect -79 365 -73 853
rect -56 365 -50 853
rect -79 359 -50 365
rect 50 853 79 859
rect 50 365 56 853
rect 73 365 79 853
rect 50 359 79 365
rect -79 244 -50 250
rect -79 -244 -73 244
rect -56 -244 -50 244
rect -79 -250 -50 -244
rect 50 244 79 250
rect 50 -244 56 244
rect 73 -244 79 244
rect 50 -250 79 -244
rect -79 -365 -50 -359
rect -79 -853 -73 -365
rect -56 -853 -50 -365
rect -79 -859 -50 -853
rect 50 -365 79 -359
rect 50 -853 56 -365
rect 73 -853 79 -365
rect 50 -859 79 -853
<< ndiffc >>
rect -73 365 -56 853
rect 56 365 73 853
rect -73 -244 -56 244
rect 56 -244 73 244
rect -73 -853 -56 -365
rect 56 -853 73 -365
<< psubdiff >>
rect -130 929 -82 946
rect 82 929 130 946
rect -130 898 -113 929
rect 113 898 130 929
rect -130 -929 -113 -898
rect 113 -929 130 -898
rect -130 -946 -82 -929
rect 82 -946 130 -929
<< psubdiffcont >>
rect -82 929 82 946
rect -130 -898 -113 898
rect 113 -898 130 898
rect -82 -946 82 -929
<< poly >>
rect -50 895 50 903
rect -50 878 -42 895
rect 42 878 50 895
rect -50 859 50 878
rect -50 340 50 359
rect -50 323 -42 340
rect 42 323 50 340
rect -50 315 50 323
rect -50 286 50 294
rect -50 269 -42 286
rect 42 269 50 286
rect -50 250 50 269
rect -50 -269 50 -250
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -50 -294 50 -286
rect -50 -323 50 -315
rect -50 -340 -42 -323
rect 42 -340 50 -323
rect -50 -359 50 -340
rect -50 -878 50 -859
rect -50 -895 -42 -878
rect 42 -895 50 -878
rect -50 -903 50 -895
<< polycont >>
rect -42 878 42 895
rect -42 323 42 340
rect -42 269 42 286
rect -42 -286 42 -269
rect -42 -340 42 -323
rect -42 -895 42 -878
<< locali >>
rect -130 929 -82 946
rect 82 929 130 946
rect -130 898 -113 929
rect 113 898 130 929
rect -50 878 -42 895
rect 42 878 50 895
rect -73 853 -56 861
rect -73 357 -56 365
rect 56 853 73 861
rect 56 357 73 365
rect -50 323 -42 340
rect 42 323 50 340
rect -50 269 -42 286
rect 42 269 50 286
rect -73 244 -56 252
rect -73 -252 -56 -244
rect 56 244 73 252
rect 56 -252 73 -244
rect -50 -286 -42 -269
rect 42 -286 50 -269
rect -50 -340 -42 -323
rect 42 -340 50 -323
rect -73 -365 -56 -357
rect -73 -861 -56 -853
rect 56 -365 73 -357
rect 56 -861 73 -853
rect -50 -895 -42 -878
rect 42 -895 50 -878
rect -130 -929 -113 -898
rect 113 -929 130 -898
rect -130 -946 -82 -929
rect 82 -946 130 -929
<< viali >>
rect -42 878 42 895
rect -73 365 -56 853
rect 56 365 73 853
rect -42 323 42 340
rect -42 269 42 286
rect -73 -244 -56 244
rect 56 -244 73 244
rect -42 -286 42 -269
rect -42 -340 42 -323
rect -73 -853 -56 -365
rect 56 -853 73 -365
rect -42 -895 42 -878
<< metal1 >>
rect -48 895 48 898
rect -48 878 -42 895
rect 42 878 48 895
rect -48 875 48 878
rect -76 853 -53 859
rect -76 365 -73 853
rect -56 365 -53 853
rect -76 359 -53 365
rect 53 853 76 859
rect 53 365 56 853
rect 73 365 76 853
rect 53 359 76 365
rect -48 340 48 343
rect -48 323 -42 340
rect 42 323 48 340
rect -48 320 48 323
rect -48 286 48 289
rect -48 269 -42 286
rect 42 269 48 286
rect -48 266 48 269
rect -76 244 -53 250
rect -76 -244 -73 244
rect -56 -244 -53 244
rect -76 -250 -53 -244
rect 53 244 76 250
rect 53 -244 56 244
rect 73 -244 76 244
rect 53 -250 76 -244
rect -48 -269 48 -266
rect -48 -286 -42 -269
rect 42 -286 48 -269
rect -48 -289 48 -286
rect -48 -323 48 -320
rect -48 -340 -42 -323
rect 42 -340 48 -323
rect -48 -343 48 -340
rect -76 -365 -53 -359
rect -76 -853 -73 -365
rect -56 -853 -53 -365
rect -76 -859 -53 -853
rect 53 -365 76 -359
rect 53 -853 56 -365
rect 73 -853 76 -365
rect 53 -859 76 -853
rect -48 -878 48 -875
rect -48 -895 -42 -878
rect 42 -895 48 -878
rect -48 -898 48 -895
<< properties >>
string FIXED_BBOX -121 -937 121 937
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 1 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
