magic
tech sky130A
magscale 1 2
timestamp 1676739250
<< pwell >>
rect -5436 3002 5436 3088
rect -5436 -3002 -5350 3002
rect 5350 -3002 5436 3002
rect -5436 -3088 5436 -3002
<< psubdiff >>
rect -5410 3028 -5287 3062
rect -5253 3028 -5219 3062
rect -5185 3028 -5151 3062
rect -5117 3028 -5083 3062
rect -5049 3028 -5015 3062
rect -4981 3028 -4947 3062
rect -4913 3028 -4879 3062
rect -4845 3028 -4811 3062
rect -4777 3028 -4743 3062
rect -4709 3028 -4675 3062
rect -4641 3028 -4607 3062
rect -4573 3028 -4539 3062
rect -4505 3028 -4471 3062
rect -4437 3028 -4403 3062
rect -4369 3028 -4335 3062
rect -4301 3028 -4267 3062
rect -4233 3028 -4199 3062
rect -4165 3028 -4131 3062
rect -4097 3028 -4063 3062
rect -4029 3028 -3995 3062
rect -3961 3028 -3927 3062
rect -3893 3028 -3859 3062
rect -3825 3028 -3791 3062
rect -3757 3028 -3723 3062
rect -3689 3028 -3655 3062
rect -3621 3028 -3587 3062
rect -3553 3028 -3519 3062
rect -3485 3028 -3451 3062
rect -3417 3028 -3383 3062
rect -3349 3028 -3315 3062
rect -3281 3028 -3247 3062
rect -3213 3028 -3179 3062
rect -3145 3028 -3111 3062
rect -3077 3028 -3043 3062
rect -3009 3028 -2975 3062
rect -2941 3028 -2907 3062
rect -2873 3028 -2839 3062
rect -2805 3028 -2771 3062
rect -2737 3028 -2703 3062
rect -2669 3028 -2635 3062
rect -2601 3028 -2567 3062
rect -2533 3028 -2499 3062
rect -2465 3028 -2431 3062
rect -2397 3028 -2363 3062
rect -2329 3028 -2295 3062
rect -2261 3028 -2227 3062
rect -2193 3028 -2159 3062
rect -2125 3028 -2091 3062
rect -2057 3028 -2023 3062
rect -1989 3028 -1955 3062
rect -1921 3028 -1887 3062
rect -1853 3028 -1819 3062
rect -1785 3028 -1751 3062
rect -1717 3028 -1683 3062
rect -1649 3028 -1615 3062
rect -1581 3028 -1547 3062
rect -1513 3028 -1479 3062
rect -1445 3028 -1411 3062
rect -1377 3028 -1343 3062
rect -1309 3028 -1275 3062
rect -1241 3028 -1207 3062
rect -1173 3028 -1139 3062
rect -1105 3028 -1071 3062
rect -1037 3028 -1003 3062
rect -969 3028 -935 3062
rect -901 3028 -867 3062
rect -833 3028 -799 3062
rect -765 3028 -731 3062
rect -697 3028 -663 3062
rect -629 3028 -595 3062
rect -561 3028 -527 3062
rect -493 3028 -459 3062
rect -425 3028 -391 3062
rect -357 3028 -323 3062
rect -289 3028 -255 3062
rect -221 3028 -187 3062
rect -153 3028 -119 3062
rect -85 3028 -51 3062
rect -17 3028 17 3062
rect 51 3028 85 3062
rect 119 3028 153 3062
rect 187 3028 221 3062
rect 255 3028 289 3062
rect 323 3028 357 3062
rect 391 3028 425 3062
rect 459 3028 493 3062
rect 527 3028 561 3062
rect 595 3028 629 3062
rect 663 3028 697 3062
rect 731 3028 765 3062
rect 799 3028 833 3062
rect 867 3028 901 3062
rect 935 3028 969 3062
rect 1003 3028 1037 3062
rect 1071 3028 1105 3062
rect 1139 3028 1173 3062
rect 1207 3028 1241 3062
rect 1275 3028 1309 3062
rect 1343 3028 1377 3062
rect 1411 3028 1445 3062
rect 1479 3028 1513 3062
rect 1547 3028 1581 3062
rect 1615 3028 1649 3062
rect 1683 3028 1717 3062
rect 1751 3028 1785 3062
rect 1819 3028 1853 3062
rect 1887 3028 1921 3062
rect 1955 3028 1989 3062
rect 2023 3028 2057 3062
rect 2091 3028 2125 3062
rect 2159 3028 2193 3062
rect 2227 3028 2261 3062
rect 2295 3028 2329 3062
rect 2363 3028 2397 3062
rect 2431 3028 2465 3062
rect 2499 3028 2533 3062
rect 2567 3028 2601 3062
rect 2635 3028 2669 3062
rect 2703 3028 2737 3062
rect 2771 3028 2805 3062
rect 2839 3028 2873 3062
rect 2907 3028 2941 3062
rect 2975 3028 3009 3062
rect 3043 3028 3077 3062
rect 3111 3028 3145 3062
rect 3179 3028 3213 3062
rect 3247 3028 3281 3062
rect 3315 3028 3349 3062
rect 3383 3028 3417 3062
rect 3451 3028 3485 3062
rect 3519 3028 3553 3062
rect 3587 3028 3621 3062
rect 3655 3028 3689 3062
rect 3723 3028 3757 3062
rect 3791 3028 3825 3062
rect 3859 3028 3893 3062
rect 3927 3028 3961 3062
rect 3995 3028 4029 3062
rect 4063 3028 4097 3062
rect 4131 3028 4165 3062
rect 4199 3028 4233 3062
rect 4267 3028 4301 3062
rect 4335 3028 4369 3062
rect 4403 3028 4437 3062
rect 4471 3028 4505 3062
rect 4539 3028 4573 3062
rect 4607 3028 4641 3062
rect 4675 3028 4709 3062
rect 4743 3028 4777 3062
rect 4811 3028 4845 3062
rect 4879 3028 4913 3062
rect 4947 3028 4981 3062
rect 5015 3028 5049 3062
rect 5083 3028 5117 3062
rect 5151 3028 5185 3062
rect 5219 3028 5253 3062
rect 5287 3028 5410 3062
rect -5410 2941 -5376 3028
rect 5376 2941 5410 3028
rect -5410 2873 -5376 2907
rect -5410 2805 -5376 2839
rect -5410 2737 -5376 2771
rect -5410 2669 -5376 2703
rect -5410 2601 -5376 2635
rect -5410 2533 -5376 2567
rect -5410 2465 -5376 2499
rect -5410 2397 -5376 2431
rect -5410 2329 -5376 2363
rect -5410 2261 -5376 2295
rect -5410 2193 -5376 2227
rect -5410 2125 -5376 2159
rect -5410 2057 -5376 2091
rect -5410 1989 -5376 2023
rect -5410 1921 -5376 1955
rect -5410 1853 -5376 1887
rect -5410 1785 -5376 1819
rect -5410 1717 -5376 1751
rect -5410 1649 -5376 1683
rect -5410 1581 -5376 1615
rect -5410 1513 -5376 1547
rect -5410 1445 -5376 1479
rect -5410 1377 -5376 1411
rect -5410 1309 -5376 1343
rect -5410 1241 -5376 1275
rect -5410 1173 -5376 1207
rect -5410 1105 -5376 1139
rect -5410 1037 -5376 1071
rect -5410 969 -5376 1003
rect -5410 901 -5376 935
rect -5410 833 -5376 867
rect -5410 765 -5376 799
rect -5410 697 -5376 731
rect -5410 629 -5376 663
rect -5410 561 -5376 595
rect -5410 493 -5376 527
rect -5410 425 -5376 459
rect -5410 357 -5376 391
rect -5410 289 -5376 323
rect -5410 221 -5376 255
rect -5410 153 -5376 187
rect -5410 85 -5376 119
rect -5410 17 -5376 51
rect -5410 -51 -5376 -17
rect -5410 -119 -5376 -85
rect -5410 -187 -5376 -153
rect -5410 -255 -5376 -221
rect -5410 -323 -5376 -289
rect -5410 -391 -5376 -357
rect -5410 -459 -5376 -425
rect -5410 -527 -5376 -493
rect -5410 -595 -5376 -561
rect -5410 -663 -5376 -629
rect -5410 -731 -5376 -697
rect -5410 -799 -5376 -765
rect -5410 -867 -5376 -833
rect -5410 -935 -5376 -901
rect -5410 -1003 -5376 -969
rect -5410 -1071 -5376 -1037
rect -5410 -1139 -5376 -1105
rect -5410 -1207 -5376 -1173
rect -5410 -1275 -5376 -1241
rect -5410 -1343 -5376 -1309
rect -5410 -1411 -5376 -1377
rect -5410 -1479 -5376 -1445
rect -5410 -1547 -5376 -1513
rect -5410 -1615 -5376 -1581
rect -5410 -1683 -5376 -1649
rect -5410 -1751 -5376 -1717
rect -5410 -1819 -5376 -1785
rect -5410 -1887 -5376 -1853
rect -5410 -1955 -5376 -1921
rect -5410 -2023 -5376 -1989
rect -5410 -2091 -5376 -2057
rect -5410 -2159 -5376 -2125
rect -5410 -2227 -5376 -2193
rect -5410 -2295 -5376 -2261
rect -5410 -2363 -5376 -2329
rect -5410 -2431 -5376 -2397
rect -5410 -2499 -5376 -2465
rect -5410 -2567 -5376 -2533
rect -5410 -2635 -5376 -2601
rect -5410 -2703 -5376 -2669
rect -5410 -2771 -5376 -2737
rect -5410 -2839 -5376 -2805
rect -5410 -2907 -5376 -2873
rect 5376 2873 5410 2907
rect 5376 2805 5410 2839
rect 5376 2737 5410 2771
rect 5376 2669 5410 2703
rect 5376 2601 5410 2635
rect 5376 2533 5410 2567
rect 5376 2465 5410 2499
rect 5376 2397 5410 2431
rect 5376 2329 5410 2363
rect 5376 2261 5410 2295
rect 5376 2193 5410 2227
rect 5376 2125 5410 2159
rect 5376 2057 5410 2091
rect 5376 1989 5410 2023
rect 5376 1921 5410 1955
rect 5376 1853 5410 1887
rect 5376 1785 5410 1819
rect 5376 1717 5410 1751
rect 5376 1649 5410 1683
rect 5376 1581 5410 1615
rect 5376 1513 5410 1547
rect 5376 1445 5410 1479
rect 5376 1377 5410 1411
rect 5376 1309 5410 1343
rect 5376 1241 5410 1275
rect 5376 1173 5410 1207
rect 5376 1105 5410 1139
rect 5376 1037 5410 1071
rect 5376 969 5410 1003
rect 5376 901 5410 935
rect 5376 833 5410 867
rect 5376 765 5410 799
rect 5376 697 5410 731
rect 5376 629 5410 663
rect 5376 561 5410 595
rect 5376 493 5410 527
rect 5376 425 5410 459
rect 5376 357 5410 391
rect 5376 289 5410 323
rect 5376 221 5410 255
rect 5376 153 5410 187
rect 5376 85 5410 119
rect 5376 17 5410 51
rect 5376 -51 5410 -17
rect 5376 -119 5410 -85
rect 5376 -187 5410 -153
rect 5376 -255 5410 -221
rect 5376 -323 5410 -289
rect 5376 -391 5410 -357
rect 5376 -459 5410 -425
rect 5376 -527 5410 -493
rect 5376 -595 5410 -561
rect 5376 -663 5410 -629
rect 5376 -731 5410 -697
rect 5376 -799 5410 -765
rect 5376 -867 5410 -833
rect 5376 -935 5410 -901
rect 5376 -1003 5410 -969
rect 5376 -1071 5410 -1037
rect 5376 -1139 5410 -1105
rect 5376 -1207 5410 -1173
rect 5376 -1275 5410 -1241
rect 5376 -1343 5410 -1309
rect 5376 -1411 5410 -1377
rect 5376 -1479 5410 -1445
rect 5376 -1547 5410 -1513
rect 5376 -1615 5410 -1581
rect 5376 -1683 5410 -1649
rect 5376 -1751 5410 -1717
rect 5376 -1819 5410 -1785
rect 5376 -1887 5410 -1853
rect 5376 -1955 5410 -1921
rect 5376 -2023 5410 -1989
rect 5376 -2091 5410 -2057
rect 5376 -2159 5410 -2125
rect 5376 -2227 5410 -2193
rect 5376 -2295 5410 -2261
rect 5376 -2363 5410 -2329
rect 5376 -2431 5410 -2397
rect 5376 -2499 5410 -2465
rect 5376 -2567 5410 -2533
rect 5376 -2635 5410 -2601
rect 5376 -2703 5410 -2669
rect 5376 -2771 5410 -2737
rect 5376 -2839 5410 -2805
rect 5376 -2907 5410 -2873
rect -5410 -3028 -5376 -2941
rect 5376 -3028 5410 -2941
rect -5410 -3062 -5287 -3028
rect -5253 -3062 -5219 -3028
rect -5185 -3062 -5151 -3028
rect -5117 -3062 -5083 -3028
rect -5049 -3062 -5015 -3028
rect -4981 -3062 -4947 -3028
rect -4913 -3062 -4879 -3028
rect -4845 -3062 -4811 -3028
rect -4777 -3062 -4743 -3028
rect -4709 -3062 -4675 -3028
rect -4641 -3062 -4607 -3028
rect -4573 -3062 -4539 -3028
rect -4505 -3062 -4471 -3028
rect -4437 -3062 -4403 -3028
rect -4369 -3062 -4335 -3028
rect -4301 -3062 -4267 -3028
rect -4233 -3062 -4199 -3028
rect -4165 -3062 -4131 -3028
rect -4097 -3062 -4063 -3028
rect -4029 -3062 -3995 -3028
rect -3961 -3062 -3927 -3028
rect -3893 -3062 -3859 -3028
rect -3825 -3062 -3791 -3028
rect -3757 -3062 -3723 -3028
rect -3689 -3062 -3655 -3028
rect -3621 -3062 -3587 -3028
rect -3553 -3062 -3519 -3028
rect -3485 -3062 -3451 -3028
rect -3417 -3062 -3383 -3028
rect -3349 -3062 -3315 -3028
rect -3281 -3062 -3247 -3028
rect -3213 -3062 -3179 -3028
rect -3145 -3062 -3111 -3028
rect -3077 -3062 -3043 -3028
rect -3009 -3062 -2975 -3028
rect -2941 -3062 -2907 -3028
rect -2873 -3062 -2839 -3028
rect -2805 -3062 -2771 -3028
rect -2737 -3062 -2703 -3028
rect -2669 -3062 -2635 -3028
rect -2601 -3062 -2567 -3028
rect -2533 -3062 -2499 -3028
rect -2465 -3062 -2431 -3028
rect -2397 -3062 -2363 -3028
rect -2329 -3062 -2295 -3028
rect -2261 -3062 -2227 -3028
rect -2193 -3062 -2159 -3028
rect -2125 -3062 -2091 -3028
rect -2057 -3062 -2023 -3028
rect -1989 -3062 -1955 -3028
rect -1921 -3062 -1887 -3028
rect -1853 -3062 -1819 -3028
rect -1785 -3062 -1751 -3028
rect -1717 -3062 -1683 -3028
rect -1649 -3062 -1615 -3028
rect -1581 -3062 -1547 -3028
rect -1513 -3062 -1479 -3028
rect -1445 -3062 -1411 -3028
rect -1377 -3062 -1343 -3028
rect -1309 -3062 -1275 -3028
rect -1241 -3062 -1207 -3028
rect -1173 -3062 -1139 -3028
rect -1105 -3062 -1071 -3028
rect -1037 -3062 -1003 -3028
rect -969 -3062 -935 -3028
rect -901 -3062 -867 -3028
rect -833 -3062 -799 -3028
rect -765 -3062 -731 -3028
rect -697 -3062 -663 -3028
rect -629 -3062 -595 -3028
rect -561 -3062 -527 -3028
rect -493 -3062 -459 -3028
rect -425 -3062 -391 -3028
rect -357 -3062 -323 -3028
rect -289 -3062 -255 -3028
rect -221 -3062 -187 -3028
rect -153 -3062 -119 -3028
rect -85 -3062 -51 -3028
rect -17 -3062 17 -3028
rect 51 -3062 85 -3028
rect 119 -3062 153 -3028
rect 187 -3062 221 -3028
rect 255 -3062 289 -3028
rect 323 -3062 357 -3028
rect 391 -3062 425 -3028
rect 459 -3062 493 -3028
rect 527 -3062 561 -3028
rect 595 -3062 629 -3028
rect 663 -3062 697 -3028
rect 731 -3062 765 -3028
rect 799 -3062 833 -3028
rect 867 -3062 901 -3028
rect 935 -3062 969 -3028
rect 1003 -3062 1037 -3028
rect 1071 -3062 1105 -3028
rect 1139 -3062 1173 -3028
rect 1207 -3062 1241 -3028
rect 1275 -3062 1309 -3028
rect 1343 -3062 1377 -3028
rect 1411 -3062 1445 -3028
rect 1479 -3062 1513 -3028
rect 1547 -3062 1581 -3028
rect 1615 -3062 1649 -3028
rect 1683 -3062 1717 -3028
rect 1751 -3062 1785 -3028
rect 1819 -3062 1853 -3028
rect 1887 -3062 1921 -3028
rect 1955 -3062 1989 -3028
rect 2023 -3062 2057 -3028
rect 2091 -3062 2125 -3028
rect 2159 -3062 2193 -3028
rect 2227 -3062 2261 -3028
rect 2295 -3062 2329 -3028
rect 2363 -3062 2397 -3028
rect 2431 -3062 2465 -3028
rect 2499 -3062 2533 -3028
rect 2567 -3062 2601 -3028
rect 2635 -3062 2669 -3028
rect 2703 -3062 2737 -3028
rect 2771 -3062 2805 -3028
rect 2839 -3062 2873 -3028
rect 2907 -3062 2941 -3028
rect 2975 -3062 3009 -3028
rect 3043 -3062 3077 -3028
rect 3111 -3062 3145 -3028
rect 3179 -3062 3213 -3028
rect 3247 -3062 3281 -3028
rect 3315 -3062 3349 -3028
rect 3383 -3062 3417 -3028
rect 3451 -3062 3485 -3028
rect 3519 -3062 3553 -3028
rect 3587 -3062 3621 -3028
rect 3655 -3062 3689 -3028
rect 3723 -3062 3757 -3028
rect 3791 -3062 3825 -3028
rect 3859 -3062 3893 -3028
rect 3927 -3062 3961 -3028
rect 3995 -3062 4029 -3028
rect 4063 -3062 4097 -3028
rect 4131 -3062 4165 -3028
rect 4199 -3062 4233 -3028
rect 4267 -3062 4301 -3028
rect 4335 -3062 4369 -3028
rect 4403 -3062 4437 -3028
rect 4471 -3062 4505 -3028
rect 4539 -3062 4573 -3028
rect 4607 -3062 4641 -3028
rect 4675 -3062 4709 -3028
rect 4743 -3062 4777 -3028
rect 4811 -3062 4845 -3028
rect 4879 -3062 4913 -3028
rect 4947 -3062 4981 -3028
rect 5015 -3062 5049 -3028
rect 5083 -3062 5117 -3028
rect 5151 -3062 5185 -3028
rect 5219 -3062 5253 -3028
rect 5287 -3062 5410 -3028
<< psubdiffcont >>
rect -5287 3028 -5253 3062
rect -5219 3028 -5185 3062
rect -5151 3028 -5117 3062
rect -5083 3028 -5049 3062
rect -5015 3028 -4981 3062
rect -4947 3028 -4913 3062
rect -4879 3028 -4845 3062
rect -4811 3028 -4777 3062
rect -4743 3028 -4709 3062
rect -4675 3028 -4641 3062
rect -4607 3028 -4573 3062
rect -4539 3028 -4505 3062
rect -4471 3028 -4437 3062
rect -4403 3028 -4369 3062
rect -4335 3028 -4301 3062
rect -4267 3028 -4233 3062
rect -4199 3028 -4165 3062
rect -4131 3028 -4097 3062
rect -4063 3028 -4029 3062
rect -3995 3028 -3961 3062
rect -3927 3028 -3893 3062
rect -3859 3028 -3825 3062
rect -3791 3028 -3757 3062
rect -3723 3028 -3689 3062
rect -3655 3028 -3621 3062
rect -3587 3028 -3553 3062
rect -3519 3028 -3485 3062
rect -3451 3028 -3417 3062
rect -3383 3028 -3349 3062
rect -3315 3028 -3281 3062
rect -3247 3028 -3213 3062
rect -3179 3028 -3145 3062
rect -3111 3028 -3077 3062
rect -3043 3028 -3009 3062
rect -2975 3028 -2941 3062
rect -2907 3028 -2873 3062
rect -2839 3028 -2805 3062
rect -2771 3028 -2737 3062
rect -2703 3028 -2669 3062
rect -2635 3028 -2601 3062
rect -2567 3028 -2533 3062
rect -2499 3028 -2465 3062
rect -2431 3028 -2397 3062
rect -2363 3028 -2329 3062
rect -2295 3028 -2261 3062
rect -2227 3028 -2193 3062
rect -2159 3028 -2125 3062
rect -2091 3028 -2057 3062
rect -2023 3028 -1989 3062
rect -1955 3028 -1921 3062
rect -1887 3028 -1853 3062
rect -1819 3028 -1785 3062
rect -1751 3028 -1717 3062
rect -1683 3028 -1649 3062
rect -1615 3028 -1581 3062
rect -1547 3028 -1513 3062
rect -1479 3028 -1445 3062
rect -1411 3028 -1377 3062
rect -1343 3028 -1309 3062
rect -1275 3028 -1241 3062
rect -1207 3028 -1173 3062
rect -1139 3028 -1105 3062
rect -1071 3028 -1037 3062
rect -1003 3028 -969 3062
rect -935 3028 -901 3062
rect -867 3028 -833 3062
rect -799 3028 -765 3062
rect -731 3028 -697 3062
rect -663 3028 -629 3062
rect -595 3028 -561 3062
rect -527 3028 -493 3062
rect -459 3028 -425 3062
rect -391 3028 -357 3062
rect -323 3028 -289 3062
rect -255 3028 -221 3062
rect -187 3028 -153 3062
rect -119 3028 -85 3062
rect -51 3028 -17 3062
rect 17 3028 51 3062
rect 85 3028 119 3062
rect 153 3028 187 3062
rect 221 3028 255 3062
rect 289 3028 323 3062
rect 357 3028 391 3062
rect 425 3028 459 3062
rect 493 3028 527 3062
rect 561 3028 595 3062
rect 629 3028 663 3062
rect 697 3028 731 3062
rect 765 3028 799 3062
rect 833 3028 867 3062
rect 901 3028 935 3062
rect 969 3028 1003 3062
rect 1037 3028 1071 3062
rect 1105 3028 1139 3062
rect 1173 3028 1207 3062
rect 1241 3028 1275 3062
rect 1309 3028 1343 3062
rect 1377 3028 1411 3062
rect 1445 3028 1479 3062
rect 1513 3028 1547 3062
rect 1581 3028 1615 3062
rect 1649 3028 1683 3062
rect 1717 3028 1751 3062
rect 1785 3028 1819 3062
rect 1853 3028 1887 3062
rect 1921 3028 1955 3062
rect 1989 3028 2023 3062
rect 2057 3028 2091 3062
rect 2125 3028 2159 3062
rect 2193 3028 2227 3062
rect 2261 3028 2295 3062
rect 2329 3028 2363 3062
rect 2397 3028 2431 3062
rect 2465 3028 2499 3062
rect 2533 3028 2567 3062
rect 2601 3028 2635 3062
rect 2669 3028 2703 3062
rect 2737 3028 2771 3062
rect 2805 3028 2839 3062
rect 2873 3028 2907 3062
rect 2941 3028 2975 3062
rect 3009 3028 3043 3062
rect 3077 3028 3111 3062
rect 3145 3028 3179 3062
rect 3213 3028 3247 3062
rect 3281 3028 3315 3062
rect 3349 3028 3383 3062
rect 3417 3028 3451 3062
rect 3485 3028 3519 3062
rect 3553 3028 3587 3062
rect 3621 3028 3655 3062
rect 3689 3028 3723 3062
rect 3757 3028 3791 3062
rect 3825 3028 3859 3062
rect 3893 3028 3927 3062
rect 3961 3028 3995 3062
rect 4029 3028 4063 3062
rect 4097 3028 4131 3062
rect 4165 3028 4199 3062
rect 4233 3028 4267 3062
rect 4301 3028 4335 3062
rect 4369 3028 4403 3062
rect 4437 3028 4471 3062
rect 4505 3028 4539 3062
rect 4573 3028 4607 3062
rect 4641 3028 4675 3062
rect 4709 3028 4743 3062
rect 4777 3028 4811 3062
rect 4845 3028 4879 3062
rect 4913 3028 4947 3062
rect 4981 3028 5015 3062
rect 5049 3028 5083 3062
rect 5117 3028 5151 3062
rect 5185 3028 5219 3062
rect 5253 3028 5287 3062
rect -5410 2907 -5376 2941
rect -5410 2839 -5376 2873
rect -5410 2771 -5376 2805
rect -5410 2703 -5376 2737
rect -5410 2635 -5376 2669
rect -5410 2567 -5376 2601
rect -5410 2499 -5376 2533
rect -5410 2431 -5376 2465
rect -5410 2363 -5376 2397
rect -5410 2295 -5376 2329
rect -5410 2227 -5376 2261
rect -5410 2159 -5376 2193
rect -5410 2091 -5376 2125
rect -5410 2023 -5376 2057
rect -5410 1955 -5376 1989
rect -5410 1887 -5376 1921
rect -5410 1819 -5376 1853
rect -5410 1751 -5376 1785
rect -5410 1683 -5376 1717
rect -5410 1615 -5376 1649
rect -5410 1547 -5376 1581
rect -5410 1479 -5376 1513
rect -5410 1411 -5376 1445
rect -5410 1343 -5376 1377
rect -5410 1275 -5376 1309
rect -5410 1207 -5376 1241
rect -5410 1139 -5376 1173
rect -5410 1071 -5376 1105
rect -5410 1003 -5376 1037
rect -5410 935 -5376 969
rect -5410 867 -5376 901
rect -5410 799 -5376 833
rect -5410 731 -5376 765
rect -5410 663 -5376 697
rect -5410 595 -5376 629
rect -5410 527 -5376 561
rect -5410 459 -5376 493
rect -5410 391 -5376 425
rect -5410 323 -5376 357
rect -5410 255 -5376 289
rect -5410 187 -5376 221
rect -5410 119 -5376 153
rect -5410 51 -5376 85
rect -5410 -17 -5376 17
rect -5410 -85 -5376 -51
rect -5410 -153 -5376 -119
rect -5410 -221 -5376 -187
rect -5410 -289 -5376 -255
rect -5410 -357 -5376 -323
rect -5410 -425 -5376 -391
rect -5410 -493 -5376 -459
rect -5410 -561 -5376 -527
rect -5410 -629 -5376 -595
rect -5410 -697 -5376 -663
rect -5410 -765 -5376 -731
rect -5410 -833 -5376 -799
rect -5410 -901 -5376 -867
rect -5410 -969 -5376 -935
rect -5410 -1037 -5376 -1003
rect -5410 -1105 -5376 -1071
rect -5410 -1173 -5376 -1139
rect -5410 -1241 -5376 -1207
rect -5410 -1309 -5376 -1275
rect -5410 -1377 -5376 -1343
rect -5410 -1445 -5376 -1411
rect -5410 -1513 -5376 -1479
rect -5410 -1581 -5376 -1547
rect -5410 -1649 -5376 -1615
rect -5410 -1717 -5376 -1683
rect -5410 -1785 -5376 -1751
rect -5410 -1853 -5376 -1819
rect -5410 -1921 -5376 -1887
rect -5410 -1989 -5376 -1955
rect -5410 -2057 -5376 -2023
rect -5410 -2125 -5376 -2091
rect -5410 -2193 -5376 -2159
rect -5410 -2261 -5376 -2227
rect -5410 -2329 -5376 -2295
rect -5410 -2397 -5376 -2363
rect -5410 -2465 -5376 -2431
rect -5410 -2533 -5376 -2499
rect -5410 -2601 -5376 -2567
rect -5410 -2669 -5376 -2635
rect -5410 -2737 -5376 -2703
rect -5410 -2805 -5376 -2771
rect -5410 -2873 -5376 -2839
rect -5410 -2941 -5376 -2907
rect 5376 2907 5410 2941
rect 5376 2839 5410 2873
rect 5376 2771 5410 2805
rect 5376 2703 5410 2737
rect 5376 2635 5410 2669
rect 5376 2567 5410 2601
rect 5376 2499 5410 2533
rect 5376 2431 5410 2465
rect 5376 2363 5410 2397
rect 5376 2295 5410 2329
rect 5376 2227 5410 2261
rect 5376 2159 5410 2193
rect 5376 2091 5410 2125
rect 5376 2023 5410 2057
rect 5376 1955 5410 1989
rect 5376 1887 5410 1921
rect 5376 1819 5410 1853
rect 5376 1751 5410 1785
rect 5376 1683 5410 1717
rect 5376 1615 5410 1649
rect 5376 1547 5410 1581
rect 5376 1479 5410 1513
rect 5376 1411 5410 1445
rect 5376 1343 5410 1377
rect 5376 1275 5410 1309
rect 5376 1207 5410 1241
rect 5376 1139 5410 1173
rect 5376 1071 5410 1105
rect 5376 1003 5410 1037
rect 5376 935 5410 969
rect 5376 867 5410 901
rect 5376 799 5410 833
rect 5376 731 5410 765
rect 5376 663 5410 697
rect 5376 595 5410 629
rect 5376 527 5410 561
rect 5376 459 5410 493
rect 5376 391 5410 425
rect 5376 323 5410 357
rect 5376 255 5410 289
rect 5376 187 5410 221
rect 5376 119 5410 153
rect 5376 51 5410 85
rect 5376 -17 5410 17
rect 5376 -85 5410 -51
rect 5376 -153 5410 -119
rect 5376 -221 5410 -187
rect 5376 -289 5410 -255
rect 5376 -357 5410 -323
rect 5376 -425 5410 -391
rect 5376 -493 5410 -459
rect 5376 -561 5410 -527
rect 5376 -629 5410 -595
rect 5376 -697 5410 -663
rect 5376 -765 5410 -731
rect 5376 -833 5410 -799
rect 5376 -901 5410 -867
rect 5376 -969 5410 -935
rect 5376 -1037 5410 -1003
rect 5376 -1105 5410 -1071
rect 5376 -1173 5410 -1139
rect 5376 -1241 5410 -1207
rect 5376 -1309 5410 -1275
rect 5376 -1377 5410 -1343
rect 5376 -1445 5410 -1411
rect 5376 -1513 5410 -1479
rect 5376 -1581 5410 -1547
rect 5376 -1649 5410 -1615
rect 5376 -1717 5410 -1683
rect 5376 -1785 5410 -1751
rect 5376 -1853 5410 -1819
rect 5376 -1921 5410 -1887
rect 5376 -1989 5410 -1955
rect 5376 -2057 5410 -2023
rect 5376 -2125 5410 -2091
rect 5376 -2193 5410 -2159
rect 5376 -2261 5410 -2227
rect 5376 -2329 5410 -2295
rect 5376 -2397 5410 -2363
rect 5376 -2465 5410 -2431
rect 5376 -2533 5410 -2499
rect 5376 -2601 5410 -2567
rect 5376 -2669 5410 -2635
rect 5376 -2737 5410 -2703
rect 5376 -2805 5410 -2771
rect 5376 -2873 5410 -2839
rect 5376 -2941 5410 -2907
rect -5287 -3062 -5253 -3028
rect -5219 -3062 -5185 -3028
rect -5151 -3062 -5117 -3028
rect -5083 -3062 -5049 -3028
rect -5015 -3062 -4981 -3028
rect -4947 -3062 -4913 -3028
rect -4879 -3062 -4845 -3028
rect -4811 -3062 -4777 -3028
rect -4743 -3062 -4709 -3028
rect -4675 -3062 -4641 -3028
rect -4607 -3062 -4573 -3028
rect -4539 -3062 -4505 -3028
rect -4471 -3062 -4437 -3028
rect -4403 -3062 -4369 -3028
rect -4335 -3062 -4301 -3028
rect -4267 -3062 -4233 -3028
rect -4199 -3062 -4165 -3028
rect -4131 -3062 -4097 -3028
rect -4063 -3062 -4029 -3028
rect -3995 -3062 -3961 -3028
rect -3927 -3062 -3893 -3028
rect -3859 -3062 -3825 -3028
rect -3791 -3062 -3757 -3028
rect -3723 -3062 -3689 -3028
rect -3655 -3062 -3621 -3028
rect -3587 -3062 -3553 -3028
rect -3519 -3062 -3485 -3028
rect -3451 -3062 -3417 -3028
rect -3383 -3062 -3349 -3028
rect -3315 -3062 -3281 -3028
rect -3247 -3062 -3213 -3028
rect -3179 -3062 -3145 -3028
rect -3111 -3062 -3077 -3028
rect -3043 -3062 -3009 -3028
rect -2975 -3062 -2941 -3028
rect -2907 -3062 -2873 -3028
rect -2839 -3062 -2805 -3028
rect -2771 -3062 -2737 -3028
rect -2703 -3062 -2669 -3028
rect -2635 -3062 -2601 -3028
rect -2567 -3062 -2533 -3028
rect -2499 -3062 -2465 -3028
rect -2431 -3062 -2397 -3028
rect -2363 -3062 -2329 -3028
rect -2295 -3062 -2261 -3028
rect -2227 -3062 -2193 -3028
rect -2159 -3062 -2125 -3028
rect -2091 -3062 -2057 -3028
rect -2023 -3062 -1989 -3028
rect -1955 -3062 -1921 -3028
rect -1887 -3062 -1853 -3028
rect -1819 -3062 -1785 -3028
rect -1751 -3062 -1717 -3028
rect -1683 -3062 -1649 -3028
rect -1615 -3062 -1581 -3028
rect -1547 -3062 -1513 -3028
rect -1479 -3062 -1445 -3028
rect -1411 -3062 -1377 -3028
rect -1343 -3062 -1309 -3028
rect -1275 -3062 -1241 -3028
rect -1207 -3062 -1173 -3028
rect -1139 -3062 -1105 -3028
rect -1071 -3062 -1037 -3028
rect -1003 -3062 -969 -3028
rect -935 -3062 -901 -3028
rect -867 -3062 -833 -3028
rect -799 -3062 -765 -3028
rect -731 -3062 -697 -3028
rect -663 -3062 -629 -3028
rect -595 -3062 -561 -3028
rect -527 -3062 -493 -3028
rect -459 -3062 -425 -3028
rect -391 -3062 -357 -3028
rect -323 -3062 -289 -3028
rect -255 -3062 -221 -3028
rect -187 -3062 -153 -3028
rect -119 -3062 -85 -3028
rect -51 -3062 -17 -3028
rect 17 -3062 51 -3028
rect 85 -3062 119 -3028
rect 153 -3062 187 -3028
rect 221 -3062 255 -3028
rect 289 -3062 323 -3028
rect 357 -3062 391 -3028
rect 425 -3062 459 -3028
rect 493 -3062 527 -3028
rect 561 -3062 595 -3028
rect 629 -3062 663 -3028
rect 697 -3062 731 -3028
rect 765 -3062 799 -3028
rect 833 -3062 867 -3028
rect 901 -3062 935 -3028
rect 969 -3062 1003 -3028
rect 1037 -3062 1071 -3028
rect 1105 -3062 1139 -3028
rect 1173 -3062 1207 -3028
rect 1241 -3062 1275 -3028
rect 1309 -3062 1343 -3028
rect 1377 -3062 1411 -3028
rect 1445 -3062 1479 -3028
rect 1513 -3062 1547 -3028
rect 1581 -3062 1615 -3028
rect 1649 -3062 1683 -3028
rect 1717 -3062 1751 -3028
rect 1785 -3062 1819 -3028
rect 1853 -3062 1887 -3028
rect 1921 -3062 1955 -3028
rect 1989 -3062 2023 -3028
rect 2057 -3062 2091 -3028
rect 2125 -3062 2159 -3028
rect 2193 -3062 2227 -3028
rect 2261 -3062 2295 -3028
rect 2329 -3062 2363 -3028
rect 2397 -3062 2431 -3028
rect 2465 -3062 2499 -3028
rect 2533 -3062 2567 -3028
rect 2601 -3062 2635 -3028
rect 2669 -3062 2703 -3028
rect 2737 -3062 2771 -3028
rect 2805 -3062 2839 -3028
rect 2873 -3062 2907 -3028
rect 2941 -3062 2975 -3028
rect 3009 -3062 3043 -3028
rect 3077 -3062 3111 -3028
rect 3145 -3062 3179 -3028
rect 3213 -3062 3247 -3028
rect 3281 -3062 3315 -3028
rect 3349 -3062 3383 -3028
rect 3417 -3062 3451 -3028
rect 3485 -3062 3519 -3028
rect 3553 -3062 3587 -3028
rect 3621 -3062 3655 -3028
rect 3689 -3062 3723 -3028
rect 3757 -3062 3791 -3028
rect 3825 -3062 3859 -3028
rect 3893 -3062 3927 -3028
rect 3961 -3062 3995 -3028
rect 4029 -3062 4063 -3028
rect 4097 -3062 4131 -3028
rect 4165 -3062 4199 -3028
rect 4233 -3062 4267 -3028
rect 4301 -3062 4335 -3028
rect 4369 -3062 4403 -3028
rect 4437 -3062 4471 -3028
rect 4505 -3062 4539 -3028
rect 4573 -3062 4607 -3028
rect 4641 -3062 4675 -3028
rect 4709 -3062 4743 -3028
rect 4777 -3062 4811 -3028
rect 4845 -3062 4879 -3028
rect 4913 -3062 4947 -3028
rect 4981 -3062 5015 -3028
rect 5049 -3062 5083 -3028
rect 5117 -3062 5151 -3028
rect 5185 -3062 5219 -3028
rect 5253 -3062 5287 -3028
<< xpolycontact >>
rect -5280 2500 -5142 2932
rect -5280 -2932 -5142 -2500
rect -4894 2500 -4756 2932
rect -4894 -2932 -4756 -2500
rect -4508 2500 -4370 2932
rect -4508 -2932 -4370 -2500
rect -4122 2500 -3984 2932
rect -4122 -2932 -3984 -2500
rect -3736 2500 -3598 2932
rect -3736 -2932 -3598 -2500
rect -3350 2500 -3212 2932
rect -3350 -2932 -3212 -2500
rect -2964 2500 -2826 2932
rect -2964 -2932 -2826 -2500
rect -2578 2500 -2440 2932
rect -2578 -2932 -2440 -2500
rect -2192 2500 -2054 2932
rect -2192 -2932 -2054 -2500
rect -1806 2500 -1668 2932
rect -1806 -2932 -1668 -2500
rect -1420 2500 -1282 2932
rect -1420 -2932 -1282 -2500
rect -1034 2500 -896 2932
rect -1034 -2932 -896 -2500
rect -648 2500 -510 2932
rect -648 -2932 -510 -2500
rect -262 2500 -124 2932
rect -262 -2932 -124 -2500
rect 124 2500 262 2932
rect 124 -2932 262 -2500
rect 510 2500 648 2932
rect 510 -2932 648 -2500
rect 896 2500 1034 2932
rect 896 -2932 1034 -2500
rect 1282 2500 1420 2932
rect 1282 -2932 1420 -2500
rect 1668 2500 1806 2932
rect 1668 -2932 1806 -2500
rect 2054 2500 2192 2932
rect 2054 -2932 2192 -2500
rect 2440 2500 2578 2932
rect 2440 -2932 2578 -2500
rect 2826 2500 2964 2932
rect 2826 -2932 2964 -2500
rect 3212 2500 3350 2932
rect 3212 -2932 3350 -2500
rect 3598 2500 3736 2932
rect 3598 -2932 3736 -2500
rect 3984 2500 4122 2932
rect 3984 -2932 4122 -2500
rect 4370 2500 4508 2932
rect 4370 -2932 4508 -2500
rect 4756 2500 4894 2932
rect 4756 -2932 4894 -2500
rect 5142 2500 5280 2932
rect 5142 -2932 5280 -2500
<< xpolyres >>
rect -5280 -2500 -5142 2500
rect -4894 -2500 -4756 2500
rect -4508 -2500 -4370 2500
rect -4122 -2500 -3984 2500
rect -3736 -2500 -3598 2500
rect -3350 -2500 -3212 2500
rect -2964 -2500 -2826 2500
rect -2578 -2500 -2440 2500
rect -2192 -2500 -2054 2500
rect -1806 -2500 -1668 2500
rect -1420 -2500 -1282 2500
rect -1034 -2500 -896 2500
rect -648 -2500 -510 2500
rect -262 -2500 -124 2500
rect 124 -2500 262 2500
rect 510 -2500 648 2500
rect 896 -2500 1034 2500
rect 1282 -2500 1420 2500
rect 1668 -2500 1806 2500
rect 2054 -2500 2192 2500
rect 2440 -2500 2578 2500
rect 2826 -2500 2964 2500
rect 3212 -2500 3350 2500
rect 3598 -2500 3736 2500
rect 3984 -2500 4122 2500
rect 4370 -2500 4508 2500
rect 4756 -2500 4894 2500
rect 5142 -2500 5280 2500
<< locali >>
rect -5410 3028 -5287 3062
rect -5253 3028 -5219 3062
rect -5185 3028 -5151 3062
rect -5117 3028 -5083 3062
rect -5049 3028 -5015 3062
rect -4981 3028 -4947 3062
rect -4913 3028 -4879 3062
rect -4845 3028 -4811 3062
rect -4777 3028 -4743 3062
rect -4709 3028 -4675 3062
rect -4641 3028 -4607 3062
rect -4573 3028 -4539 3062
rect -4505 3028 -4471 3062
rect -4437 3028 -4403 3062
rect -4369 3028 -4335 3062
rect -4301 3028 -4267 3062
rect -4233 3028 -4199 3062
rect -4165 3028 -4131 3062
rect -4097 3028 -4063 3062
rect -4029 3028 -3995 3062
rect -3961 3028 -3927 3062
rect -3893 3028 -3859 3062
rect -3825 3028 -3791 3062
rect -3757 3028 -3723 3062
rect -3689 3028 -3655 3062
rect -3621 3028 -3587 3062
rect -3553 3028 -3519 3062
rect -3485 3028 -3451 3062
rect -3417 3028 -3383 3062
rect -3349 3028 -3315 3062
rect -3281 3028 -3247 3062
rect -3213 3028 -3179 3062
rect -3145 3028 -3111 3062
rect -3077 3028 -3043 3062
rect -3009 3028 -2975 3062
rect -2941 3028 -2907 3062
rect -2873 3028 -2839 3062
rect -2805 3028 -2771 3062
rect -2737 3028 -2703 3062
rect -2669 3028 -2635 3062
rect -2601 3028 -2567 3062
rect -2533 3028 -2499 3062
rect -2465 3028 -2431 3062
rect -2397 3028 -2363 3062
rect -2329 3028 -2295 3062
rect -2261 3028 -2227 3062
rect -2193 3028 -2159 3062
rect -2125 3028 -2091 3062
rect -2057 3028 -2023 3062
rect -1989 3028 -1955 3062
rect -1921 3028 -1887 3062
rect -1853 3028 -1819 3062
rect -1785 3028 -1751 3062
rect -1717 3028 -1683 3062
rect -1649 3028 -1615 3062
rect -1581 3028 -1547 3062
rect -1513 3028 -1479 3062
rect -1445 3028 -1411 3062
rect -1377 3028 -1343 3062
rect -1309 3028 -1275 3062
rect -1241 3028 -1207 3062
rect -1173 3028 -1139 3062
rect -1105 3028 -1071 3062
rect -1037 3028 -1003 3062
rect -969 3028 -935 3062
rect -901 3028 -867 3062
rect -833 3028 -799 3062
rect -765 3028 -731 3062
rect -697 3028 -663 3062
rect -629 3028 -595 3062
rect -561 3028 -527 3062
rect -493 3028 -459 3062
rect -425 3028 -391 3062
rect -357 3028 -323 3062
rect -289 3028 -255 3062
rect -221 3028 -187 3062
rect -153 3028 -119 3062
rect -85 3028 -51 3062
rect -17 3028 17 3062
rect 51 3028 85 3062
rect 119 3028 153 3062
rect 187 3028 221 3062
rect 255 3028 289 3062
rect 323 3028 357 3062
rect 391 3028 425 3062
rect 459 3028 493 3062
rect 527 3028 561 3062
rect 595 3028 629 3062
rect 663 3028 697 3062
rect 731 3028 765 3062
rect 799 3028 833 3062
rect 867 3028 901 3062
rect 935 3028 969 3062
rect 1003 3028 1037 3062
rect 1071 3028 1105 3062
rect 1139 3028 1173 3062
rect 1207 3028 1241 3062
rect 1275 3028 1309 3062
rect 1343 3028 1377 3062
rect 1411 3028 1445 3062
rect 1479 3028 1513 3062
rect 1547 3028 1581 3062
rect 1615 3028 1649 3062
rect 1683 3028 1717 3062
rect 1751 3028 1785 3062
rect 1819 3028 1853 3062
rect 1887 3028 1921 3062
rect 1955 3028 1989 3062
rect 2023 3028 2057 3062
rect 2091 3028 2125 3062
rect 2159 3028 2193 3062
rect 2227 3028 2261 3062
rect 2295 3028 2329 3062
rect 2363 3028 2397 3062
rect 2431 3028 2465 3062
rect 2499 3028 2533 3062
rect 2567 3028 2601 3062
rect 2635 3028 2669 3062
rect 2703 3028 2737 3062
rect 2771 3028 2805 3062
rect 2839 3028 2873 3062
rect 2907 3028 2941 3062
rect 2975 3028 3009 3062
rect 3043 3028 3077 3062
rect 3111 3028 3145 3062
rect 3179 3028 3213 3062
rect 3247 3028 3281 3062
rect 3315 3028 3349 3062
rect 3383 3028 3417 3062
rect 3451 3028 3485 3062
rect 3519 3028 3553 3062
rect 3587 3028 3621 3062
rect 3655 3028 3689 3062
rect 3723 3028 3757 3062
rect 3791 3028 3825 3062
rect 3859 3028 3893 3062
rect 3927 3028 3961 3062
rect 3995 3028 4029 3062
rect 4063 3028 4097 3062
rect 4131 3028 4165 3062
rect 4199 3028 4233 3062
rect 4267 3028 4301 3062
rect 4335 3028 4369 3062
rect 4403 3028 4437 3062
rect 4471 3028 4505 3062
rect 4539 3028 4573 3062
rect 4607 3028 4641 3062
rect 4675 3028 4709 3062
rect 4743 3028 4777 3062
rect 4811 3028 4845 3062
rect 4879 3028 4913 3062
rect 4947 3028 4981 3062
rect 5015 3028 5049 3062
rect 5083 3028 5117 3062
rect 5151 3028 5185 3062
rect 5219 3028 5253 3062
rect 5287 3028 5410 3062
rect -5410 2941 -5376 3028
rect 5376 2941 5410 3028
rect -5410 2873 -5376 2907
rect -5410 2805 -5376 2839
rect -5410 2737 -5376 2771
rect -5410 2669 -5376 2683
rect -5410 2601 -5376 2611
rect -5410 2533 -5376 2539
rect 5376 2873 5410 2907
rect 5376 2805 5410 2839
rect 5376 2737 5410 2771
rect 5376 2669 5410 2683
rect 5376 2601 5410 2611
rect 5376 2533 5410 2539
rect -5410 2465 -5376 2467
rect -5410 2429 -5376 2431
rect -5410 2357 -5376 2363
rect -5410 2285 -5376 2295
rect -5410 2213 -5376 2227
rect -5410 2141 -5376 2159
rect -5410 2069 -5376 2091
rect -5410 1997 -5376 2023
rect -5410 1925 -5376 1955
rect -5410 1853 -5376 1887
rect -5410 1785 -5376 1819
rect -5410 1717 -5376 1747
rect -5410 1649 -5376 1675
rect -5410 1581 -5376 1603
rect -5410 1513 -5376 1531
rect -5410 1445 -5376 1459
rect -5410 1377 -5376 1387
rect -5410 1309 -5376 1315
rect -5410 1241 -5376 1243
rect -5410 1205 -5376 1207
rect -5410 1133 -5376 1139
rect -5410 1061 -5376 1071
rect -5410 989 -5376 1003
rect -5410 917 -5376 935
rect -5410 845 -5376 867
rect -5410 773 -5376 799
rect -5410 701 -5376 731
rect -5410 629 -5376 663
rect -5410 561 -5376 595
rect -5410 493 -5376 523
rect -5410 425 -5376 451
rect -5410 357 -5376 379
rect -5410 289 -5376 307
rect -5410 221 -5376 235
rect -5410 153 -5376 163
rect -5410 85 -5376 91
rect -5410 17 -5376 19
rect -5410 -19 -5376 -17
rect -5410 -91 -5376 -85
rect -5410 -163 -5376 -153
rect -5410 -235 -5376 -221
rect -5410 -307 -5376 -289
rect -5410 -379 -5376 -357
rect -5410 -451 -5376 -425
rect -5410 -523 -5376 -493
rect -5410 -595 -5376 -561
rect -5410 -663 -5376 -629
rect -5410 -731 -5376 -701
rect -5410 -799 -5376 -773
rect -5410 -867 -5376 -845
rect -5410 -935 -5376 -917
rect -5410 -1003 -5376 -989
rect -5410 -1071 -5376 -1061
rect -5410 -1139 -5376 -1133
rect -5410 -1207 -5376 -1205
rect -5410 -1243 -5376 -1241
rect -5410 -1315 -5376 -1309
rect -5410 -1387 -5376 -1377
rect -5410 -1459 -5376 -1445
rect -5410 -1531 -5376 -1513
rect -5410 -1603 -5376 -1581
rect -5410 -1675 -5376 -1649
rect -5410 -1747 -5376 -1717
rect -5410 -1819 -5376 -1785
rect -5410 -1887 -5376 -1853
rect -5410 -1955 -5376 -1925
rect -5410 -2023 -5376 -1997
rect -5410 -2091 -5376 -2069
rect -5410 -2159 -5376 -2141
rect -5410 -2227 -5376 -2213
rect -5410 -2295 -5376 -2285
rect -5410 -2363 -5376 -2357
rect -5410 -2431 -5376 -2429
rect -5410 -2467 -5376 -2465
rect 5376 2465 5410 2467
rect 5376 2429 5410 2431
rect 5376 2357 5410 2363
rect 5376 2285 5410 2295
rect 5376 2213 5410 2227
rect 5376 2141 5410 2159
rect 5376 2069 5410 2091
rect 5376 1997 5410 2023
rect 5376 1925 5410 1955
rect 5376 1853 5410 1887
rect 5376 1785 5410 1819
rect 5376 1717 5410 1747
rect 5376 1649 5410 1675
rect 5376 1581 5410 1603
rect 5376 1513 5410 1531
rect 5376 1445 5410 1459
rect 5376 1377 5410 1387
rect 5376 1309 5410 1315
rect 5376 1241 5410 1243
rect 5376 1205 5410 1207
rect 5376 1133 5410 1139
rect 5376 1061 5410 1071
rect 5376 989 5410 1003
rect 5376 917 5410 935
rect 5376 845 5410 867
rect 5376 773 5410 799
rect 5376 701 5410 731
rect 5376 629 5410 663
rect 5376 561 5410 595
rect 5376 493 5410 523
rect 5376 425 5410 451
rect 5376 357 5410 379
rect 5376 289 5410 307
rect 5376 221 5410 235
rect 5376 153 5410 163
rect 5376 85 5410 91
rect 5376 17 5410 19
rect 5376 -19 5410 -17
rect 5376 -91 5410 -85
rect 5376 -163 5410 -153
rect 5376 -235 5410 -221
rect 5376 -307 5410 -289
rect 5376 -379 5410 -357
rect 5376 -451 5410 -425
rect 5376 -523 5410 -493
rect 5376 -595 5410 -561
rect 5376 -663 5410 -629
rect 5376 -731 5410 -701
rect 5376 -799 5410 -773
rect 5376 -867 5410 -845
rect 5376 -935 5410 -917
rect 5376 -1003 5410 -989
rect 5376 -1071 5410 -1061
rect 5376 -1139 5410 -1133
rect 5376 -1207 5410 -1205
rect 5376 -1243 5410 -1241
rect 5376 -1315 5410 -1309
rect 5376 -1387 5410 -1377
rect 5376 -1459 5410 -1445
rect 5376 -1531 5410 -1513
rect 5376 -1603 5410 -1581
rect 5376 -1675 5410 -1649
rect 5376 -1747 5410 -1717
rect 5376 -1819 5410 -1785
rect 5376 -1887 5410 -1853
rect 5376 -1955 5410 -1925
rect 5376 -2023 5410 -1997
rect 5376 -2091 5410 -2069
rect 5376 -2159 5410 -2141
rect 5376 -2227 5410 -2213
rect 5376 -2295 5410 -2285
rect 5376 -2363 5410 -2357
rect 5376 -2431 5410 -2429
rect 5376 -2467 5410 -2465
rect -5410 -2539 -5376 -2533
rect -5410 -2611 -5376 -2601
rect -5410 -2683 -5376 -2669
rect -5410 -2771 -5376 -2737
rect -5410 -2839 -5376 -2805
rect -5410 -2907 -5376 -2873
rect 5376 -2539 5410 -2533
rect 5376 -2611 5410 -2601
rect 5376 -2683 5410 -2669
rect 5376 -2771 5410 -2737
rect 5376 -2839 5410 -2805
rect 5376 -2907 5410 -2873
rect -5410 -3028 -5376 -2941
rect 5376 -3028 5410 -2941
rect -5410 -3062 -5287 -3028
rect -5253 -3062 -5219 -3028
rect -5185 -3062 -5151 -3028
rect -5117 -3062 -5083 -3028
rect -5049 -3062 -5015 -3028
rect -4981 -3062 -4947 -3028
rect -4913 -3062 -4879 -3028
rect -4845 -3062 -4811 -3028
rect -4771 -3062 -4743 -3028
rect -4699 -3062 -4675 -3028
rect -4627 -3062 -4607 -3028
rect -4555 -3062 -4539 -3028
rect -4483 -3062 -4471 -3028
rect -4411 -3062 -4403 -3028
rect -4339 -3062 -4335 -3028
rect -4233 -3062 -4229 -3028
rect -4165 -3062 -4157 -3028
rect -4097 -3062 -4085 -3028
rect -4029 -3062 -4013 -3028
rect -3961 -3062 -3941 -3028
rect -3893 -3062 -3869 -3028
rect -3825 -3062 -3797 -3028
rect -3757 -3062 -3725 -3028
rect -3689 -3062 -3655 -3028
rect -3619 -3062 -3587 -3028
rect -3547 -3062 -3519 -3028
rect -3475 -3062 -3451 -3028
rect -3403 -3062 -3383 -3028
rect -3331 -3062 -3315 -3028
rect -3259 -3062 -3247 -3028
rect -3187 -3062 -3179 -3028
rect -3115 -3062 -3111 -3028
rect -3009 -3062 -3005 -3028
rect -2941 -3062 -2933 -3028
rect -2873 -3062 -2861 -3028
rect -2805 -3062 -2789 -3028
rect -2737 -3062 -2717 -3028
rect -2669 -3062 -2645 -3028
rect -2601 -3062 -2573 -3028
rect -2533 -3062 -2501 -3028
rect -2465 -3062 -2431 -3028
rect -2395 -3062 -2363 -3028
rect -2323 -3062 -2295 -3028
rect -2251 -3062 -2227 -3028
rect -2179 -3062 -2159 -3028
rect -2107 -3062 -2091 -3028
rect -2035 -3062 -2023 -3028
rect -1963 -3062 -1955 -3028
rect -1891 -3062 -1887 -3028
rect -1785 -3062 -1781 -3028
rect -1717 -3062 -1709 -3028
rect -1649 -3062 -1637 -3028
rect -1581 -3062 -1565 -3028
rect -1513 -3062 -1493 -3028
rect -1445 -3062 -1421 -3028
rect -1377 -3062 -1349 -3028
rect -1309 -3062 -1277 -3028
rect -1241 -3062 -1207 -3028
rect -1171 -3062 -1139 -3028
rect -1099 -3062 -1071 -3028
rect -1027 -3062 -1003 -3028
rect -955 -3062 -935 -3028
rect -883 -3062 -867 -3028
rect -811 -3062 -799 -3028
rect -739 -3062 -731 -3028
rect -667 -3062 -663 -3028
rect -561 -3062 -557 -3028
rect -493 -3062 -485 -3028
rect -425 -3062 -413 -3028
rect -357 -3062 -341 -3028
rect -289 -3062 -269 -3028
rect -221 -3062 -197 -3028
rect -153 -3062 -125 -3028
rect -85 -3062 -53 -3028
rect -17 -3062 17 -3028
rect 53 -3062 85 -3028
rect 125 -3062 153 -3028
rect 197 -3062 221 -3028
rect 269 -3062 289 -3028
rect 341 -3062 357 -3028
rect 413 -3062 425 -3028
rect 485 -3062 493 -3028
rect 557 -3062 561 -3028
rect 663 -3062 667 -3028
rect 731 -3062 739 -3028
rect 799 -3062 811 -3028
rect 867 -3062 883 -3028
rect 935 -3062 955 -3028
rect 1003 -3062 1027 -3028
rect 1071 -3062 1099 -3028
rect 1139 -3062 1171 -3028
rect 1207 -3062 1241 -3028
rect 1277 -3062 1309 -3028
rect 1349 -3062 1377 -3028
rect 1421 -3062 1445 -3028
rect 1493 -3062 1513 -3028
rect 1565 -3062 1581 -3028
rect 1637 -3062 1649 -3028
rect 1709 -3062 1717 -3028
rect 1781 -3062 1785 -3028
rect 1887 -3062 1891 -3028
rect 1955 -3062 1963 -3028
rect 2023 -3062 2035 -3028
rect 2091 -3062 2107 -3028
rect 2159 -3062 2179 -3028
rect 2227 -3062 2251 -3028
rect 2295 -3062 2323 -3028
rect 2363 -3062 2395 -3028
rect 2431 -3062 2465 -3028
rect 2501 -3062 2533 -3028
rect 2573 -3062 2601 -3028
rect 2645 -3062 2669 -3028
rect 2717 -3062 2737 -3028
rect 2789 -3062 2805 -3028
rect 2861 -3062 2873 -3028
rect 2933 -3062 2941 -3028
rect 3005 -3062 3009 -3028
rect 3111 -3062 3115 -3028
rect 3179 -3062 3187 -3028
rect 3247 -3062 3259 -3028
rect 3315 -3062 3331 -3028
rect 3383 -3062 3403 -3028
rect 3451 -3062 3475 -3028
rect 3519 -3062 3547 -3028
rect 3587 -3062 3619 -3028
rect 3655 -3062 3689 -3028
rect 3725 -3062 3757 -3028
rect 3797 -3062 3825 -3028
rect 3869 -3062 3893 -3028
rect 3941 -3062 3961 -3028
rect 4013 -3062 4029 -3028
rect 4085 -3062 4097 -3028
rect 4157 -3062 4165 -3028
rect 4229 -3062 4233 -3028
rect 4335 -3062 4339 -3028
rect 4403 -3062 4411 -3028
rect 4471 -3062 4483 -3028
rect 4539 -3062 4555 -3028
rect 4607 -3062 4627 -3028
rect 4675 -3062 4699 -3028
rect 4743 -3062 4771 -3028
rect 4811 -3062 4845 -3028
rect 4879 -3062 4913 -3028
rect 4947 -3062 4981 -3028
rect 5015 -3062 5049 -3028
rect 5083 -3062 5117 -3028
rect 5151 -3062 5185 -3028
rect 5219 -3062 5253 -3028
rect 5287 -3062 5410 -3028
<< viali >>
rect -5410 2703 -5376 2717
rect -5410 2683 -5376 2703
rect -5410 2635 -5376 2645
rect -5410 2611 -5376 2635
rect -5410 2567 -5376 2573
rect -5410 2539 -5376 2567
rect -5410 2499 -5376 2501
rect 5376 2703 5410 2717
rect 5376 2683 5410 2703
rect 5376 2635 5410 2645
rect 5376 2611 5410 2635
rect 5376 2567 5410 2573
rect 5376 2539 5410 2567
rect -5410 2467 -5376 2499
rect -5410 2397 -5376 2429
rect -5410 2395 -5376 2397
rect -5410 2329 -5376 2357
rect -5410 2323 -5376 2329
rect -5410 2261 -5376 2285
rect -5410 2251 -5376 2261
rect -5410 2193 -5376 2213
rect -5410 2179 -5376 2193
rect -5410 2125 -5376 2141
rect -5410 2107 -5376 2125
rect -5410 2057 -5376 2069
rect -5410 2035 -5376 2057
rect -5410 1989 -5376 1997
rect -5410 1963 -5376 1989
rect -5410 1921 -5376 1925
rect -5410 1891 -5376 1921
rect -5410 1819 -5376 1853
rect -5410 1751 -5376 1781
rect -5410 1747 -5376 1751
rect -5410 1683 -5376 1709
rect -5410 1675 -5376 1683
rect -5410 1615 -5376 1637
rect -5410 1603 -5376 1615
rect -5410 1547 -5376 1565
rect -5410 1531 -5376 1547
rect -5410 1479 -5376 1493
rect -5410 1459 -5376 1479
rect -5410 1411 -5376 1421
rect -5410 1387 -5376 1411
rect -5410 1343 -5376 1349
rect -5410 1315 -5376 1343
rect -5410 1275 -5376 1277
rect -5410 1243 -5376 1275
rect -5410 1173 -5376 1205
rect -5410 1171 -5376 1173
rect -5410 1105 -5376 1133
rect -5410 1099 -5376 1105
rect -5410 1037 -5376 1061
rect -5410 1027 -5376 1037
rect -5410 969 -5376 989
rect -5410 955 -5376 969
rect -5410 901 -5376 917
rect -5410 883 -5376 901
rect -5410 833 -5376 845
rect -5410 811 -5376 833
rect -5410 765 -5376 773
rect -5410 739 -5376 765
rect -5410 697 -5376 701
rect -5410 667 -5376 697
rect -5410 595 -5376 629
rect -5410 527 -5376 557
rect -5410 523 -5376 527
rect -5410 459 -5376 485
rect -5410 451 -5376 459
rect -5410 391 -5376 413
rect -5410 379 -5376 391
rect -5410 323 -5376 341
rect -5410 307 -5376 323
rect -5410 255 -5376 269
rect -5410 235 -5376 255
rect -5410 187 -5376 197
rect -5410 163 -5376 187
rect -5410 119 -5376 125
rect -5410 91 -5376 119
rect -5410 51 -5376 53
rect -5410 19 -5376 51
rect -5410 -51 -5376 -19
rect -5410 -53 -5376 -51
rect -5410 -119 -5376 -91
rect -5410 -125 -5376 -119
rect -5410 -187 -5376 -163
rect -5410 -197 -5376 -187
rect -5410 -255 -5376 -235
rect -5410 -269 -5376 -255
rect -5410 -323 -5376 -307
rect -5410 -341 -5376 -323
rect -5410 -391 -5376 -379
rect -5410 -413 -5376 -391
rect -5410 -459 -5376 -451
rect -5410 -485 -5376 -459
rect -5410 -527 -5376 -523
rect -5410 -557 -5376 -527
rect -5410 -629 -5376 -595
rect -5410 -697 -5376 -667
rect -5410 -701 -5376 -697
rect -5410 -765 -5376 -739
rect -5410 -773 -5376 -765
rect -5410 -833 -5376 -811
rect -5410 -845 -5376 -833
rect -5410 -901 -5376 -883
rect -5410 -917 -5376 -901
rect -5410 -969 -5376 -955
rect -5410 -989 -5376 -969
rect -5410 -1037 -5376 -1027
rect -5410 -1061 -5376 -1037
rect -5410 -1105 -5376 -1099
rect -5410 -1133 -5376 -1105
rect -5410 -1173 -5376 -1171
rect -5410 -1205 -5376 -1173
rect -5410 -1275 -5376 -1243
rect -5410 -1277 -5376 -1275
rect -5410 -1343 -5376 -1315
rect -5410 -1349 -5376 -1343
rect -5410 -1411 -5376 -1387
rect -5410 -1421 -5376 -1411
rect -5410 -1479 -5376 -1459
rect -5410 -1493 -5376 -1479
rect -5410 -1547 -5376 -1531
rect -5410 -1565 -5376 -1547
rect -5410 -1615 -5376 -1603
rect -5410 -1637 -5376 -1615
rect -5410 -1683 -5376 -1675
rect -5410 -1709 -5376 -1683
rect -5410 -1751 -5376 -1747
rect -5410 -1781 -5376 -1751
rect -5410 -1853 -5376 -1819
rect -5410 -1921 -5376 -1891
rect -5410 -1925 -5376 -1921
rect -5410 -1989 -5376 -1963
rect -5410 -1997 -5376 -1989
rect -5410 -2057 -5376 -2035
rect -5410 -2069 -5376 -2057
rect -5410 -2125 -5376 -2107
rect -5410 -2141 -5376 -2125
rect -5410 -2193 -5376 -2179
rect -5410 -2213 -5376 -2193
rect -5410 -2261 -5376 -2251
rect -5410 -2285 -5376 -2261
rect -5410 -2329 -5376 -2323
rect -5410 -2357 -5376 -2329
rect -5410 -2397 -5376 -2395
rect -5410 -2429 -5376 -2397
rect -5410 -2499 -5376 -2467
rect -5410 -2501 -5376 -2499
rect 5376 2499 5410 2501
rect 5376 2467 5410 2499
rect 5376 2397 5410 2429
rect 5376 2395 5410 2397
rect 5376 2329 5410 2357
rect 5376 2323 5410 2329
rect 5376 2261 5410 2285
rect 5376 2251 5410 2261
rect 5376 2193 5410 2213
rect 5376 2179 5410 2193
rect 5376 2125 5410 2141
rect 5376 2107 5410 2125
rect 5376 2057 5410 2069
rect 5376 2035 5410 2057
rect 5376 1989 5410 1997
rect 5376 1963 5410 1989
rect 5376 1921 5410 1925
rect 5376 1891 5410 1921
rect 5376 1819 5410 1853
rect 5376 1751 5410 1781
rect 5376 1747 5410 1751
rect 5376 1683 5410 1709
rect 5376 1675 5410 1683
rect 5376 1615 5410 1637
rect 5376 1603 5410 1615
rect 5376 1547 5410 1565
rect 5376 1531 5410 1547
rect 5376 1479 5410 1493
rect 5376 1459 5410 1479
rect 5376 1411 5410 1421
rect 5376 1387 5410 1411
rect 5376 1343 5410 1349
rect 5376 1315 5410 1343
rect 5376 1275 5410 1277
rect 5376 1243 5410 1275
rect 5376 1173 5410 1205
rect 5376 1171 5410 1173
rect 5376 1105 5410 1133
rect 5376 1099 5410 1105
rect 5376 1037 5410 1061
rect 5376 1027 5410 1037
rect 5376 969 5410 989
rect 5376 955 5410 969
rect 5376 901 5410 917
rect 5376 883 5410 901
rect 5376 833 5410 845
rect 5376 811 5410 833
rect 5376 765 5410 773
rect 5376 739 5410 765
rect 5376 697 5410 701
rect 5376 667 5410 697
rect 5376 595 5410 629
rect 5376 527 5410 557
rect 5376 523 5410 527
rect 5376 459 5410 485
rect 5376 451 5410 459
rect 5376 391 5410 413
rect 5376 379 5410 391
rect 5376 323 5410 341
rect 5376 307 5410 323
rect 5376 255 5410 269
rect 5376 235 5410 255
rect 5376 187 5410 197
rect 5376 163 5410 187
rect 5376 119 5410 125
rect 5376 91 5410 119
rect 5376 51 5410 53
rect 5376 19 5410 51
rect 5376 -51 5410 -19
rect 5376 -53 5410 -51
rect 5376 -119 5410 -91
rect 5376 -125 5410 -119
rect 5376 -187 5410 -163
rect 5376 -197 5410 -187
rect 5376 -255 5410 -235
rect 5376 -269 5410 -255
rect 5376 -323 5410 -307
rect 5376 -341 5410 -323
rect 5376 -391 5410 -379
rect 5376 -413 5410 -391
rect 5376 -459 5410 -451
rect 5376 -485 5410 -459
rect 5376 -527 5410 -523
rect 5376 -557 5410 -527
rect 5376 -629 5410 -595
rect 5376 -697 5410 -667
rect 5376 -701 5410 -697
rect 5376 -765 5410 -739
rect 5376 -773 5410 -765
rect 5376 -833 5410 -811
rect 5376 -845 5410 -833
rect 5376 -901 5410 -883
rect 5376 -917 5410 -901
rect 5376 -969 5410 -955
rect 5376 -989 5410 -969
rect 5376 -1037 5410 -1027
rect 5376 -1061 5410 -1037
rect 5376 -1105 5410 -1099
rect 5376 -1133 5410 -1105
rect 5376 -1173 5410 -1171
rect 5376 -1205 5410 -1173
rect 5376 -1275 5410 -1243
rect 5376 -1277 5410 -1275
rect 5376 -1343 5410 -1315
rect 5376 -1349 5410 -1343
rect 5376 -1411 5410 -1387
rect 5376 -1421 5410 -1411
rect 5376 -1479 5410 -1459
rect 5376 -1493 5410 -1479
rect 5376 -1547 5410 -1531
rect 5376 -1565 5410 -1547
rect 5376 -1615 5410 -1603
rect 5376 -1637 5410 -1615
rect 5376 -1683 5410 -1675
rect 5376 -1709 5410 -1683
rect 5376 -1751 5410 -1747
rect 5376 -1781 5410 -1751
rect 5376 -1853 5410 -1819
rect 5376 -1921 5410 -1891
rect 5376 -1925 5410 -1921
rect 5376 -1989 5410 -1963
rect 5376 -1997 5410 -1989
rect 5376 -2057 5410 -2035
rect 5376 -2069 5410 -2057
rect 5376 -2125 5410 -2107
rect 5376 -2141 5410 -2125
rect 5376 -2193 5410 -2179
rect 5376 -2213 5410 -2193
rect 5376 -2261 5410 -2251
rect 5376 -2285 5410 -2261
rect 5376 -2329 5410 -2323
rect 5376 -2357 5410 -2329
rect 5376 -2397 5410 -2395
rect 5376 -2429 5410 -2397
rect 5376 -2499 5410 -2467
rect -5410 -2567 -5376 -2539
rect -5410 -2573 -5376 -2567
rect -5410 -2635 -5376 -2611
rect -5410 -2645 -5376 -2635
rect -5410 -2703 -5376 -2683
rect -5410 -2717 -5376 -2703
rect 5376 -2501 5410 -2499
rect 5376 -2567 5410 -2539
rect 5376 -2573 5410 -2567
rect 5376 -2635 5410 -2611
rect 5376 -2645 5410 -2635
rect 5376 -2703 5410 -2683
rect 5376 -2717 5410 -2703
rect -4805 -3062 -4777 -3028
rect -4777 -3062 -4771 -3028
rect -4733 -3062 -4709 -3028
rect -4709 -3062 -4699 -3028
rect -4661 -3062 -4641 -3028
rect -4641 -3062 -4627 -3028
rect -4589 -3062 -4573 -3028
rect -4573 -3062 -4555 -3028
rect -4517 -3062 -4505 -3028
rect -4505 -3062 -4483 -3028
rect -4445 -3062 -4437 -3028
rect -4437 -3062 -4411 -3028
rect -4373 -3062 -4369 -3028
rect -4369 -3062 -4339 -3028
rect -4301 -3062 -4267 -3028
rect -4229 -3062 -4199 -3028
rect -4199 -3062 -4195 -3028
rect -4157 -3062 -4131 -3028
rect -4131 -3062 -4123 -3028
rect -4085 -3062 -4063 -3028
rect -4063 -3062 -4051 -3028
rect -4013 -3062 -3995 -3028
rect -3995 -3062 -3979 -3028
rect -3941 -3062 -3927 -3028
rect -3927 -3062 -3907 -3028
rect -3869 -3062 -3859 -3028
rect -3859 -3062 -3835 -3028
rect -3797 -3062 -3791 -3028
rect -3791 -3062 -3763 -3028
rect -3725 -3062 -3723 -3028
rect -3723 -3062 -3691 -3028
rect -3653 -3062 -3621 -3028
rect -3621 -3062 -3619 -3028
rect -3581 -3062 -3553 -3028
rect -3553 -3062 -3547 -3028
rect -3509 -3062 -3485 -3028
rect -3485 -3062 -3475 -3028
rect -3437 -3062 -3417 -3028
rect -3417 -3062 -3403 -3028
rect -3365 -3062 -3349 -3028
rect -3349 -3062 -3331 -3028
rect -3293 -3062 -3281 -3028
rect -3281 -3062 -3259 -3028
rect -3221 -3062 -3213 -3028
rect -3213 -3062 -3187 -3028
rect -3149 -3062 -3145 -3028
rect -3145 -3062 -3115 -3028
rect -3077 -3062 -3043 -3028
rect -3005 -3062 -2975 -3028
rect -2975 -3062 -2971 -3028
rect -2933 -3062 -2907 -3028
rect -2907 -3062 -2899 -3028
rect -2861 -3062 -2839 -3028
rect -2839 -3062 -2827 -3028
rect -2789 -3062 -2771 -3028
rect -2771 -3062 -2755 -3028
rect -2717 -3062 -2703 -3028
rect -2703 -3062 -2683 -3028
rect -2645 -3062 -2635 -3028
rect -2635 -3062 -2611 -3028
rect -2573 -3062 -2567 -3028
rect -2567 -3062 -2539 -3028
rect -2501 -3062 -2499 -3028
rect -2499 -3062 -2467 -3028
rect -2429 -3062 -2397 -3028
rect -2397 -3062 -2395 -3028
rect -2357 -3062 -2329 -3028
rect -2329 -3062 -2323 -3028
rect -2285 -3062 -2261 -3028
rect -2261 -3062 -2251 -3028
rect -2213 -3062 -2193 -3028
rect -2193 -3062 -2179 -3028
rect -2141 -3062 -2125 -3028
rect -2125 -3062 -2107 -3028
rect -2069 -3062 -2057 -3028
rect -2057 -3062 -2035 -3028
rect -1997 -3062 -1989 -3028
rect -1989 -3062 -1963 -3028
rect -1925 -3062 -1921 -3028
rect -1921 -3062 -1891 -3028
rect -1853 -3062 -1819 -3028
rect -1781 -3062 -1751 -3028
rect -1751 -3062 -1747 -3028
rect -1709 -3062 -1683 -3028
rect -1683 -3062 -1675 -3028
rect -1637 -3062 -1615 -3028
rect -1615 -3062 -1603 -3028
rect -1565 -3062 -1547 -3028
rect -1547 -3062 -1531 -3028
rect -1493 -3062 -1479 -3028
rect -1479 -3062 -1459 -3028
rect -1421 -3062 -1411 -3028
rect -1411 -3062 -1387 -3028
rect -1349 -3062 -1343 -3028
rect -1343 -3062 -1315 -3028
rect -1277 -3062 -1275 -3028
rect -1275 -3062 -1243 -3028
rect -1205 -3062 -1173 -3028
rect -1173 -3062 -1171 -3028
rect -1133 -3062 -1105 -3028
rect -1105 -3062 -1099 -3028
rect -1061 -3062 -1037 -3028
rect -1037 -3062 -1027 -3028
rect -989 -3062 -969 -3028
rect -969 -3062 -955 -3028
rect -917 -3062 -901 -3028
rect -901 -3062 -883 -3028
rect -845 -3062 -833 -3028
rect -833 -3062 -811 -3028
rect -773 -3062 -765 -3028
rect -765 -3062 -739 -3028
rect -701 -3062 -697 -3028
rect -697 -3062 -667 -3028
rect -629 -3062 -595 -3028
rect -557 -3062 -527 -3028
rect -527 -3062 -523 -3028
rect -485 -3062 -459 -3028
rect -459 -3062 -451 -3028
rect -413 -3062 -391 -3028
rect -391 -3062 -379 -3028
rect -341 -3062 -323 -3028
rect -323 -3062 -307 -3028
rect -269 -3062 -255 -3028
rect -255 -3062 -235 -3028
rect -197 -3062 -187 -3028
rect -187 -3062 -163 -3028
rect -125 -3062 -119 -3028
rect -119 -3062 -91 -3028
rect -53 -3062 -51 -3028
rect -51 -3062 -19 -3028
rect 19 -3062 51 -3028
rect 51 -3062 53 -3028
rect 91 -3062 119 -3028
rect 119 -3062 125 -3028
rect 163 -3062 187 -3028
rect 187 -3062 197 -3028
rect 235 -3062 255 -3028
rect 255 -3062 269 -3028
rect 307 -3062 323 -3028
rect 323 -3062 341 -3028
rect 379 -3062 391 -3028
rect 391 -3062 413 -3028
rect 451 -3062 459 -3028
rect 459 -3062 485 -3028
rect 523 -3062 527 -3028
rect 527 -3062 557 -3028
rect 595 -3062 629 -3028
rect 667 -3062 697 -3028
rect 697 -3062 701 -3028
rect 739 -3062 765 -3028
rect 765 -3062 773 -3028
rect 811 -3062 833 -3028
rect 833 -3062 845 -3028
rect 883 -3062 901 -3028
rect 901 -3062 917 -3028
rect 955 -3062 969 -3028
rect 969 -3062 989 -3028
rect 1027 -3062 1037 -3028
rect 1037 -3062 1061 -3028
rect 1099 -3062 1105 -3028
rect 1105 -3062 1133 -3028
rect 1171 -3062 1173 -3028
rect 1173 -3062 1205 -3028
rect 1243 -3062 1275 -3028
rect 1275 -3062 1277 -3028
rect 1315 -3062 1343 -3028
rect 1343 -3062 1349 -3028
rect 1387 -3062 1411 -3028
rect 1411 -3062 1421 -3028
rect 1459 -3062 1479 -3028
rect 1479 -3062 1493 -3028
rect 1531 -3062 1547 -3028
rect 1547 -3062 1565 -3028
rect 1603 -3062 1615 -3028
rect 1615 -3062 1637 -3028
rect 1675 -3062 1683 -3028
rect 1683 -3062 1709 -3028
rect 1747 -3062 1751 -3028
rect 1751 -3062 1781 -3028
rect 1819 -3062 1853 -3028
rect 1891 -3062 1921 -3028
rect 1921 -3062 1925 -3028
rect 1963 -3062 1989 -3028
rect 1989 -3062 1997 -3028
rect 2035 -3062 2057 -3028
rect 2057 -3062 2069 -3028
rect 2107 -3062 2125 -3028
rect 2125 -3062 2141 -3028
rect 2179 -3062 2193 -3028
rect 2193 -3062 2213 -3028
rect 2251 -3062 2261 -3028
rect 2261 -3062 2285 -3028
rect 2323 -3062 2329 -3028
rect 2329 -3062 2357 -3028
rect 2395 -3062 2397 -3028
rect 2397 -3062 2429 -3028
rect 2467 -3062 2499 -3028
rect 2499 -3062 2501 -3028
rect 2539 -3062 2567 -3028
rect 2567 -3062 2573 -3028
rect 2611 -3062 2635 -3028
rect 2635 -3062 2645 -3028
rect 2683 -3062 2703 -3028
rect 2703 -3062 2717 -3028
rect 2755 -3062 2771 -3028
rect 2771 -3062 2789 -3028
rect 2827 -3062 2839 -3028
rect 2839 -3062 2861 -3028
rect 2899 -3062 2907 -3028
rect 2907 -3062 2933 -3028
rect 2971 -3062 2975 -3028
rect 2975 -3062 3005 -3028
rect 3043 -3062 3077 -3028
rect 3115 -3062 3145 -3028
rect 3145 -3062 3149 -3028
rect 3187 -3062 3213 -3028
rect 3213 -3062 3221 -3028
rect 3259 -3062 3281 -3028
rect 3281 -3062 3293 -3028
rect 3331 -3062 3349 -3028
rect 3349 -3062 3365 -3028
rect 3403 -3062 3417 -3028
rect 3417 -3062 3437 -3028
rect 3475 -3062 3485 -3028
rect 3485 -3062 3509 -3028
rect 3547 -3062 3553 -3028
rect 3553 -3062 3581 -3028
rect 3619 -3062 3621 -3028
rect 3621 -3062 3653 -3028
rect 3691 -3062 3723 -3028
rect 3723 -3062 3725 -3028
rect 3763 -3062 3791 -3028
rect 3791 -3062 3797 -3028
rect 3835 -3062 3859 -3028
rect 3859 -3062 3869 -3028
rect 3907 -3062 3927 -3028
rect 3927 -3062 3941 -3028
rect 3979 -3062 3995 -3028
rect 3995 -3062 4013 -3028
rect 4051 -3062 4063 -3028
rect 4063 -3062 4085 -3028
rect 4123 -3062 4131 -3028
rect 4131 -3062 4157 -3028
rect 4195 -3062 4199 -3028
rect 4199 -3062 4229 -3028
rect 4267 -3062 4301 -3028
rect 4339 -3062 4369 -3028
rect 4369 -3062 4373 -3028
rect 4411 -3062 4437 -3028
rect 4437 -3062 4445 -3028
rect 4483 -3062 4505 -3028
rect 4505 -3062 4517 -3028
rect 4555 -3062 4573 -3028
rect 4573 -3062 4589 -3028
rect 4627 -3062 4641 -3028
rect 4641 -3062 4661 -3028
rect 4699 -3062 4709 -3028
rect 4709 -3062 4733 -3028
rect 4771 -3062 4777 -3028
rect 4777 -3062 4805 -3028
<< metal1 >>
rect -5416 2717 -5370 2737
rect -5416 2683 -5410 2717
rect -5376 2683 -5370 2717
rect -5416 2645 -5370 2683
rect -5416 2611 -5410 2645
rect -5376 2611 -5370 2645
rect -5416 2573 -5370 2611
rect -5416 2539 -5410 2573
rect -5376 2539 -5370 2573
rect -5416 2501 -5370 2539
rect -5416 2467 -5410 2501
rect -5376 2467 -5370 2501
rect -5416 2429 -5370 2467
rect -5416 2395 -5410 2429
rect -5376 2395 -5370 2429
rect -5416 2357 -5370 2395
rect -5416 2323 -5410 2357
rect -5376 2323 -5370 2357
rect -5416 2285 -5370 2323
rect -5416 2251 -5410 2285
rect -5376 2251 -5370 2285
rect -5416 2213 -5370 2251
rect -5416 2179 -5410 2213
rect -5376 2179 -5370 2213
rect -5416 2141 -5370 2179
rect -5416 2107 -5410 2141
rect -5376 2107 -5370 2141
rect -5416 2069 -5370 2107
rect -5416 2035 -5410 2069
rect -5376 2035 -5370 2069
rect -5416 1997 -5370 2035
rect -5416 1963 -5410 1997
rect -5376 1963 -5370 1997
rect -5416 1925 -5370 1963
rect -5416 1891 -5410 1925
rect -5376 1891 -5370 1925
rect -5416 1853 -5370 1891
rect -5416 1819 -5410 1853
rect -5376 1819 -5370 1853
rect -5416 1781 -5370 1819
rect -5416 1747 -5410 1781
rect -5376 1747 -5370 1781
rect -5416 1709 -5370 1747
rect -5416 1675 -5410 1709
rect -5376 1675 -5370 1709
rect -5416 1637 -5370 1675
rect -5416 1603 -5410 1637
rect -5376 1603 -5370 1637
rect -5416 1565 -5370 1603
rect -5416 1531 -5410 1565
rect -5376 1531 -5370 1565
rect -5416 1493 -5370 1531
rect -5416 1459 -5410 1493
rect -5376 1459 -5370 1493
rect -5416 1421 -5370 1459
rect -5416 1387 -5410 1421
rect -5376 1387 -5370 1421
rect -5416 1349 -5370 1387
rect -5416 1315 -5410 1349
rect -5376 1315 -5370 1349
rect -5416 1277 -5370 1315
rect -5416 1243 -5410 1277
rect -5376 1243 -5370 1277
rect -5416 1205 -5370 1243
rect -5416 1171 -5410 1205
rect -5376 1171 -5370 1205
rect -5416 1133 -5370 1171
rect -5416 1099 -5410 1133
rect -5376 1099 -5370 1133
rect -5416 1061 -5370 1099
rect -5416 1027 -5410 1061
rect -5376 1027 -5370 1061
rect -5416 989 -5370 1027
rect -5416 955 -5410 989
rect -5376 955 -5370 989
rect -5416 917 -5370 955
rect -5416 883 -5410 917
rect -5376 883 -5370 917
rect -5416 845 -5370 883
rect -5416 811 -5410 845
rect -5376 811 -5370 845
rect -5416 773 -5370 811
rect -5416 739 -5410 773
rect -5376 739 -5370 773
rect -5416 701 -5370 739
rect -5416 667 -5410 701
rect -5376 667 -5370 701
rect -5416 629 -5370 667
rect -5416 595 -5410 629
rect -5376 595 -5370 629
rect -5416 557 -5370 595
rect -5416 523 -5410 557
rect -5376 523 -5370 557
rect -5416 485 -5370 523
rect -5416 451 -5410 485
rect -5376 451 -5370 485
rect -5416 413 -5370 451
rect -5416 379 -5410 413
rect -5376 379 -5370 413
rect -5416 341 -5370 379
rect -5416 307 -5410 341
rect -5376 307 -5370 341
rect -5416 269 -5370 307
rect -5416 235 -5410 269
rect -5376 235 -5370 269
rect -5416 197 -5370 235
rect -5416 163 -5410 197
rect -5376 163 -5370 197
rect -5416 125 -5370 163
rect -5416 91 -5410 125
rect -5376 91 -5370 125
rect -5416 53 -5370 91
rect -5416 19 -5410 53
rect -5376 19 -5370 53
rect -5416 -19 -5370 19
rect -5416 -53 -5410 -19
rect -5376 -53 -5370 -19
rect -5416 -91 -5370 -53
rect -5416 -125 -5410 -91
rect -5376 -125 -5370 -91
rect -5416 -163 -5370 -125
rect -5416 -197 -5410 -163
rect -5376 -197 -5370 -163
rect -5416 -235 -5370 -197
rect -5416 -269 -5410 -235
rect -5376 -269 -5370 -235
rect -5416 -307 -5370 -269
rect -5416 -341 -5410 -307
rect -5376 -341 -5370 -307
rect -5416 -379 -5370 -341
rect -5416 -413 -5410 -379
rect -5376 -413 -5370 -379
rect -5416 -451 -5370 -413
rect -5416 -485 -5410 -451
rect -5376 -485 -5370 -451
rect -5416 -523 -5370 -485
rect -5416 -557 -5410 -523
rect -5376 -557 -5370 -523
rect -5416 -595 -5370 -557
rect -5416 -629 -5410 -595
rect -5376 -629 -5370 -595
rect -5416 -667 -5370 -629
rect -5416 -701 -5410 -667
rect -5376 -701 -5370 -667
rect -5416 -739 -5370 -701
rect -5416 -773 -5410 -739
rect -5376 -773 -5370 -739
rect -5416 -811 -5370 -773
rect -5416 -845 -5410 -811
rect -5376 -845 -5370 -811
rect -5416 -883 -5370 -845
rect -5416 -917 -5410 -883
rect -5376 -917 -5370 -883
rect -5416 -955 -5370 -917
rect -5416 -989 -5410 -955
rect -5376 -989 -5370 -955
rect -5416 -1027 -5370 -989
rect -5416 -1061 -5410 -1027
rect -5376 -1061 -5370 -1027
rect -5416 -1099 -5370 -1061
rect -5416 -1133 -5410 -1099
rect -5376 -1133 -5370 -1099
rect -5416 -1171 -5370 -1133
rect -5416 -1205 -5410 -1171
rect -5376 -1205 -5370 -1171
rect -5416 -1243 -5370 -1205
rect -5416 -1277 -5410 -1243
rect -5376 -1277 -5370 -1243
rect -5416 -1315 -5370 -1277
rect -5416 -1349 -5410 -1315
rect -5376 -1349 -5370 -1315
rect -5416 -1387 -5370 -1349
rect -5416 -1421 -5410 -1387
rect -5376 -1421 -5370 -1387
rect -5416 -1459 -5370 -1421
rect -5416 -1493 -5410 -1459
rect -5376 -1493 -5370 -1459
rect -5416 -1531 -5370 -1493
rect -5416 -1565 -5410 -1531
rect -5376 -1565 -5370 -1531
rect -5416 -1603 -5370 -1565
rect -5416 -1637 -5410 -1603
rect -5376 -1637 -5370 -1603
rect -5416 -1675 -5370 -1637
rect -5416 -1709 -5410 -1675
rect -5376 -1709 -5370 -1675
rect -5416 -1747 -5370 -1709
rect -5416 -1781 -5410 -1747
rect -5376 -1781 -5370 -1747
rect -5416 -1819 -5370 -1781
rect -5416 -1853 -5410 -1819
rect -5376 -1853 -5370 -1819
rect -5416 -1891 -5370 -1853
rect -5416 -1925 -5410 -1891
rect -5376 -1925 -5370 -1891
rect -5416 -1963 -5370 -1925
rect -5416 -1997 -5410 -1963
rect -5376 -1997 -5370 -1963
rect -5416 -2035 -5370 -1997
rect -5416 -2069 -5410 -2035
rect -5376 -2069 -5370 -2035
rect -5416 -2107 -5370 -2069
rect -5416 -2141 -5410 -2107
rect -5376 -2141 -5370 -2107
rect -5416 -2179 -5370 -2141
rect -5416 -2213 -5410 -2179
rect -5376 -2213 -5370 -2179
rect -5416 -2251 -5370 -2213
rect -5416 -2285 -5410 -2251
rect -5376 -2285 -5370 -2251
rect -5416 -2323 -5370 -2285
rect -5416 -2357 -5410 -2323
rect -5376 -2357 -5370 -2323
rect -5416 -2395 -5370 -2357
rect -5416 -2429 -5410 -2395
rect -5376 -2429 -5370 -2395
rect -5416 -2467 -5370 -2429
rect -5416 -2501 -5410 -2467
rect -5376 -2501 -5370 -2467
rect -5416 -2539 -5370 -2501
rect -5416 -2573 -5410 -2539
rect -5376 -2573 -5370 -2539
rect -5416 -2611 -5370 -2573
rect -5416 -2645 -5410 -2611
rect -5376 -2645 -5370 -2611
rect -5416 -2683 -5370 -2645
rect -5416 -2717 -5410 -2683
rect -5376 -2717 -5370 -2683
rect -5416 -2737 -5370 -2717
rect 5370 2717 5416 2737
rect 5370 2683 5376 2717
rect 5410 2683 5416 2717
rect 5370 2645 5416 2683
rect 5370 2611 5376 2645
rect 5410 2611 5416 2645
rect 5370 2573 5416 2611
rect 5370 2539 5376 2573
rect 5410 2539 5416 2573
rect 5370 2501 5416 2539
rect 5370 2467 5376 2501
rect 5410 2467 5416 2501
rect 5370 2429 5416 2467
rect 5370 2395 5376 2429
rect 5410 2395 5416 2429
rect 5370 2357 5416 2395
rect 5370 2323 5376 2357
rect 5410 2323 5416 2357
rect 5370 2285 5416 2323
rect 5370 2251 5376 2285
rect 5410 2251 5416 2285
rect 5370 2213 5416 2251
rect 5370 2179 5376 2213
rect 5410 2179 5416 2213
rect 5370 2141 5416 2179
rect 5370 2107 5376 2141
rect 5410 2107 5416 2141
rect 5370 2069 5416 2107
rect 5370 2035 5376 2069
rect 5410 2035 5416 2069
rect 5370 1997 5416 2035
rect 5370 1963 5376 1997
rect 5410 1963 5416 1997
rect 5370 1925 5416 1963
rect 5370 1891 5376 1925
rect 5410 1891 5416 1925
rect 5370 1853 5416 1891
rect 5370 1819 5376 1853
rect 5410 1819 5416 1853
rect 5370 1781 5416 1819
rect 5370 1747 5376 1781
rect 5410 1747 5416 1781
rect 5370 1709 5416 1747
rect 5370 1675 5376 1709
rect 5410 1675 5416 1709
rect 5370 1637 5416 1675
rect 5370 1603 5376 1637
rect 5410 1603 5416 1637
rect 5370 1565 5416 1603
rect 5370 1531 5376 1565
rect 5410 1531 5416 1565
rect 5370 1493 5416 1531
rect 5370 1459 5376 1493
rect 5410 1459 5416 1493
rect 5370 1421 5416 1459
rect 5370 1387 5376 1421
rect 5410 1387 5416 1421
rect 5370 1349 5416 1387
rect 5370 1315 5376 1349
rect 5410 1315 5416 1349
rect 5370 1277 5416 1315
rect 5370 1243 5376 1277
rect 5410 1243 5416 1277
rect 5370 1205 5416 1243
rect 5370 1171 5376 1205
rect 5410 1171 5416 1205
rect 5370 1133 5416 1171
rect 5370 1099 5376 1133
rect 5410 1099 5416 1133
rect 5370 1061 5416 1099
rect 5370 1027 5376 1061
rect 5410 1027 5416 1061
rect 5370 989 5416 1027
rect 5370 955 5376 989
rect 5410 955 5416 989
rect 5370 917 5416 955
rect 5370 883 5376 917
rect 5410 883 5416 917
rect 5370 845 5416 883
rect 5370 811 5376 845
rect 5410 811 5416 845
rect 5370 773 5416 811
rect 5370 739 5376 773
rect 5410 739 5416 773
rect 5370 701 5416 739
rect 5370 667 5376 701
rect 5410 667 5416 701
rect 5370 629 5416 667
rect 5370 595 5376 629
rect 5410 595 5416 629
rect 5370 557 5416 595
rect 5370 523 5376 557
rect 5410 523 5416 557
rect 5370 485 5416 523
rect 5370 451 5376 485
rect 5410 451 5416 485
rect 5370 413 5416 451
rect 5370 379 5376 413
rect 5410 379 5416 413
rect 5370 341 5416 379
rect 5370 307 5376 341
rect 5410 307 5416 341
rect 5370 269 5416 307
rect 5370 235 5376 269
rect 5410 235 5416 269
rect 5370 197 5416 235
rect 5370 163 5376 197
rect 5410 163 5416 197
rect 5370 125 5416 163
rect 5370 91 5376 125
rect 5410 91 5416 125
rect 5370 53 5416 91
rect 5370 19 5376 53
rect 5410 19 5416 53
rect 5370 -19 5416 19
rect 5370 -53 5376 -19
rect 5410 -53 5416 -19
rect 5370 -91 5416 -53
rect 5370 -125 5376 -91
rect 5410 -125 5416 -91
rect 5370 -163 5416 -125
rect 5370 -197 5376 -163
rect 5410 -197 5416 -163
rect 5370 -235 5416 -197
rect 5370 -269 5376 -235
rect 5410 -269 5416 -235
rect 5370 -307 5416 -269
rect 5370 -341 5376 -307
rect 5410 -341 5416 -307
rect 5370 -379 5416 -341
rect 5370 -413 5376 -379
rect 5410 -413 5416 -379
rect 5370 -451 5416 -413
rect 5370 -485 5376 -451
rect 5410 -485 5416 -451
rect 5370 -523 5416 -485
rect 5370 -557 5376 -523
rect 5410 -557 5416 -523
rect 5370 -595 5416 -557
rect 5370 -629 5376 -595
rect 5410 -629 5416 -595
rect 5370 -667 5416 -629
rect 5370 -701 5376 -667
rect 5410 -701 5416 -667
rect 5370 -739 5416 -701
rect 5370 -773 5376 -739
rect 5410 -773 5416 -739
rect 5370 -811 5416 -773
rect 5370 -845 5376 -811
rect 5410 -845 5416 -811
rect 5370 -883 5416 -845
rect 5370 -917 5376 -883
rect 5410 -917 5416 -883
rect 5370 -955 5416 -917
rect 5370 -989 5376 -955
rect 5410 -989 5416 -955
rect 5370 -1027 5416 -989
rect 5370 -1061 5376 -1027
rect 5410 -1061 5416 -1027
rect 5370 -1099 5416 -1061
rect 5370 -1133 5376 -1099
rect 5410 -1133 5416 -1099
rect 5370 -1171 5416 -1133
rect 5370 -1205 5376 -1171
rect 5410 -1205 5416 -1171
rect 5370 -1243 5416 -1205
rect 5370 -1277 5376 -1243
rect 5410 -1277 5416 -1243
rect 5370 -1315 5416 -1277
rect 5370 -1349 5376 -1315
rect 5410 -1349 5416 -1315
rect 5370 -1387 5416 -1349
rect 5370 -1421 5376 -1387
rect 5410 -1421 5416 -1387
rect 5370 -1459 5416 -1421
rect 5370 -1493 5376 -1459
rect 5410 -1493 5416 -1459
rect 5370 -1531 5416 -1493
rect 5370 -1565 5376 -1531
rect 5410 -1565 5416 -1531
rect 5370 -1603 5416 -1565
rect 5370 -1637 5376 -1603
rect 5410 -1637 5416 -1603
rect 5370 -1675 5416 -1637
rect 5370 -1709 5376 -1675
rect 5410 -1709 5416 -1675
rect 5370 -1747 5416 -1709
rect 5370 -1781 5376 -1747
rect 5410 -1781 5416 -1747
rect 5370 -1819 5416 -1781
rect 5370 -1853 5376 -1819
rect 5410 -1853 5416 -1819
rect 5370 -1891 5416 -1853
rect 5370 -1925 5376 -1891
rect 5410 -1925 5416 -1891
rect 5370 -1963 5416 -1925
rect 5370 -1997 5376 -1963
rect 5410 -1997 5416 -1963
rect 5370 -2035 5416 -1997
rect 5370 -2069 5376 -2035
rect 5410 -2069 5416 -2035
rect 5370 -2107 5416 -2069
rect 5370 -2141 5376 -2107
rect 5410 -2141 5416 -2107
rect 5370 -2179 5416 -2141
rect 5370 -2213 5376 -2179
rect 5410 -2213 5416 -2179
rect 5370 -2251 5416 -2213
rect 5370 -2285 5376 -2251
rect 5410 -2285 5416 -2251
rect 5370 -2323 5416 -2285
rect 5370 -2357 5376 -2323
rect 5410 -2357 5416 -2323
rect 5370 -2395 5416 -2357
rect 5370 -2429 5376 -2395
rect 5410 -2429 5416 -2395
rect 5370 -2467 5416 -2429
rect 5370 -2501 5376 -2467
rect 5410 -2501 5416 -2467
rect 5370 -2539 5416 -2501
rect 5370 -2573 5376 -2539
rect 5410 -2573 5416 -2539
rect 5370 -2611 5416 -2573
rect 5370 -2645 5376 -2611
rect 5410 -2645 5416 -2611
rect 5370 -2683 5416 -2645
rect 5370 -2717 5376 -2683
rect 5410 -2717 5416 -2683
rect 5370 -2737 5416 -2717
rect -4850 -3028 4850 -3022
rect -4850 -3062 -4805 -3028
rect -4771 -3062 -4733 -3028
rect -4699 -3062 -4661 -3028
rect -4627 -3062 -4589 -3028
rect -4555 -3062 -4517 -3028
rect -4483 -3062 -4445 -3028
rect -4411 -3062 -4373 -3028
rect -4339 -3062 -4301 -3028
rect -4267 -3062 -4229 -3028
rect -4195 -3062 -4157 -3028
rect -4123 -3062 -4085 -3028
rect -4051 -3062 -4013 -3028
rect -3979 -3062 -3941 -3028
rect -3907 -3062 -3869 -3028
rect -3835 -3062 -3797 -3028
rect -3763 -3062 -3725 -3028
rect -3691 -3062 -3653 -3028
rect -3619 -3062 -3581 -3028
rect -3547 -3062 -3509 -3028
rect -3475 -3062 -3437 -3028
rect -3403 -3062 -3365 -3028
rect -3331 -3062 -3293 -3028
rect -3259 -3062 -3221 -3028
rect -3187 -3062 -3149 -3028
rect -3115 -3062 -3077 -3028
rect -3043 -3062 -3005 -3028
rect -2971 -3062 -2933 -3028
rect -2899 -3062 -2861 -3028
rect -2827 -3062 -2789 -3028
rect -2755 -3062 -2717 -3028
rect -2683 -3062 -2645 -3028
rect -2611 -3062 -2573 -3028
rect -2539 -3062 -2501 -3028
rect -2467 -3062 -2429 -3028
rect -2395 -3062 -2357 -3028
rect -2323 -3062 -2285 -3028
rect -2251 -3062 -2213 -3028
rect -2179 -3062 -2141 -3028
rect -2107 -3062 -2069 -3028
rect -2035 -3062 -1997 -3028
rect -1963 -3062 -1925 -3028
rect -1891 -3062 -1853 -3028
rect -1819 -3062 -1781 -3028
rect -1747 -3062 -1709 -3028
rect -1675 -3062 -1637 -3028
rect -1603 -3062 -1565 -3028
rect -1531 -3062 -1493 -3028
rect -1459 -3062 -1421 -3028
rect -1387 -3062 -1349 -3028
rect -1315 -3062 -1277 -3028
rect -1243 -3062 -1205 -3028
rect -1171 -3062 -1133 -3028
rect -1099 -3062 -1061 -3028
rect -1027 -3062 -989 -3028
rect -955 -3062 -917 -3028
rect -883 -3062 -845 -3028
rect -811 -3062 -773 -3028
rect -739 -3062 -701 -3028
rect -667 -3062 -629 -3028
rect -595 -3062 -557 -3028
rect -523 -3062 -485 -3028
rect -451 -3062 -413 -3028
rect -379 -3062 -341 -3028
rect -307 -3062 -269 -3028
rect -235 -3062 -197 -3028
rect -163 -3062 -125 -3028
rect -91 -3062 -53 -3028
rect -19 -3062 19 -3028
rect 53 -3062 91 -3028
rect 125 -3062 163 -3028
rect 197 -3062 235 -3028
rect 269 -3062 307 -3028
rect 341 -3062 379 -3028
rect 413 -3062 451 -3028
rect 485 -3062 523 -3028
rect 557 -3062 595 -3028
rect 629 -3062 667 -3028
rect 701 -3062 739 -3028
rect 773 -3062 811 -3028
rect 845 -3062 883 -3028
rect 917 -3062 955 -3028
rect 989 -3062 1027 -3028
rect 1061 -3062 1099 -3028
rect 1133 -3062 1171 -3028
rect 1205 -3062 1243 -3028
rect 1277 -3062 1315 -3028
rect 1349 -3062 1387 -3028
rect 1421 -3062 1459 -3028
rect 1493 -3062 1531 -3028
rect 1565 -3062 1603 -3028
rect 1637 -3062 1675 -3028
rect 1709 -3062 1747 -3028
rect 1781 -3062 1819 -3028
rect 1853 -3062 1891 -3028
rect 1925 -3062 1963 -3028
rect 1997 -3062 2035 -3028
rect 2069 -3062 2107 -3028
rect 2141 -3062 2179 -3028
rect 2213 -3062 2251 -3028
rect 2285 -3062 2323 -3028
rect 2357 -3062 2395 -3028
rect 2429 -3062 2467 -3028
rect 2501 -3062 2539 -3028
rect 2573 -3062 2611 -3028
rect 2645 -3062 2683 -3028
rect 2717 -3062 2755 -3028
rect 2789 -3062 2827 -3028
rect 2861 -3062 2899 -3028
rect 2933 -3062 2971 -3028
rect 3005 -3062 3043 -3028
rect 3077 -3062 3115 -3028
rect 3149 -3062 3187 -3028
rect 3221 -3062 3259 -3028
rect 3293 -3062 3331 -3028
rect 3365 -3062 3403 -3028
rect 3437 -3062 3475 -3028
rect 3509 -3062 3547 -3028
rect 3581 -3062 3619 -3028
rect 3653 -3062 3691 -3028
rect 3725 -3062 3763 -3028
rect 3797 -3062 3835 -3028
rect 3869 -3062 3907 -3028
rect 3941 -3062 3979 -3028
rect 4013 -3062 4051 -3028
rect 4085 -3062 4123 -3028
rect 4157 -3062 4195 -3028
rect 4229 -3062 4267 -3028
rect 4301 -3062 4339 -3028
rect 4373 -3062 4411 -3028
rect 4445 -3062 4483 -3028
rect 4517 -3062 4555 -3028
rect 4589 -3062 4627 -3028
rect 4661 -3062 4699 -3028
rect 4733 -3062 4771 -3028
rect 4805 -3062 4850 -3028
rect -4850 -3068 4850 -3062
<< properties >>
string FIXED_BBOX -5393 -3045 5393 3045
<< end >>
