magic
tech sky130A
magscale 1 2
timestamp 1683391037
<< nwell >>
rect -941 -719 941 719
<< pmos >>
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
<< pdiff >>
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
<< pdiffc >>
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
<< nsubdiff >>
rect -905 649 -809 683
rect 809 649 905 683
rect -905 587 -871 649
rect 871 587 905 649
rect -905 -649 -871 -587
rect 871 -649 905 -587
rect -905 -683 -809 -649
rect 809 -683 905 -649
<< nsubdiffcont >>
rect -809 649 809 683
rect -905 -587 -871 587
rect 871 -587 905 587
rect -809 -683 809 -649
<< poly >>
rect -745 581 -545 597
rect -745 547 -729 581
rect -561 547 -545 581
rect -745 500 -545 547
rect -487 581 -287 597
rect -487 547 -471 581
rect -303 547 -287 581
rect -487 500 -287 547
rect -229 581 -29 597
rect -229 547 -213 581
rect -45 547 -29 581
rect -229 500 -29 547
rect 29 581 229 597
rect 29 547 45 581
rect 213 547 229 581
rect 29 500 229 547
rect 287 581 487 597
rect 287 547 303 581
rect 471 547 487 581
rect 287 500 487 547
rect 545 581 745 597
rect 545 547 561 581
rect 729 547 745 581
rect 545 500 745 547
rect -745 -547 -545 -500
rect -745 -581 -729 -547
rect -561 -581 -545 -547
rect -745 -597 -545 -581
rect -487 -547 -287 -500
rect -487 -581 -471 -547
rect -303 -581 -287 -547
rect -487 -597 -287 -581
rect -229 -547 -29 -500
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect -229 -597 -29 -581
rect 29 -547 229 -500
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 29 -597 229 -581
rect 287 -547 487 -500
rect 287 -581 303 -547
rect 471 -581 487 -547
rect 287 -597 487 -581
rect 545 -547 745 -500
rect 545 -581 561 -547
rect 729 -581 745 -547
rect 545 -597 745 -581
<< polycont >>
rect -729 547 -561 581
rect -471 547 -303 581
rect -213 547 -45 581
rect 45 547 213 581
rect 303 547 471 581
rect 561 547 729 581
rect -729 -581 -561 -547
rect -471 -581 -303 -547
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect 303 -581 471 -547
rect 561 -581 729 -547
<< locali >>
rect -905 649 -809 683
rect 809 649 905 683
rect -905 587 -871 649
rect 871 587 905 649
rect -745 547 -729 581
rect -561 547 -545 581
rect -487 547 -471 581
rect -303 547 -287 581
rect -229 547 -213 581
rect -45 547 -29 581
rect 29 547 45 581
rect 213 547 229 581
rect 287 547 303 581
rect 471 547 487 581
rect 545 547 561 581
rect 729 547 745 581
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect -745 -581 -729 -547
rect -561 -581 -545 -547
rect -487 -581 -471 -547
rect -303 -581 -287 -547
rect -229 -581 -213 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 213 -581 229 -547
rect 287 -581 303 -547
rect 471 -581 487 -547
rect 545 -581 561 -547
rect 729 -581 745 -547
rect -905 -649 -871 -587
rect 871 -649 905 -587
rect -905 -683 -809 -649
rect 809 -683 905 -649
<< viali >>
rect -729 547 -561 581
rect -471 547 -303 581
rect -213 547 -45 581
rect 45 547 213 581
rect 303 547 471 581
rect 561 547 729 581
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect -729 -581 -561 -547
rect -471 -581 -303 -547
rect -213 -581 -45 -547
rect 45 -581 213 -547
rect 303 -581 471 -547
rect 561 -581 729 -547
<< metal1 >>
rect -741 581 -549 587
rect -741 547 -729 581
rect -561 547 -549 581
rect -741 541 -549 547
rect -483 581 -291 587
rect -483 547 -471 581
rect -303 547 -291 581
rect -483 541 -291 547
rect -225 581 -33 587
rect -225 547 -213 581
rect -45 547 -33 581
rect -225 541 -33 547
rect 33 581 225 587
rect 33 547 45 581
rect 213 547 225 581
rect 33 541 225 547
rect 291 581 483 587
rect 291 547 303 581
rect 471 547 483 581
rect 291 541 483 547
rect 549 581 741 587
rect 549 547 561 581
rect 729 547 741 581
rect 549 541 741 547
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect -741 -547 -549 -541
rect -741 -581 -729 -547
rect -561 -581 -549 -547
rect -741 -587 -549 -581
rect -483 -547 -291 -541
rect -483 -581 -471 -547
rect -303 -581 -291 -547
rect -483 -587 -291 -581
rect -225 -547 -33 -541
rect -225 -581 -213 -547
rect -45 -581 -33 -547
rect -225 -587 -33 -581
rect 33 -547 225 -541
rect 33 -581 45 -547
rect 213 -581 225 -547
rect 33 -587 225 -581
rect 291 -547 483 -541
rect 291 -581 303 -547
rect 471 -581 483 -547
rect 291 -587 483 -581
rect 549 -547 741 -541
rect 549 -581 561 -547
rect 729 -581 741 -547
rect 549 -587 741 -581
<< properties >>
string FIXED_BBOX -888 -666 888 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 1 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
