magic
tech sky130A
magscale 1 2
timestamp 1685420127
<< error_s >>
rect 37390 700890 37391 700891
rect 37389 700889 37390 700890
rect 37389 697770 37390 697771
rect 37390 697769 37391 697770
rect 41527 694199 41627 694200
rect 41685 694199 41785 694200
rect 41843 694199 41943 694200
rect 42001 694199 42101 694200
rect 42159 694199 42259 694200
rect 42317 694199 42417 694200
rect 42475 694199 42575 694200
rect 42633 694199 42733 694200
rect 42791 694199 42891 694200
rect 42949 694199 43049 694200
rect 43107 694199 43207 694200
rect 43265 694199 43365 694200
rect 43423 694199 43523 694200
rect 43581 694199 43681 694200
rect 43739 694199 43839 694200
rect 43897 694199 43997 694200
rect 44055 694199 44155 694200
rect 44213 694199 44313 694200
rect 44371 694199 44471 694200
rect 44529 694199 44629 694200
rect 44673 694195 44675 694320
rect 44685 694199 44785 694200
rect 44843 694199 44943 694200
rect 45001 694199 45101 694200
rect 45159 694199 45259 694200
rect 45317 694199 45417 694200
rect 45475 694199 45575 694200
rect 45633 694199 45733 694200
rect 45791 694199 45891 694200
rect 45949 694199 46049 694200
rect 46107 694199 46207 694200
rect 46265 694199 46365 694200
rect 46423 694199 46523 694200
rect 46581 694199 46681 694200
rect 46739 694199 46839 694200
rect 46897 694199 46997 694200
rect 47055 694199 47155 694200
rect 47213 694199 47313 694200
rect 47371 694199 47471 694200
rect 47529 694199 47629 694200
rect 47687 694199 47787 694200
rect 43042 693575 43110 693576
rect 43200 693575 43268 693576
rect 43358 693575 43426 693576
rect 43516 693575 43584 693576
rect 43674 693575 43742 693576
rect 43832 693575 43900 693576
rect 43990 693575 44058 693576
rect 44148 693575 44216 693576
rect 44306 693575 44374 693576
rect 44464 693575 44532 693576
rect 44622 693575 44690 693576
rect 44780 693575 44848 693576
rect 44938 693575 45006 693576
rect 45096 693575 45164 693576
rect 45254 693575 45322 693576
rect 45412 693575 45480 693576
rect 45570 693575 45638 693576
rect 45728 693575 45796 693576
rect 45886 693575 45954 693576
rect 46044 693575 46112 693576
rect 46202 693575 46270 693576
rect 43026 692529 43126 692530
rect 43184 692529 43284 692530
rect 43342 692529 43442 692530
rect 43500 692529 43600 692530
rect 43658 692529 43758 692530
rect 43816 692529 43916 692530
rect 43974 692529 44074 692530
rect 44132 692529 44232 692530
rect 44290 692529 44390 692530
rect 44448 692529 44548 692530
rect 44606 692529 44706 692530
rect 44764 692529 44864 692530
rect 44922 692529 45022 692530
rect 45080 692529 45180 692530
rect 45238 692529 45338 692530
rect 45396 692529 45496 692530
rect 45554 692529 45654 692530
rect 45712 692529 45812 692530
rect 45870 692529 45970 692530
rect 46028 692529 46128 692530
rect 46186 692529 46286 692530
rect 43042 692035 43110 692036
rect 43200 692035 43268 692036
rect 43358 692035 43426 692036
rect 43516 692035 43584 692036
rect 43674 692035 43742 692036
rect 43832 692035 43900 692036
rect 43990 692035 44058 692036
rect 44148 692035 44216 692036
rect 44306 692035 44374 692036
rect 44464 692035 44532 692036
rect 44622 692035 44690 692036
rect 44780 692035 44848 692036
rect 44938 692035 45006 692036
rect 45096 692035 45164 692036
rect 45254 692035 45322 692036
rect 45412 692035 45480 692036
rect 45570 692035 45638 692036
rect 45728 692035 45796 692036
rect 45886 692035 45954 692036
rect 46044 692035 46112 692036
rect 46202 692035 46270 692036
rect 43412 692029 43438 692030
rect 43440 692001 43466 692030
rect 43476 692001 43500 692030
rect 43504 692029 43528 692030
rect 43732 692029 43754 692030
rect 43760 692001 43782 692030
rect 45688 692001 45710 692030
rect 45716 692029 45738 692030
rect 45942 692029 45966 692030
rect 45970 692001 45994 692030
rect 46004 692001 46030 692030
rect 46032 692029 46058 692030
rect 43026 690989 43126 690990
rect 43184 690989 43284 690990
rect 43342 690989 43442 690990
rect 43500 690989 43600 690990
rect 43658 690989 43758 690990
rect 43816 690989 43916 690990
rect 43974 690989 44074 690990
rect 44132 690989 44232 690990
rect 44290 690989 44390 690990
rect 44448 690989 44548 690990
rect 44606 690989 44706 690990
rect 44764 690989 44864 690990
rect 44922 690989 45022 690990
rect 45080 690989 45180 690990
rect 45238 690989 45338 690990
rect 45396 690989 45496 690990
rect 45554 690989 45654 690990
rect 45712 690989 45812 690990
rect 45870 690989 45970 690990
rect 46028 690989 46128 690990
rect 46186 690989 46286 690990
rect 44669 684856 44671 685864
rect 44651 680206 44653 680714
rect 44649 679457 44651 679713
rect 44870 679710 44920 679737
rect 44867 679682 44913 679709
rect 44652 677956 44654 678964
<< nwell >>
rect 534289 289502 546909 294942
rect 536434 284239 544644 285480
rect 536794 284238 544412 284239
rect 12500 269330 17250 275990
rect 23960 271710 26900 273600
<< pwell >>
rect 541314 677258 547888 678108
rect 541312 663278 547884 664522
rect 5780 303200 16200 304514
rect 559800 295600 561114 306020
rect 569000 295600 570314 306020
rect 5780 292800 16200 294114
rect 530556 289189 533752 292137
rect 536249 288722 544977 289214
rect 547616 289189 550812 292137
rect 536249 288222 544977 288714
rect 536809 287622 544319 288214
rect 536809 287002 544319 287594
rect 568080 287580 578500 288894
rect 536249 286402 544977 286994
rect 536249 285802 544977 286394
rect 539564 283448 541638 284040
rect 539784 282923 541422 283415
rect 536849 282298 544359 282890
rect 537314 281290 543888 282108
rect 11705 276597 14643 279793
rect 17369 271931 18789 273371
rect 18889 271931 20309 273371
rect 20410 270940 21830 274370
rect 21930 270680 23350 274626
rect 27080 272310 28000 272960
rect 28080 271950 28750 273316
rect 28830 271695 30250 273577
rect 30390 269150 45200 276180
rect 537314 275978 543894 281290
rect 568100 280100 578520 281414
rect 11705 265527 14643 268723
rect 537314 268522 543884 275978
rect 537312 267278 543884 268522
rect 5780 251200 16200 252514
rect 5780 240800 16200 242114
<< nmos >>
rect 5990 304278 15990 304318
rect 5990 304180 15990 304220
rect 5990 304082 15990 304122
rect 5990 303984 15990 304024
rect 5990 303886 15990 303926
rect 5990 303788 15990 303828
rect 5990 303690 15990 303730
rect 5990 303592 15990 303632
rect 5990 303494 15990 303534
rect 5990 303396 15990 303436
rect 559996 295810 560036 305810
rect 560094 295810 560134 305810
rect 560192 295810 560232 305810
rect 560290 295810 560330 305810
rect 560388 295810 560428 305810
rect 560486 295810 560526 305810
rect 560584 295810 560624 305810
rect 560682 295810 560722 305810
rect 560780 295810 560820 305810
rect 560878 295810 560918 305810
rect 569196 295810 569236 305810
rect 569294 295810 569334 305810
rect 569392 295810 569432 305810
rect 569490 295810 569530 305810
rect 569588 295810 569628 305810
rect 569686 295810 569726 305810
rect 569784 295810 569824 305810
rect 569882 295810 569922 305810
rect 569980 295810 570020 305810
rect 570078 295810 570118 305810
rect 5990 293878 15990 293918
rect 5990 293780 15990 293820
rect 5990 293682 15990 293722
rect 5990 293584 15990 293624
rect 5990 293486 15990 293526
rect 5990 293388 15990 293428
rect 5990 293290 15990 293330
rect 5990 293192 15990 293232
rect 5990 293094 15990 293134
rect 5990 292996 15990 293036
rect 536459 288918 537459 289018
rect 537677 288918 538677 289018
rect 538895 288918 539895 289018
rect 540113 288918 541113 289018
rect 541331 288918 542331 289018
rect 542549 288918 543549 289018
rect 543767 288918 544767 289018
rect 536459 288418 537459 288518
rect 537677 288418 538677 288518
rect 538895 288418 539895 288518
rect 540113 288418 541113 288518
rect 541331 288418 542331 288518
rect 542549 288418 543549 288518
rect 543767 288418 544767 288518
rect 537019 287818 538019 288018
rect 538237 287818 539237 288018
rect 539455 287818 540455 288018
rect 540673 287818 541673 288018
rect 541891 287818 542891 288018
rect 543109 287818 544109 288018
rect 568290 288658 578290 288698
rect 568290 288560 578290 288600
rect 568290 288462 578290 288502
rect 568290 288364 578290 288404
rect 568290 288266 578290 288306
rect 568290 288168 578290 288208
rect 568290 288070 578290 288110
rect 568290 287972 578290 288012
rect 568290 287874 578290 287914
rect 568290 287776 578290 287816
rect 537019 287198 538019 287398
rect 538237 287198 539237 287398
rect 539455 287198 540455 287398
rect 540673 287198 541673 287398
rect 541891 287198 542891 287398
rect 543109 287198 544109 287398
rect 536459 286598 537459 286798
rect 537677 286598 538677 286798
rect 538895 286598 539895 286798
rect 540113 286598 541113 286798
rect 541331 286598 542331 286798
rect 542549 286598 543549 286798
rect 543767 286598 544767 286798
rect 536459 285998 537459 286198
rect 537677 285998 538677 286198
rect 538895 285998 539895 286198
rect 540113 285998 541113 286198
rect 541331 285998 542331 286198
rect 542549 285998 543549 286198
rect 543767 285998 544767 286198
rect 539774 283644 540024 283844
rect 540242 283644 540492 283844
rect 540710 283644 540960 283844
rect 541178 283644 541428 283844
rect 539994 283119 540494 283219
rect 540712 283119 541212 283219
rect 537059 282494 538059 282694
rect 538277 282494 539277 282694
rect 539495 282494 540495 282694
rect 540713 282494 541713 282694
rect 541931 282494 542931 282694
rect 543149 282494 544149 282694
rect 568310 281178 578310 281218
rect 568310 281080 578310 281120
rect 568310 280982 578310 281022
rect 568310 280884 578310 280924
rect 568310 280786 578310 280826
rect 568310 280688 578310 280728
rect 568310 280590 578310 280630
rect 568310 280492 578310 280532
rect 568310 280394 578310 280434
rect 568310 280296 578310 280336
rect 17579 273075 18579 273175
rect 17579 272917 18579 273017
rect 17579 272759 18579 272859
rect 17579 272601 18579 272701
rect 17579 272443 18579 272543
rect 17579 272285 18579 272385
rect 17579 272127 18579 272227
rect 19099 273075 20099 273175
rect 19099 272917 20099 273017
rect 19099 272759 20099 272859
rect 19099 272601 20099 272701
rect 19099 272443 20099 272543
rect 19099 272285 20099 272385
rect 19099 272127 20099 272227
rect 20620 273974 21620 274174
rect 20620 273716 21620 273916
rect 20620 273458 21620 273658
rect 20620 273200 21620 273400
rect 20620 272942 21620 273142
rect 20620 272684 21620 272884
rect 20620 272426 21620 272626
rect 20620 272168 21620 272368
rect 20620 271910 21620 272110
rect 20620 271652 21620 271852
rect 20620 271394 21620 271594
rect 20620 271136 21620 271336
rect 22140 274230 23140 274430
rect 22140 273972 23140 274172
rect 22140 273714 23140 273914
rect 22140 273456 23140 273656
rect 22140 273198 23140 273398
rect 22140 272940 23140 273140
rect 22140 272682 23140 272882
rect 22140 272424 23140 272624
rect 22140 272166 23140 272366
rect 22140 271908 23140 272108
rect 22140 271650 23140 271850
rect 22140 271392 23140 271592
rect 22140 271134 23140 271334
rect 22140 270876 23140 271076
rect 27290 272664 27790 272764
rect 27290 272506 27790 272606
rect 28290 272920 28540 273120
rect 28290 272662 28540 272862
rect 28290 272404 28540 272604
rect 28290 272146 28540 272346
rect 29040 273181 30040 273381
rect 29040 272923 30040 273123
rect 29040 272665 30040 272865
rect 29040 272407 30040 272607
rect 29040 272149 30040 272349
rect 29040 271891 30040 272091
rect 5990 252278 15990 252318
rect 5990 252180 15990 252220
rect 5990 252082 15990 252122
rect 5990 251984 15990 252024
rect 5990 251886 15990 251926
rect 5990 251788 15990 251828
rect 5990 251690 15990 251730
rect 5990 251592 15990 251632
rect 5990 251494 15990 251534
rect 5990 251396 15990 251436
rect 5990 241878 15990 241918
rect 5990 241780 15990 241820
rect 5990 241682 15990 241722
rect 5990 241584 15990 241624
rect 5990 241486 15990 241526
rect 5990 241388 15990 241428
rect 5990 241290 15990 241330
rect 5990 241192 15990 241232
rect 5990 241094 15990 241134
rect 5990 240996 15990 241036
<< pmos >>
rect 536368 294638 537368 294738
rect 537604 294638 538604 294738
rect 538840 294638 539840 294738
rect 540076 294638 541076 294738
rect 541312 294638 542312 294738
rect 542548 294638 543548 294738
rect 543784 294638 544784 294738
rect 536368 294098 537368 294198
rect 537604 294098 538604 294198
rect 538840 294098 539840 294198
rect 540076 294098 541076 294198
rect 541312 294098 542312 294198
rect 542548 294098 543548 294198
rect 543784 294098 544784 294198
rect 536368 293558 537368 293658
rect 537604 293558 538604 293658
rect 538840 293558 539840 293658
rect 540076 293558 541076 293658
rect 541312 293558 542312 293658
rect 542548 293558 543548 293658
rect 543784 293558 544784 293658
rect 536368 293018 537368 293118
rect 537604 293018 538604 293118
rect 538840 293018 539840 293118
rect 540076 293018 541076 293118
rect 541312 293018 542312 293118
rect 542548 293018 543548 293118
rect 543784 293018 544784 293118
rect 536368 292438 537368 292538
rect 537604 292438 538604 292538
rect 538840 292438 539840 292538
rect 540076 292438 541076 292538
rect 541312 292438 542312 292538
rect 542548 292438 543548 292538
rect 543784 292438 544784 292538
rect 536368 291858 537368 291958
rect 537604 291858 538604 291958
rect 538840 291858 539840 291958
rect 540076 291858 541076 291958
rect 541312 291858 542312 291958
rect 542548 291858 543548 291958
rect 543784 291858 544784 291958
rect 534528 291318 535528 291418
rect 535764 291318 536764 291418
rect 537000 291318 538000 291418
rect 538236 291318 539236 291418
rect 539472 291318 540472 291418
rect 540708 291318 541708 291418
rect 541944 291318 542944 291418
rect 543180 291318 544180 291418
rect 544416 291318 545416 291418
rect 545652 291318 546652 291418
rect 534528 290778 535528 290878
rect 535764 290778 536764 290878
rect 537000 290778 538000 290878
rect 538236 290778 539236 290878
rect 539472 290778 540472 290878
rect 540708 290778 541708 290878
rect 541944 290778 542944 290878
rect 543180 290778 544180 290878
rect 544416 290778 545416 290878
rect 545652 290778 546652 290878
rect 534528 290238 535528 290338
rect 535764 290238 536764 290338
rect 537000 290238 538000 290338
rect 538236 290238 539236 290338
rect 539472 290238 540472 290338
rect 540708 290238 541708 290338
rect 541944 290238 542944 290338
rect 543180 290238 544180 290338
rect 544416 290238 545416 290338
rect 545652 290238 546652 290338
rect 534528 289698 535528 289798
rect 535764 289698 536764 289798
rect 537000 289698 538000 289798
rect 538236 289698 539236 289798
rect 539472 289698 540472 289798
rect 540708 289698 541708 289798
rect 541944 289698 542944 289798
rect 543180 289698 544180 289798
rect 544416 289698 545416 289798
rect 545652 289698 546652 289798
rect 537013 285024 538013 285224
rect 538249 285024 539249 285224
rect 539485 285024 540485 285224
rect 540721 285024 541721 285224
rect 541957 285024 542957 285224
rect 543193 285024 544193 285224
rect 537013 284434 538013 284634
rect 538249 284434 539249 284634
rect 539485 284434 540485 284634
rect 540721 284434 541721 284634
rect 541957 284434 542957 284634
rect 543193 284434 544193 284634
rect 12801 275688 13801 275788
rect 12801 275530 13801 275630
rect 12801 275372 13801 275472
rect 12801 275214 13801 275314
rect 12801 275056 13801 275156
rect 12801 274898 13801 274998
rect 12801 274740 13801 274840
rect 12801 274582 13801 274682
rect 12801 274424 13801 274524
rect 12801 274266 13801 274366
rect 12801 274108 13801 274208
rect 12801 273950 13801 274050
rect 12801 273792 13801 273892
rect 12801 273634 13801 273734
rect 12801 273476 13801 273576
rect 12801 273318 13801 273418
rect 12801 273160 13801 273260
rect 12801 273002 13801 273102
rect 12801 272844 13801 272944
rect 12801 272686 13801 272786
rect 12801 272528 13801 272628
rect 12801 272370 13801 272470
rect 12801 272212 13801 272312
rect 12801 272054 13801 272154
rect 12801 271896 13801 271996
rect 12801 271738 13801 271838
rect 12801 271580 13801 271680
rect 12801 271422 13801 271522
rect 12801 271264 13801 271364
rect 12801 271106 13801 271206
rect 12801 270948 13801 271048
rect 12801 270790 13801 270890
rect 12801 270632 13801 270732
rect 12801 270474 13801 270574
rect 12801 270316 13801 270416
rect 12801 270158 13801 270258
rect 12801 270000 13801 270100
rect 12801 269842 13801 269942
rect 12801 269684 13801 269784
rect 12801 269526 13801 269626
rect 14471 274186 15471 274286
rect 14471 274028 15471 274128
rect 14471 273870 15471 273970
rect 14471 273712 15471 273812
rect 14471 273554 15471 273654
rect 14471 273396 15471 273496
rect 14471 273238 15471 273338
rect 14471 273080 15471 273180
rect 14471 272922 15471 273022
rect 14471 272764 15471 272864
rect 14471 272606 15471 272706
rect 14471 272448 15471 272548
rect 14471 272290 15471 272390
rect 14471 272132 15471 272232
rect 14471 271974 15471 272074
rect 14471 271816 15471 271916
rect 14471 271658 15471 271758
rect 14471 271500 15471 271600
rect 14471 271342 15471 271442
rect 14471 271184 15471 271284
rect 14471 271026 15471 271126
rect 16011 274186 17011 274286
rect 16011 274028 17011 274128
rect 16011 273870 17011 273970
rect 16011 273712 17011 273812
rect 16011 273554 17011 273654
rect 16011 273396 17011 273496
rect 16011 273238 17011 273338
rect 16011 273080 17011 273180
rect 16011 272922 17011 273022
rect 16011 272764 17011 272864
rect 16011 272606 17011 272706
rect 16011 272448 17011 272548
rect 16011 272290 17011 272390
rect 16011 272132 17011 272232
rect 16011 271974 17011 272074
rect 16011 271816 17011 271916
rect 16011 271658 17011 271758
rect 16011 271500 17011 271600
rect 16011 271342 17011 271442
rect 16011 271184 17011 271284
rect 16011 271026 17011 271126
rect 24181 273196 25181 273396
rect 24181 272938 25181 273138
rect 24181 272680 25181 272880
rect 24181 272422 25181 272622
rect 24181 272164 25181 272364
rect 24181 271906 25181 272106
rect 25681 273196 26681 273396
rect 25681 272938 26681 273138
rect 25681 272680 26681 272880
rect 25681 272422 26681 272622
rect 25681 272164 26681 272364
rect 25681 271906 26681 272106
<< ndiff >>
rect 5990 304364 15990 304376
rect 5990 304330 6002 304364
rect 15978 304330 15990 304364
rect 5990 304318 15990 304330
rect 5990 304266 15990 304278
rect 5990 304232 6002 304266
rect 15978 304232 15990 304266
rect 5990 304220 15990 304232
rect 5990 304168 15990 304180
rect 5990 304134 6002 304168
rect 15978 304134 15990 304168
rect 5990 304122 15990 304134
rect 5990 304070 15990 304082
rect 5990 304036 6002 304070
rect 15978 304036 15990 304070
rect 5990 304024 15990 304036
rect 5990 303972 15990 303984
rect 5990 303938 6002 303972
rect 15978 303938 15990 303972
rect 5990 303926 15990 303938
rect 5990 303874 15990 303886
rect 5990 303840 6002 303874
rect 15978 303840 15990 303874
rect 5990 303828 15990 303840
rect 5990 303776 15990 303788
rect 5990 303742 6002 303776
rect 15978 303742 15990 303776
rect 5990 303730 15990 303742
rect 5990 303678 15990 303690
rect 5990 303644 6002 303678
rect 15978 303644 15990 303678
rect 5990 303632 15990 303644
rect 5990 303580 15990 303592
rect 5990 303546 6002 303580
rect 15978 303546 15990 303580
rect 5990 303534 15990 303546
rect 5990 303482 15990 303494
rect 5990 303448 6002 303482
rect 15978 303448 15990 303482
rect 5990 303436 15990 303448
rect 5990 303384 15990 303396
rect 5990 303350 6002 303384
rect 15978 303350 15990 303384
rect 5990 303338 15990 303350
rect 559938 305798 559996 305810
rect 559938 295822 559950 305798
rect 559984 295822 559996 305798
rect 559938 295810 559996 295822
rect 560036 305798 560094 305810
rect 560036 295822 560048 305798
rect 560082 295822 560094 305798
rect 560036 295810 560094 295822
rect 560134 305798 560192 305810
rect 560134 295822 560146 305798
rect 560180 295822 560192 305798
rect 560134 295810 560192 295822
rect 560232 305798 560290 305810
rect 560232 295822 560244 305798
rect 560278 295822 560290 305798
rect 560232 295810 560290 295822
rect 560330 305798 560388 305810
rect 560330 295822 560342 305798
rect 560376 295822 560388 305798
rect 560330 295810 560388 295822
rect 560428 305798 560486 305810
rect 560428 295822 560440 305798
rect 560474 295822 560486 305798
rect 560428 295810 560486 295822
rect 560526 305798 560584 305810
rect 560526 295822 560538 305798
rect 560572 295822 560584 305798
rect 560526 295810 560584 295822
rect 560624 305798 560682 305810
rect 560624 295822 560636 305798
rect 560670 295822 560682 305798
rect 560624 295810 560682 295822
rect 560722 305798 560780 305810
rect 560722 295822 560734 305798
rect 560768 295822 560780 305798
rect 560722 295810 560780 295822
rect 560820 305798 560878 305810
rect 560820 295822 560832 305798
rect 560866 295822 560878 305798
rect 560820 295810 560878 295822
rect 560918 305798 560976 305810
rect 560918 295822 560930 305798
rect 560964 295822 560976 305798
rect 560918 295810 560976 295822
rect 569138 305798 569196 305810
rect 569138 295822 569150 305798
rect 569184 295822 569196 305798
rect 569138 295810 569196 295822
rect 569236 305798 569294 305810
rect 569236 295822 569248 305798
rect 569282 295822 569294 305798
rect 569236 295810 569294 295822
rect 569334 305798 569392 305810
rect 569334 295822 569346 305798
rect 569380 295822 569392 305798
rect 569334 295810 569392 295822
rect 569432 305798 569490 305810
rect 569432 295822 569444 305798
rect 569478 295822 569490 305798
rect 569432 295810 569490 295822
rect 569530 305798 569588 305810
rect 569530 295822 569542 305798
rect 569576 295822 569588 305798
rect 569530 295810 569588 295822
rect 569628 305798 569686 305810
rect 569628 295822 569640 305798
rect 569674 295822 569686 305798
rect 569628 295810 569686 295822
rect 569726 305798 569784 305810
rect 569726 295822 569738 305798
rect 569772 295822 569784 305798
rect 569726 295810 569784 295822
rect 569824 305798 569882 305810
rect 569824 295822 569836 305798
rect 569870 295822 569882 305798
rect 569824 295810 569882 295822
rect 569922 305798 569980 305810
rect 569922 295822 569934 305798
rect 569968 295822 569980 305798
rect 569922 295810 569980 295822
rect 570020 305798 570078 305810
rect 570020 295822 570032 305798
rect 570066 295822 570078 305798
rect 570020 295810 570078 295822
rect 570118 305798 570176 305810
rect 570118 295822 570130 305798
rect 570164 295822 570176 305798
rect 570118 295810 570176 295822
rect 5990 293964 15990 293976
rect 5990 293930 6002 293964
rect 15978 293930 15990 293964
rect 5990 293918 15990 293930
rect 5990 293866 15990 293878
rect 5990 293832 6002 293866
rect 15978 293832 15990 293866
rect 5990 293820 15990 293832
rect 5990 293768 15990 293780
rect 5990 293734 6002 293768
rect 15978 293734 15990 293768
rect 5990 293722 15990 293734
rect 5990 293670 15990 293682
rect 5990 293636 6002 293670
rect 15978 293636 15990 293670
rect 5990 293624 15990 293636
rect 5990 293572 15990 293584
rect 5990 293538 6002 293572
rect 15978 293538 15990 293572
rect 5990 293526 15990 293538
rect 5990 293474 15990 293486
rect 5990 293440 6002 293474
rect 15978 293440 15990 293474
rect 5990 293428 15990 293440
rect 5990 293376 15990 293388
rect 5990 293342 6002 293376
rect 15978 293342 15990 293376
rect 5990 293330 15990 293342
rect 5990 293278 15990 293290
rect 5990 293244 6002 293278
rect 15978 293244 15990 293278
rect 5990 293232 15990 293244
rect 5990 293180 15990 293192
rect 5990 293146 6002 293180
rect 15978 293146 15990 293180
rect 5990 293134 15990 293146
rect 5990 293082 15990 293094
rect 5990 293048 6002 293082
rect 15978 293048 15990 293082
rect 5990 293036 15990 293048
rect 5990 292984 15990 292996
rect 5990 292950 6002 292984
rect 15978 292950 15990 292984
rect 5990 292938 15990 292950
rect 536459 289064 537459 289076
rect 536459 289030 536471 289064
rect 537447 289030 537459 289064
rect 536459 289018 537459 289030
rect 537677 289064 538677 289076
rect 537677 289030 537689 289064
rect 538665 289030 538677 289064
rect 537677 289018 538677 289030
rect 538895 289064 539895 289076
rect 538895 289030 538907 289064
rect 539883 289030 539895 289064
rect 538895 289018 539895 289030
rect 540113 289064 541113 289076
rect 540113 289030 540125 289064
rect 541101 289030 541113 289064
rect 540113 289018 541113 289030
rect 541331 289064 542331 289076
rect 541331 289030 541343 289064
rect 542319 289030 542331 289064
rect 541331 289018 542331 289030
rect 542549 289064 543549 289076
rect 542549 289030 542561 289064
rect 543537 289030 543549 289064
rect 542549 289018 543549 289030
rect 543767 289064 544767 289076
rect 543767 289030 543779 289064
rect 544755 289030 544767 289064
rect 543767 289018 544767 289030
rect 536459 288906 537459 288918
rect 536459 288872 536471 288906
rect 537447 288872 537459 288906
rect 536459 288860 537459 288872
rect 537677 288906 538677 288918
rect 537677 288872 537689 288906
rect 538665 288872 538677 288906
rect 537677 288860 538677 288872
rect 538895 288906 539895 288918
rect 538895 288872 538907 288906
rect 539883 288872 539895 288906
rect 538895 288860 539895 288872
rect 540113 288906 541113 288918
rect 540113 288872 540125 288906
rect 541101 288872 541113 288906
rect 540113 288860 541113 288872
rect 541331 288906 542331 288918
rect 541331 288872 541343 288906
rect 542319 288872 542331 288906
rect 541331 288860 542331 288872
rect 542549 288906 543549 288918
rect 542549 288872 542561 288906
rect 543537 288872 543549 288906
rect 542549 288860 543549 288872
rect 543767 288906 544767 288918
rect 543767 288872 543779 288906
rect 544755 288872 544767 288906
rect 543767 288860 544767 288872
rect 536459 288564 537459 288576
rect 536459 288530 536471 288564
rect 537447 288530 537459 288564
rect 536459 288518 537459 288530
rect 537677 288564 538677 288576
rect 537677 288530 537689 288564
rect 538665 288530 538677 288564
rect 537677 288518 538677 288530
rect 538895 288564 539895 288576
rect 538895 288530 538907 288564
rect 539883 288530 539895 288564
rect 538895 288518 539895 288530
rect 540113 288564 541113 288576
rect 540113 288530 540125 288564
rect 541101 288530 541113 288564
rect 540113 288518 541113 288530
rect 541331 288564 542331 288576
rect 541331 288530 541343 288564
rect 542319 288530 542331 288564
rect 541331 288518 542331 288530
rect 542549 288564 543549 288576
rect 542549 288530 542561 288564
rect 543537 288530 543549 288564
rect 542549 288518 543549 288530
rect 543767 288564 544767 288576
rect 543767 288530 543779 288564
rect 544755 288530 544767 288564
rect 543767 288518 544767 288530
rect 536459 288406 537459 288418
rect 536459 288372 536471 288406
rect 537447 288372 537459 288406
rect 536459 288360 537459 288372
rect 537677 288406 538677 288418
rect 537677 288372 537689 288406
rect 538665 288372 538677 288406
rect 537677 288360 538677 288372
rect 538895 288406 539895 288418
rect 538895 288372 538907 288406
rect 539883 288372 539895 288406
rect 538895 288360 539895 288372
rect 540113 288406 541113 288418
rect 540113 288372 540125 288406
rect 541101 288372 541113 288406
rect 540113 288360 541113 288372
rect 541331 288406 542331 288418
rect 541331 288372 541343 288406
rect 542319 288372 542331 288406
rect 541331 288360 542331 288372
rect 542549 288406 543549 288418
rect 542549 288372 542561 288406
rect 543537 288372 543549 288406
rect 542549 288360 543549 288372
rect 543767 288406 544767 288418
rect 543767 288372 543779 288406
rect 544755 288372 544767 288406
rect 543767 288360 544767 288372
rect 537019 288064 538019 288076
rect 537019 288030 537031 288064
rect 538007 288030 538019 288064
rect 537019 288018 538019 288030
rect 538237 288064 539237 288076
rect 538237 288030 538249 288064
rect 539225 288030 539237 288064
rect 538237 288018 539237 288030
rect 539455 288064 540455 288076
rect 539455 288030 539467 288064
rect 540443 288030 540455 288064
rect 539455 288018 540455 288030
rect 540673 288064 541673 288076
rect 540673 288030 540685 288064
rect 541661 288030 541673 288064
rect 540673 288018 541673 288030
rect 541891 288064 542891 288076
rect 541891 288030 541903 288064
rect 542879 288030 542891 288064
rect 541891 288018 542891 288030
rect 543109 288064 544109 288076
rect 543109 288030 543121 288064
rect 544097 288030 544109 288064
rect 543109 288018 544109 288030
rect 537019 287806 538019 287818
rect 537019 287772 537031 287806
rect 538007 287772 538019 287806
rect 537019 287760 538019 287772
rect 538237 287806 539237 287818
rect 538237 287772 538249 287806
rect 539225 287772 539237 287806
rect 538237 287760 539237 287772
rect 539455 287806 540455 287818
rect 539455 287772 539467 287806
rect 540443 287772 540455 287806
rect 539455 287760 540455 287772
rect 540673 287806 541673 287818
rect 540673 287772 540685 287806
rect 541661 287772 541673 287806
rect 540673 287760 541673 287772
rect 541891 287806 542891 287818
rect 541891 287772 541903 287806
rect 542879 287772 542891 287806
rect 541891 287760 542891 287772
rect 543109 287806 544109 287818
rect 543109 287772 543121 287806
rect 544097 287772 544109 287806
rect 543109 287760 544109 287772
rect 568290 288744 578290 288756
rect 568290 288710 568302 288744
rect 578278 288710 578290 288744
rect 568290 288698 578290 288710
rect 568290 288646 578290 288658
rect 568290 288612 568302 288646
rect 578278 288612 578290 288646
rect 568290 288600 578290 288612
rect 568290 288548 578290 288560
rect 568290 288514 568302 288548
rect 578278 288514 578290 288548
rect 568290 288502 578290 288514
rect 568290 288450 578290 288462
rect 568290 288416 568302 288450
rect 578278 288416 578290 288450
rect 568290 288404 578290 288416
rect 568290 288352 578290 288364
rect 568290 288318 568302 288352
rect 578278 288318 578290 288352
rect 568290 288306 578290 288318
rect 568290 288254 578290 288266
rect 568290 288220 568302 288254
rect 578278 288220 578290 288254
rect 568290 288208 578290 288220
rect 568290 288156 578290 288168
rect 568290 288122 568302 288156
rect 578278 288122 578290 288156
rect 568290 288110 578290 288122
rect 568290 288058 578290 288070
rect 568290 288024 568302 288058
rect 578278 288024 578290 288058
rect 568290 288012 578290 288024
rect 568290 287960 578290 287972
rect 568290 287926 568302 287960
rect 578278 287926 578290 287960
rect 568290 287914 578290 287926
rect 568290 287862 578290 287874
rect 568290 287828 568302 287862
rect 578278 287828 578290 287862
rect 568290 287816 578290 287828
rect 568290 287764 578290 287776
rect 568290 287730 568302 287764
rect 578278 287730 578290 287764
rect 568290 287718 578290 287730
rect 537019 287444 538019 287456
rect 537019 287410 537031 287444
rect 538007 287410 538019 287444
rect 537019 287398 538019 287410
rect 538237 287444 539237 287456
rect 538237 287410 538249 287444
rect 539225 287410 539237 287444
rect 538237 287398 539237 287410
rect 539455 287444 540455 287456
rect 539455 287410 539467 287444
rect 540443 287410 540455 287444
rect 539455 287398 540455 287410
rect 540673 287444 541673 287456
rect 540673 287410 540685 287444
rect 541661 287410 541673 287444
rect 540673 287398 541673 287410
rect 541891 287444 542891 287456
rect 541891 287410 541903 287444
rect 542879 287410 542891 287444
rect 541891 287398 542891 287410
rect 543109 287444 544109 287456
rect 543109 287410 543121 287444
rect 544097 287410 544109 287444
rect 543109 287398 544109 287410
rect 537019 287186 538019 287198
rect 537019 287152 537031 287186
rect 538007 287152 538019 287186
rect 537019 287140 538019 287152
rect 538237 287186 539237 287198
rect 538237 287152 538249 287186
rect 539225 287152 539237 287186
rect 538237 287140 539237 287152
rect 539455 287186 540455 287198
rect 539455 287152 539467 287186
rect 540443 287152 540455 287186
rect 539455 287140 540455 287152
rect 540673 287186 541673 287198
rect 540673 287152 540685 287186
rect 541661 287152 541673 287186
rect 540673 287140 541673 287152
rect 541891 287186 542891 287198
rect 541891 287152 541903 287186
rect 542879 287152 542891 287186
rect 541891 287140 542891 287152
rect 543109 287186 544109 287198
rect 543109 287152 543121 287186
rect 544097 287152 544109 287186
rect 543109 287140 544109 287152
rect 536459 286844 537459 286856
rect 536459 286810 536471 286844
rect 537447 286810 537459 286844
rect 536459 286798 537459 286810
rect 537677 286844 538677 286856
rect 537677 286810 537689 286844
rect 538665 286810 538677 286844
rect 537677 286798 538677 286810
rect 538895 286844 539895 286856
rect 538895 286810 538907 286844
rect 539883 286810 539895 286844
rect 538895 286798 539895 286810
rect 540113 286844 541113 286856
rect 540113 286810 540125 286844
rect 541101 286810 541113 286844
rect 540113 286798 541113 286810
rect 541331 286844 542331 286856
rect 541331 286810 541343 286844
rect 542319 286810 542331 286844
rect 541331 286798 542331 286810
rect 542549 286844 543549 286856
rect 542549 286810 542561 286844
rect 543537 286810 543549 286844
rect 542549 286798 543549 286810
rect 543767 286844 544767 286856
rect 543767 286810 543779 286844
rect 544755 286810 544767 286844
rect 543767 286798 544767 286810
rect 536459 286586 537459 286598
rect 536459 286552 536471 286586
rect 537447 286552 537459 286586
rect 536459 286540 537459 286552
rect 537677 286586 538677 286598
rect 537677 286552 537689 286586
rect 538665 286552 538677 286586
rect 537677 286540 538677 286552
rect 538895 286586 539895 286598
rect 538895 286552 538907 286586
rect 539883 286552 539895 286586
rect 538895 286540 539895 286552
rect 540113 286586 541113 286598
rect 540113 286552 540125 286586
rect 541101 286552 541113 286586
rect 540113 286540 541113 286552
rect 541331 286586 542331 286598
rect 541331 286552 541343 286586
rect 542319 286552 542331 286586
rect 541331 286540 542331 286552
rect 542549 286586 543549 286598
rect 542549 286552 542561 286586
rect 543537 286552 543549 286586
rect 542549 286540 543549 286552
rect 543767 286586 544767 286598
rect 543767 286552 543779 286586
rect 544755 286552 544767 286586
rect 543767 286540 544767 286552
rect 536459 286244 537459 286256
rect 536459 286210 536471 286244
rect 537447 286210 537459 286244
rect 536459 286198 537459 286210
rect 537677 286244 538677 286256
rect 537677 286210 537689 286244
rect 538665 286210 538677 286244
rect 537677 286198 538677 286210
rect 538895 286244 539895 286256
rect 538895 286210 538907 286244
rect 539883 286210 539895 286244
rect 538895 286198 539895 286210
rect 540113 286244 541113 286256
rect 540113 286210 540125 286244
rect 541101 286210 541113 286244
rect 540113 286198 541113 286210
rect 541331 286244 542331 286256
rect 541331 286210 541343 286244
rect 542319 286210 542331 286244
rect 541331 286198 542331 286210
rect 542549 286244 543549 286256
rect 542549 286210 542561 286244
rect 543537 286210 543549 286244
rect 542549 286198 543549 286210
rect 543767 286244 544767 286256
rect 543767 286210 543779 286244
rect 544755 286210 544767 286244
rect 543767 286198 544767 286210
rect 536459 285986 537459 285998
rect 536459 285952 536471 285986
rect 537447 285952 537459 285986
rect 536459 285940 537459 285952
rect 537677 285986 538677 285998
rect 537677 285952 537689 285986
rect 538665 285952 538677 285986
rect 537677 285940 538677 285952
rect 538895 285986 539895 285998
rect 538895 285952 538907 285986
rect 539883 285952 539895 285986
rect 538895 285940 539895 285952
rect 540113 285986 541113 285998
rect 540113 285952 540125 285986
rect 541101 285952 541113 285986
rect 540113 285940 541113 285952
rect 541331 285986 542331 285998
rect 541331 285952 541343 285986
rect 542319 285952 542331 285986
rect 541331 285940 542331 285952
rect 542549 285986 543549 285998
rect 542549 285952 542561 285986
rect 543537 285952 543549 285986
rect 542549 285940 543549 285952
rect 543767 285986 544767 285998
rect 543767 285952 543779 285986
rect 544755 285952 544767 285986
rect 543767 285940 544767 285952
rect 539774 283890 540024 283902
rect 539774 283856 539786 283890
rect 540012 283856 540024 283890
rect 539774 283844 540024 283856
rect 540242 283890 540492 283902
rect 540242 283856 540254 283890
rect 540480 283856 540492 283890
rect 540242 283844 540492 283856
rect 540710 283890 540960 283902
rect 540710 283856 540722 283890
rect 540948 283856 540960 283890
rect 540710 283844 540960 283856
rect 541178 283890 541428 283902
rect 541178 283856 541190 283890
rect 541416 283856 541428 283890
rect 541178 283844 541428 283856
rect 539774 283632 540024 283644
rect 539774 283598 539786 283632
rect 540012 283598 540024 283632
rect 539774 283586 540024 283598
rect 540242 283632 540492 283644
rect 540242 283598 540254 283632
rect 540480 283598 540492 283632
rect 540242 283586 540492 283598
rect 540710 283632 540960 283644
rect 540710 283598 540722 283632
rect 540948 283598 540960 283632
rect 540710 283586 540960 283598
rect 541178 283632 541428 283644
rect 541178 283598 541190 283632
rect 541416 283598 541428 283632
rect 541178 283586 541428 283598
rect 539994 283265 540494 283277
rect 539994 283231 540006 283265
rect 540482 283231 540494 283265
rect 539994 283219 540494 283231
rect 540712 283265 541212 283277
rect 540712 283231 540724 283265
rect 541200 283231 541212 283265
rect 540712 283219 541212 283231
rect 539994 283107 540494 283119
rect 539994 283073 540006 283107
rect 540482 283073 540494 283107
rect 539994 283061 540494 283073
rect 540712 283107 541212 283119
rect 540712 283073 540724 283107
rect 541200 283073 541212 283107
rect 540712 283061 541212 283073
rect 537059 282740 538059 282752
rect 537059 282706 537071 282740
rect 538047 282706 538059 282740
rect 537059 282694 538059 282706
rect 538277 282740 539277 282752
rect 538277 282706 538289 282740
rect 539265 282706 539277 282740
rect 538277 282694 539277 282706
rect 539495 282740 540495 282752
rect 539495 282706 539507 282740
rect 540483 282706 540495 282740
rect 539495 282694 540495 282706
rect 540713 282740 541713 282752
rect 540713 282706 540725 282740
rect 541701 282706 541713 282740
rect 540713 282694 541713 282706
rect 541931 282740 542931 282752
rect 541931 282706 541943 282740
rect 542919 282706 542931 282740
rect 541931 282694 542931 282706
rect 543149 282740 544149 282752
rect 543149 282706 543161 282740
rect 544137 282706 544149 282740
rect 543149 282694 544149 282706
rect 537059 282482 538059 282494
rect 537059 282448 537071 282482
rect 538047 282448 538059 282482
rect 537059 282436 538059 282448
rect 538277 282482 539277 282494
rect 538277 282448 538289 282482
rect 539265 282448 539277 282482
rect 538277 282436 539277 282448
rect 539495 282482 540495 282494
rect 539495 282448 539507 282482
rect 540483 282448 540495 282482
rect 539495 282436 540495 282448
rect 540713 282482 541713 282494
rect 540713 282448 540725 282482
rect 541701 282448 541713 282482
rect 540713 282436 541713 282448
rect 541931 282482 542931 282494
rect 541931 282448 541943 282482
rect 542919 282448 542931 282482
rect 541931 282436 542931 282448
rect 543149 282482 544149 282494
rect 543149 282448 543161 282482
rect 544137 282448 544149 282482
rect 543149 282436 544149 282448
rect 568310 281264 578310 281276
rect 568310 281230 568322 281264
rect 578298 281230 578310 281264
rect 568310 281218 578310 281230
rect 568310 281166 578310 281178
rect 568310 281132 568322 281166
rect 578298 281132 578310 281166
rect 568310 281120 578310 281132
rect 568310 281068 578310 281080
rect 568310 281034 568322 281068
rect 578298 281034 578310 281068
rect 568310 281022 578310 281034
rect 568310 280970 578310 280982
rect 568310 280936 568322 280970
rect 578298 280936 578310 280970
rect 568310 280924 578310 280936
rect 568310 280872 578310 280884
rect 568310 280838 568322 280872
rect 578298 280838 578310 280872
rect 568310 280826 578310 280838
rect 568310 280774 578310 280786
rect 568310 280740 568322 280774
rect 578298 280740 578310 280774
rect 568310 280728 578310 280740
rect 568310 280676 578310 280688
rect 568310 280642 568322 280676
rect 578298 280642 578310 280676
rect 568310 280630 578310 280642
rect 568310 280578 578310 280590
rect 568310 280544 568322 280578
rect 578298 280544 578310 280578
rect 568310 280532 578310 280544
rect 568310 280480 578310 280492
rect 568310 280446 568322 280480
rect 578298 280446 578310 280480
rect 568310 280434 578310 280446
rect 568310 280382 578310 280394
rect 568310 280348 568322 280382
rect 578298 280348 578310 280382
rect 568310 280336 578310 280348
rect 568310 280284 578310 280296
rect 568310 280250 568322 280284
rect 578298 280250 578310 280284
rect 568310 280238 578310 280250
rect 17579 273221 18579 273233
rect 17579 273187 17591 273221
rect 18567 273187 18579 273221
rect 17579 273175 18579 273187
rect 17579 273063 18579 273075
rect 17579 273029 17591 273063
rect 18567 273029 18579 273063
rect 17579 273017 18579 273029
rect 17579 272905 18579 272917
rect 17579 272871 17591 272905
rect 18567 272871 18579 272905
rect 17579 272859 18579 272871
rect 17579 272747 18579 272759
rect 17579 272713 17591 272747
rect 18567 272713 18579 272747
rect 17579 272701 18579 272713
rect 17579 272589 18579 272601
rect 17579 272555 17591 272589
rect 18567 272555 18579 272589
rect 17579 272543 18579 272555
rect 17579 272431 18579 272443
rect 17579 272397 17591 272431
rect 18567 272397 18579 272431
rect 17579 272385 18579 272397
rect 17579 272273 18579 272285
rect 17579 272239 17591 272273
rect 18567 272239 18579 272273
rect 17579 272227 18579 272239
rect 17579 272115 18579 272127
rect 17579 272081 17591 272115
rect 18567 272081 18579 272115
rect 17579 272069 18579 272081
rect 19099 273221 20099 273233
rect 19099 273187 19111 273221
rect 20087 273187 20099 273221
rect 19099 273175 20099 273187
rect 19099 273063 20099 273075
rect 19099 273029 19111 273063
rect 20087 273029 20099 273063
rect 19099 273017 20099 273029
rect 19099 272905 20099 272917
rect 19099 272871 19111 272905
rect 20087 272871 20099 272905
rect 19099 272859 20099 272871
rect 19099 272747 20099 272759
rect 19099 272713 19111 272747
rect 20087 272713 20099 272747
rect 19099 272701 20099 272713
rect 19099 272589 20099 272601
rect 19099 272555 19111 272589
rect 20087 272555 20099 272589
rect 19099 272543 20099 272555
rect 19099 272431 20099 272443
rect 19099 272397 19111 272431
rect 20087 272397 20099 272431
rect 19099 272385 20099 272397
rect 19099 272273 20099 272285
rect 19099 272239 19111 272273
rect 20087 272239 20099 272273
rect 19099 272227 20099 272239
rect 19099 272115 20099 272127
rect 19099 272081 19111 272115
rect 20087 272081 20099 272115
rect 19099 272069 20099 272081
rect 20620 274220 21620 274232
rect 20620 274186 20632 274220
rect 21608 274186 21620 274220
rect 20620 274174 21620 274186
rect 20620 273962 21620 273974
rect 20620 273928 20632 273962
rect 21608 273928 21620 273962
rect 20620 273916 21620 273928
rect 20620 273704 21620 273716
rect 20620 273670 20632 273704
rect 21608 273670 21620 273704
rect 20620 273658 21620 273670
rect 20620 273446 21620 273458
rect 20620 273412 20632 273446
rect 21608 273412 21620 273446
rect 20620 273400 21620 273412
rect 20620 273188 21620 273200
rect 20620 273154 20632 273188
rect 21608 273154 21620 273188
rect 20620 273142 21620 273154
rect 20620 272930 21620 272942
rect 20620 272896 20632 272930
rect 21608 272896 21620 272930
rect 20620 272884 21620 272896
rect 20620 272672 21620 272684
rect 20620 272638 20632 272672
rect 21608 272638 21620 272672
rect 20620 272626 21620 272638
rect 20620 272414 21620 272426
rect 20620 272380 20632 272414
rect 21608 272380 21620 272414
rect 20620 272368 21620 272380
rect 20620 272156 21620 272168
rect 20620 272122 20632 272156
rect 21608 272122 21620 272156
rect 20620 272110 21620 272122
rect 20620 271898 21620 271910
rect 20620 271864 20632 271898
rect 21608 271864 21620 271898
rect 20620 271852 21620 271864
rect 20620 271640 21620 271652
rect 20620 271606 20632 271640
rect 21608 271606 21620 271640
rect 20620 271594 21620 271606
rect 20620 271382 21620 271394
rect 20620 271348 20632 271382
rect 21608 271348 21620 271382
rect 20620 271336 21620 271348
rect 20620 271124 21620 271136
rect 20620 271090 20632 271124
rect 21608 271090 21620 271124
rect 20620 271078 21620 271090
rect 22140 274476 23140 274488
rect 22140 274442 22152 274476
rect 23128 274442 23140 274476
rect 22140 274430 23140 274442
rect 22140 274218 23140 274230
rect 22140 274184 22152 274218
rect 23128 274184 23140 274218
rect 22140 274172 23140 274184
rect 22140 273960 23140 273972
rect 22140 273926 22152 273960
rect 23128 273926 23140 273960
rect 22140 273914 23140 273926
rect 22140 273702 23140 273714
rect 22140 273668 22152 273702
rect 23128 273668 23140 273702
rect 22140 273656 23140 273668
rect 22140 273444 23140 273456
rect 22140 273410 22152 273444
rect 23128 273410 23140 273444
rect 22140 273398 23140 273410
rect 22140 273186 23140 273198
rect 22140 273152 22152 273186
rect 23128 273152 23140 273186
rect 22140 273140 23140 273152
rect 22140 272928 23140 272940
rect 22140 272894 22152 272928
rect 23128 272894 23140 272928
rect 22140 272882 23140 272894
rect 22140 272670 23140 272682
rect 22140 272636 22152 272670
rect 23128 272636 23140 272670
rect 22140 272624 23140 272636
rect 22140 272412 23140 272424
rect 22140 272378 22152 272412
rect 23128 272378 23140 272412
rect 22140 272366 23140 272378
rect 22140 272154 23140 272166
rect 22140 272120 22152 272154
rect 23128 272120 23140 272154
rect 22140 272108 23140 272120
rect 22140 271896 23140 271908
rect 22140 271862 22152 271896
rect 23128 271862 23140 271896
rect 22140 271850 23140 271862
rect 22140 271638 23140 271650
rect 22140 271604 22152 271638
rect 23128 271604 23140 271638
rect 22140 271592 23140 271604
rect 22140 271380 23140 271392
rect 22140 271346 22152 271380
rect 23128 271346 23140 271380
rect 22140 271334 23140 271346
rect 22140 271122 23140 271134
rect 22140 271088 22152 271122
rect 23128 271088 23140 271122
rect 22140 271076 23140 271088
rect 22140 270864 23140 270876
rect 22140 270830 22152 270864
rect 23128 270830 23140 270864
rect 22140 270818 23140 270830
rect 27290 272810 27790 272822
rect 27290 272776 27302 272810
rect 27778 272776 27790 272810
rect 27290 272764 27790 272776
rect 27290 272652 27790 272664
rect 27290 272618 27302 272652
rect 27778 272618 27790 272652
rect 27290 272606 27790 272618
rect 27290 272494 27790 272506
rect 27290 272460 27302 272494
rect 27778 272460 27790 272494
rect 27290 272448 27790 272460
rect 28290 273166 28540 273178
rect 28290 273132 28302 273166
rect 28528 273132 28540 273166
rect 28290 273120 28540 273132
rect 28290 272908 28540 272920
rect 28290 272874 28302 272908
rect 28528 272874 28540 272908
rect 28290 272862 28540 272874
rect 28290 272650 28540 272662
rect 28290 272616 28302 272650
rect 28528 272616 28540 272650
rect 28290 272604 28540 272616
rect 28290 272392 28540 272404
rect 28290 272358 28302 272392
rect 28528 272358 28540 272392
rect 28290 272346 28540 272358
rect 28290 272134 28540 272146
rect 28290 272100 28302 272134
rect 28528 272100 28540 272134
rect 28290 272088 28540 272100
rect 29040 273427 30040 273439
rect 29040 273393 29052 273427
rect 30028 273393 30040 273427
rect 29040 273381 30040 273393
rect 29040 273169 30040 273181
rect 29040 273135 29052 273169
rect 30028 273135 30040 273169
rect 29040 273123 30040 273135
rect 29040 272911 30040 272923
rect 29040 272877 29052 272911
rect 30028 272877 30040 272911
rect 29040 272865 30040 272877
rect 29040 272653 30040 272665
rect 29040 272619 29052 272653
rect 30028 272619 30040 272653
rect 29040 272607 30040 272619
rect 29040 272395 30040 272407
rect 29040 272361 29052 272395
rect 30028 272361 30040 272395
rect 29040 272349 30040 272361
rect 29040 272137 30040 272149
rect 29040 272103 29052 272137
rect 30028 272103 30040 272137
rect 29040 272091 30040 272103
rect 29040 271879 30040 271891
rect 29040 271845 29052 271879
rect 30028 271845 30040 271879
rect 29040 271833 30040 271845
rect 5990 252364 15990 252376
rect 5990 252330 6002 252364
rect 15978 252330 15990 252364
rect 5990 252318 15990 252330
rect 5990 252266 15990 252278
rect 5990 252232 6002 252266
rect 15978 252232 15990 252266
rect 5990 252220 15990 252232
rect 5990 252168 15990 252180
rect 5990 252134 6002 252168
rect 15978 252134 15990 252168
rect 5990 252122 15990 252134
rect 5990 252070 15990 252082
rect 5990 252036 6002 252070
rect 15978 252036 15990 252070
rect 5990 252024 15990 252036
rect 5990 251972 15990 251984
rect 5990 251938 6002 251972
rect 15978 251938 15990 251972
rect 5990 251926 15990 251938
rect 5990 251874 15990 251886
rect 5990 251840 6002 251874
rect 15978 251840 15990 251874
rect 5990 251828 15990 251840
rect 5990 251776 15990 251788
rect 5990 251742 6002 251776
rect 15978 251742 15990 251776
rect 5990 251730 15990 251742
rect 5990 251678 15990 251690
rect 5990 251644 6002 251678
rect 15978 251644 15990 251678
rect 5990 251632 15990 251644
rect 5990 251580 15990 251592
rect 5990 251546 6002 251580
rect 15978 251546 15990 251580
rect 5990 251534 15990 251546
rect 5990 251482 15990 251494
rect 5990 251448 6002 251482
rect 15978 251448 15990 251482
rect 5990 251436 15990 251448
rect 5990 251384 15990 251396
rect 5990 251350 6002 251384
rect 15978 251350 15990 251384
rect 5990 251338 15990 251350
rect 5990 241964 15990 241976
rect 5990 241930 6002 241964
rect 15978 241930 15990 241964
rect 5990 241918 15990 241930
rect 5990 241866 15990 241878
rect 5990 241832 6002 241866
rect 15978 241832 15990 241866
rect 5990 241820 15990 241832
rect 5990 241768 15990 241780
rect 5990 241734 6002 241768
rect 15978 241734 15990 241768
rect 5990 241722 15990 241734
rect 5990 241670 15990 241682
rect 5990 241636 6002 241670
rect 15978 241636 15990 241670
rect 5990 241624 15990 241636
rect 5990 241572 15990 241584
rect 5990 241538 6002 241572
rect 15978 241538 15990 241572
rect 5990 241526 15990 241538
rect 5990 241474 15990 241486
rect 5990 241440 6002 241474
rect 15978 241440 15990 241474
rect 5990 241428 15990 241440
rect 5990 241376 15990 241388
rect 5990 241342 6002 241376
rect 15978 241342 15990 241376
rect 5990 241330 15990 241342
rect 5990 241278 15990 241290
rect 5990 241244 6002 241278
rect 15978 241244 15990 241278
rect 5990 241232 15990 241244
rect 5990 241180 15990 241192
rect 5990 241146 6002 241180
rect 15978 241146 15990 241180
rect 5990 241134 15990 241146
rect 5990 241082 15990 241094
rect 5990 241048 6002 241082
rect 15978 241048 15990 241082
rect 5990 241036 15990 241048
rect 5990 240984 15990 240996
rect 5990 240950 6002 240984
rect 15978 240950 15990 240984
rect 5990 240938 15990 240950
<< pdiff >>
rect 536368 294784 537368 294796
rect 536368 294750 536380 294784
rect 537356 294750 537368 294784
rect 536368 294738 537368 294750
rect 537604 294784 538604 294796
rect 537604 294750 537616 294784
rect 538592 294750 538604 294784
rect 537604 294738 538604 294750
rect 538840 294784 539840 294796
rect 538840 294750 538852 294784
rect 539828 294750 539840 294784
rect 538840 294738 539840 294750
rect 540076 294784 541076 294796
rect 540076 294750 540088 294784
rect 541064 294750 541076 294784
rect 540076 294738 541076 294750
rect 541312 294784 542312 294796
rect 541312 294750 541324 294784
rect 542300 294750 542312 294784
rect 541312 294738 542312 294750
rect 542548 294784 543548 294796
rect 542548 294750 542560 294784
rect 543536 294750 543548 294784
rect 542548 294738 543548 294750
rect 543784 294784 544784 294796
rect 543784 294750 543796 294784
rect 544772 294750 544784 294784
rect 543784 294738 544784 294750
rect 536368 294626 537368 294638
rect 536368 294592 536380 294626
rect 537356 294592 537368 294626
rect 536368 294580 537368 294592
rect 537604 294626 538604 294638
rect 537604 294592 537616 294626
rect 538592 294592 538604 294626
rect 537604 294580 538604 294592
rect 538840 294626 539840 294638
rect 538840 294592 538852 294626
rect 539828 294592 539840 294626
rect 538840 294580 539840 294592
rect 540076 294626 541076 294638
rect 540076 294592 540088 294626
rect 541064 294592 541076 294626
rect 540076 294580 541076 294592
rect 541312 294626 542312 294638
rect 541312 294592 541324 294626
rect 542300 294592 542312 294626
rect 541312 294580 542312 294592
rect 542548 294626 543548 294638
rect 542548 294592 542560 294626
rect 543536 294592 543548 294626
rect 542548 294580 543548 294592
rect 543784 294626 544784 294638
rect 543784 294592 543796 294626
rect 544772 294592 544784 294626
rect 543784 294580 544784 294592
rect 536368 294244 537368 294256
rect 536368 294210 536380 294244
rect 537356 294210 537368 294244
rect 536368 294198 537368 294210
rect 537604 294244 538604 294256
rect 537604 294210 537616 294244
rect 538592 294210 538604 294244
rect 537604 294198 538604 294210
rect 538840 294244 539840 294256
rect 538840 294210 538852 294244
rect 539828 294210 539840 294244
rect 538840 294198 539840 294210
rect 540076 294244 541076 294256
rect 540076 294210 540088 294244
rect 541064 294210 541076 294244
rect 540076 294198 541076 294210
rect 541312 294244 542312 294256
rect 541312 294210 541324 294244
rect 542300 294210 542312 294244
rect 541312 294198 542312 294210
rect 542548 294244 543548 294256
rect 542548 294210 542560 294244
rect 543536 294210 543548 294244
rect 542548 294198 543548 294210
rect 543784 294244 544784 294256
rect 543784 294210 543796 294244
rect 544772 294210 544784 294244
rect 543784 294198 544784 294210
rect 536368 294086 537368 294098
rect 536368 294052 536380 294086
rect 537356 294052 537368 294086
rect 536368 294040 537368 294052
rect 537604 294086 538604 294098
rect 537604 294052 537616 294086
rect 538592 294052 538604 294086
rect 537604 294040 538604 294052
rect 538840 294086 539840 294098
rect 538840 294052 538852 294086
rect 539828 294052 539840 294086
rect 538840 294040 539840 294052
rect 540076 294086 541076 294098
rect 540076 294052 540088 294086
rect 541064 294052 541076 294086
rect 540076 294040 541076 294052
rect 541312 294086 542312 294098
rect 541312 294052 541324 294086
rect 542300 294052 542312 294086
rect 541312 294040 542312 294052
rect 542548 294086 543548 294098
rect 542548 294052 542560 294086
rect 543536 294052 543548 294086
rect 542548 294040 543548 294052
rect 543784 294086 544784 294098
rect 543784 294052 543796 294086
rect 544772 294052 544784 294086
rect 543784 294040 544784 294052
rect 536368 293704 537368 293716
rect 536368 293670 536380 293704
rect 537356 293670 537368 293704
rect 536368 293658 537368 293670
rect 537604 293704 538604 293716
rect 537604 293670 537616 293704
rect 538592 293670 538604 293704
rect 537604 293658 538604 293670
rect 538840 293704 539840 293716
rect 538840 293670 538852 293704
rect 539828 293670 539840 293704
rect 538840 293658 539840 293670
rect 540076 293704 541076 293716
rect 540076 293670 540088 293704
rect 541064 293670 541076 293704
rect 540076 293658 541076 293670
rect 541312 293704 542312 293716
rect 541312 293670 541324 293704
rect 542300 293670 542312 293704
rect 541312 293658 542312 293670
rect 542548 293704 543548 293716
rect 542548 293670 542560 293704
rect 543536 293670 543548 293704
rect 542548 293658 543548 293670
rect 543784 293704 544784 293716
rect 543784 293670 543796 293704
rect 544772 293670 544784 293704
rect 543784 293658 544784 293670
rect 536368 293546 537368 293558
rect 536368 293512 536380 293546
rect 537356 293512 537368 293546
rect 536368 293500 537368 293512
rect 537604 293546 538604 293558
rect 537604 293512 537616 293546
rect 538592 293512 538604 293546
rect 537604 293500 538604 293512
rect 538840 293546 539840 293558
rect 538840 293512 538852 293546
rect 539828 293512 539840 293546
rect 538840 293500 539840 293512
rect 540076 293546 541076 293558
rect 540076 293512 540088 293546
rect 541064 293512 541076 293546
rect 540076 293500 541076 293512
rect 541312 293546 542312 293558
rect 541312 293512 541324 293546
rect 542300 293512 542312 293546
rect 541312 293500 542312 293512
rect 542548 293546 543548 293558
rect 542548 293512 542560 293546
rect 543536 293512 543548 293546
rect 542548 293500 543548 293512
rect 543784 293546 544784 293558
rect 543784 293512 543796 293546
rect 544772 293512 544784 293546
rect 543784 293500 544784 293512
rect 536368 293164 537368 293176
rect 536368 293130 536380 293164
rect 537356 293130 537368 293164
rect 536368 293118 537368 293130
rect 537604 293164 538604 293176
rect 537604 293130 537616 293164
rect 538592 293130 538604 293164
rect 537604 293118 538604 293130
rect 538840 293164 539840 293176
rect 538840 293130 538852 293164
rect 539828 293130 539840 293164
rect 538840 293118 539840 293130
rect 540076 293164 541076 293176
rect 540076 293130 540088 293164
rect 541064 293130 541076 293164
rect 540076 293118 541076 293130
rect 541312 293164 542312 293176
rect 541312 293130 541324 293164
rect 542300 293130 542312 293164
rect 541312 293118 542312 293130
rect 542548 293164 543548 293176
rect 542548 293130 542560 293164
rect 543536 293130 543548 293164
rect 542548 293118 543548 293130
rect 543784 293164 544784 293176
rect 543784 293130 543796 293164
rect 544772 293130 544784 293164
rect 543784 293118 544784 293130
rect 536368 293006 537368 293018
rect 536368 292972 536380 293006
rect 537356 292972 537368 293006
rect 536368 292960 537368 292972
rect 537604 293006 538604 293018
rect 537604 292972 537616 293006
rect 538592 292972 538604 293006
rect 537604 292960 538604 292972
rect 538840 293006 539840 293018
rect 538840 292972 538852 293006
rect 539828 292972 539840 293006
rect 538840 292960 539840 292972
rect 540076 293006 541076 293018
rect 540076 292972 540088 293006
rect 541064 292972 541076 293006
rect 540076 292960 541076 292972
rect 541312 293006 542312 293018
rect 541312 292972 541324 293006
rect 542300 292972 542312 293006
rect 541312 292960 542312 292972
rect 542548 293006 543548 293018
rect 542548 292972 542560 293006
rect 543536 292972 543548 293006
rect 542548 292960 543548 292972
rect 543784 293006 544784 293018
rect 543784 292972 543796 293006
rect 544772 292972 544784 293006
rect 543784 292960 544784 292972
rect 536368 292584 537368 292596
rect 536368 292550 536380 292584
rect 537356 292550 537368 292584
rect 536368 292538 537368 292550
rect 537604 292584 538604 292596
rect 537604 292550 537616 292584
rect 538592 292550 538604 292584
rect 537604 292538 538604 292550
rect 538840 292584 539840 292596
rect 538840 292550 538852 292584
rect 539828 292550 539840 292584
rect 538840 292538 539840 292550
rect 540076 292584 541076 292596
rect 540076 292550 540088 292584
rect 541064 292550 541076 292584
rect 540076 292538 541076 292550
rect 541312 292584 542312 292596
rect 541312 292550 541324 292584
rect 542300 292550 542312 292584
rect 541312 292538 542312 292550
rect 542548 292584 543548 292596
rect 542548 292550 542560 292584
rect 543536 292550 543548 292584
rect 542548 292538 543548 292550
rect 543784 292584 544784 292596
rect 543784 292550 543796 292584
rect 544772 292550 544784 292584
rect 543784 292538 544784 292550
rect 536368 292426 537368 292438
rect 536368 292392 536380 292426
rect 537356 292392 537368 292426
rect 536368 292380 537368 292392
rect 537604 292426 538604 292438
rect 537604 292392 537616 292426
rect 538592 292392 538604 292426
rect 537604 292380 538604 292392
rect 538840 292426 539840 292438
rect 538840 292392 538852 292426
rect 539828 292392 539840 292426
rect 538840 292380 539840 292392
rect 540076 292426 541076 292438
rect 540076 292392 540088 292426
rect 541064 292392 541076 292426
rect 540076 292380 541076 292392
rect 541312 292426 542312 292438
rect 541312 292392 541324 292426
rect 542300 292392 542312 292426
rect 541312 292380 542312 292392
rect 542548 292426 543548 292438
rect 542548 292392 542560 292426
rect 543536 292392 543548 292426
rect 542548 292380 543548 292392
rect 543784 292426 544784 292438
rect 543784 292392 543796 292426
rect 544772 292392 544784 292426
rect 543784 292380 544784 292392
rect 536368 292004 537368 292016
rect 536368 291970 536380 292004
rect 537356 291970 537368 292004
rect 536368 291958 537368 291970
rect 537604 292004 538604 292016
rect 537604 291970 537616 292004
rect 538592 291970 538604 292004
rect 537604 291958 538604 291970
rect 538840 292004 539840 292016
rect 538840 291970 538852 292004
rect 539828 291970 539840 292004
rect 538840 291958 539840 291970
rect 540076 292004 541076 292016
rect 540076 291970 540088 292004
rect 541064 291970 541076 292004
rect 540076 291958 541076 291970
rect 541312 292004 542312 292016
rect 541312 291970 541324 292004
rect 542300 291970 542312 292004
rect 541312 291958 542312 291970
rect 542548 292004 543548 292016
rect 542548 291970 542560 292004
rect 543536 291970 543548 292004
rect 542548 291958 543548 291970
rect 543784 292004 544784 292016
rect 543784 291970 543796 292004
rect 544772 291970 544784 292004
rect 543784 291958 544784 291970
rect 536368 291846 537368 291858
rect 536368 291812 536380 291846
rect 537356 291812 537368 291846
rect 536368 291800 537368 291812
rect 537604 291846 538604 291858
rect 537604 291812 537616 291846
rect 538592 291812 538604 291846
rect 537604 291800 538604 291812
rect 538840 291846 539840 291858
rect 538840 291812 538852 291846
rect 539828 291812 539840 291846
rect 538840 291800 539840 291812
rect 540076 291846 541076 291858
rect 540076 291812 540088 291846
rect 541064 291812 541076 291846
rect 540076 291800 541076 291812
rect 541312 291846 542312 291858
rect 541312 291812 541324 291846
rect 542300 291812 542312 291846
rect 541312 291800 542312 291812
rect 542548 291846 543548 291858
rect 542548 291812 542560 291846
rect 543536 291812 543548 291846
rect 542548 291800 543548 291812
rect 543784 291846 544784 291858
rect 543784 291812 543796 291846
rect 544772 291812 544784 291846
rect 543784 291800 544784 291812
rect 534528 291464 535528 291476
rect 534528 291430 534540 291464
rect 535516 291430 535528 291464
rect 534528 291418 535528 291430
rect 535764 291464 536764 291476
rect 535764 291430 535776 291464
rect 536752 291430 536764 291464
rect 535764 291418 536764 291430
rect 537000 291464 538000 291476
rect 537000 291430 537012 291464
rect 537988 291430 538000 291464
rect 537000 291418 538000 291430
rect 538236 291464 539236 291476
rect 538236 291430 538248 291464
rect 539224 291430 539236 291464
rect 538236 291418 539236 291430
rect 539472 291464 540472 291476
rect 539472 291430 539484 291464
rect 540460 291430 540472 291464
rect 539472 291418 540472 291430
rect 540708 291464 541708 291476
rect 540708 291430 540720 291464
rect 541696 291430 541708 291464
rect 540708 291418 541708 291430
rect 541944 291464 542944 291476
rect 541944 291430 541956 291464
rect 542932 291430 542944 291464
rect 541944 291418 542944 291430
rect 543180 291464 544180 291476
rect 543180 291430 543192 291464
rect 544168 291430 544180 291464
rect 543180 291418 544180 291430
rect 544416 291464 545416 291476
rect 544416 291430 544428 291464
rect 545404 291430 545416 291464
rect 544416 291418 545416 291430
rect 545652 291464 546652 291476
rect 545652 291430 545664 291464
rect 546640 291430 546652 291464
rect 545652 291418 546652 291430
rect 534528 291306 535528 291318
rect 534528 291272 534540 291306
rect 535516 291272 535528 291306
rect 534528 291260 535528 291272
rect 535764 291306 536764 291318
rect 535764 291272 535776 291306
rect 536752 291272 536764 291306
rect 535764 291260 536764 291272
rect 537000 291306 538000 291318
rect 537000 291272 537012 291306
rect 537988 291272 538000 291306
rect 537000 291260 538000 291272
rect 538236 291306 539236 291318
rect 538236 291272 538248 291306
rect 539224 291272 539236 291306
rect 538236 291260 539236 291272
rect 539472 291306 540472 291318
rect 539472 291272 539484 291306
rect 540460 291272 540472 291306
rect 539472 291260 540472 291272
rect 540708 291306 541708 291318
rect 540708 291272 540720 291306
rect 541696 291272 541708 291306
rect 540708 291260 541708 291272
rect 541944 291306 542944 291318
rect 541944 291272 541956 291306
rect 542932 291272 542944 291306
rect 541944 291260 542944 291272
rect 543180 291306 544180 291318
rect 543180 291272 543192 291306
rect 544168 291272 544180 291306
rect 543180 291260 544180 291272
rect 544416 291306 545416 291318
rect 544416 291272 544428 291306
rect 545404 291272 545416 291306
rect 544416 291260 545416 291272
rect 545652 291306 546652 291318
rect 545652 291272 545664 291306
rect 546640 291272 546652 291306
rect 545652 291260 546652 291272
rect 534528 290924 535528 290936
rect 534528 290890 534540 290924
rect 535516 290890 535528 290924
rect 534528 290878 535528 290890
rect 535764 290924 536764 290936
rect 535764 290890 535776 290924
rect 536752 290890 536764 290924
rect 535764 290878 536764 290890
rect 537000 290924 538000 290936
rect 537000 290890 537012 290924
rect 537988 290890 538000 290924
rect 537000 290878 538000 290890
rect 538236 290924 539236 290936
rect 538236 290890 538248 290924
rect 539224 290890 539236 290924
rect 538236 290878 539236 290890
rect 539472 290924 540472 290936
rect 539472 290890 539484 290924
rect 540460 290890 540472 290924
rect 539472 290878 540472 290890
rect 540708 290924 541708 290936
rect 540708 290890 540720 290924
rect 541696 290890 541708 290924
rect 540708 290878 541708 290890
rect 541944 290924 542944 290936
rect 541944 290890 541956 290924
rect 542932 290890 542944 290924
rect 541944 290878 542944 290890
rect 543180 290924 544180 290936
rect 543180 290890 543192 290924
rect 544168 290890 544180 290924
rect 543180 290878 544180 290890
rect 544416 290924 545416 290936
rect 544416 290890 544428 290924
rect 545404 290890 545416 290924
rect 544416 290878 545416 290890
rect 545652 290924 546652 290936
rect 545652 290890 545664 290924
rect 546640 290890 546652 290924
rect 545652 290878 546652 290890
rect 534528 290766 535528 290778
rect 534528 290732 534540 290766
rect 535516 290732 535528 290766
rect 534528 290720 535528 290732
rect 535764 290766 536764 290778
rect 535764 290732 535776 290766
rect 536752 290732 536764 290766
rect 535764 290720 536764 290732
rect 537000 290766 538000 290778
rect 537000 290732 537012 290766
rect 537988 290732 538000 290766
rect 537000 290720 538000 290732
rect 538236 290766 539236 290778
rect 538236 290732 538248 290766
rect 539224 290732 539236 290766
rect 538236 290720 539236 290732
rect 539472 290766 540472 290778
rect 539472 290732 539484 290766
rect 540460 290732 540472 290766
rect 539472 290720 540472 290732
rect 540708 290766 541708 290778
rect 540708 290732 540720 290766
rect 541696 290732 541708 290766
rect 540708 290720 541708 290732
rect 541944 290766 542944 290778
rect 541944 290732 541956 290766
rect 542932 290732 542944 290766
rect 541944 290720 542944 290732
rect 543180 290766 544180 290778
rect 543180 290732 543192 290766
rect 544168 290732 544180 290766
rect 543180 290720 544180 290732
rect 544416 290766 545416 290778
rect 544416 290732 544428 290766
rect 545404 290732 545416 290766
rect 544416 290720 545416 290732
rect 545652 290766 546652 290778
rect 545652 290732 545664 290766
rect 546640 290732 546652 290766
rect 545652 290720 546652 290732
rect 534528 290384 535528 290396
rect 534528 290350 534540 290384
rect 535516 290350 535528 290384
rect 534528 290338 535528 290350
rect 535764 290384 536764 290396
rect 535764 290350 535776 290384
rect 536752 290350 536764 290384
rect 535764 290338 536764 290350
rect 537000 290384 538000 290396
rect 537000 290350 537012 290384
rect 537988 290350 538000 290384
rect 537000 290338 538000 290350
rect 538236 290384 539236 290396
rect 538236 290350 538248 290384
rect 539224 290350 539236 290384
rect 538236 290338 539236 290350
rect 539472 290384 540472 290396
rect 539472 290350 539484 290384
rect 540460 290350 540472 290384
rect 539472 290338 540472 290350
rect 540708 290384 541708 290396
rect 540708 290350 540720 290384
rect 541696 290350 541708 290384
rect 540708 290338 541708 290350
rect 541944 290384 542944 290396
rect 541944 290350 541956 290384
rect 542932 290350 542944 290384
rect 541944 290338 542944 290350
rect 543180 290384 544180 290396
rect 543180 290350 543192 290384
rect 544168 290350 544180 290384
rect 543180 290338 544180 290350
rect 544416 290384 545416 290396
rect 544416 290350 544428 290384
rect 545404 290350 545416 290384
rect 544416 290338 545416 290350
rect 545652 290384 546652 290396
rect 545652 290350 545664 290384
rect 546640 290350 546652 290384
rect 545652 290338 546652 290350
rect 534528 290226 535528 290238
rect 534528 290192 534540 290226
rect 535516 290192 535528 290226
rect 534528 290180 535528 290192
rect 535764 290226 536764 290238
rect 535764 290192 535776 290226
rect 536752 290192 536764 290226
rect 535764 290180 536764 290192
rect 537000 290226 538000 290238
rect 537000 290192 537012 290226
rect 537988 290192 538000 290226
rect 537000 290180 538000 290192
rect 538236 290226 539236 290238
rect 538236 290192 538248 290226
rect 539224 290192 539236 290226
rect 538236 290180 539236 290192
rect 539472 290226 540472 290238
rect 539472 290192 539484 290226
rect 540460 290192 540472 290226
rect 539472 290180 540472 290192
rect 540708 290226 541708 290238
rect 540708 290192 540720 290226
rect 541696 290192 541708 290226
rect 540708 290180 541708 290192
rect 541944 290226 542944 290238
rect 541944 290192 541956 290226
rect 542932 290192 542944 290226
rect 541944 290180 542944 290192
rect 543180 290226 544180 290238
rect 543180 290192 543192 290226
rect 544168 290192 544180 290226
rect 543180 290180 544180 290192
rect 544416 290226 545416 290238
rect 544416 290192 544428 290226
rect 545404 290192 545416 290226
rect 544416 290180 545416 290192
rect 545652 290226 546652 290238
rect 545652 290192 545664 290226
rect 546640 290192 546652 290226
rect 545652 290180 546652 290192
rect 534528 289844 535528 289856
rect 534528 289810 534540 289844
rect 535516 289810 535528 289844
rect 534528 289798 535528 289810
rect 535764 289844 536764 289856
rect 535764 289810 535776 289844
rect 536752 289810 536764 289844
rect 535764 289798 536764 289810
rect 537000 289844 538000 289856
rect 537000 289810 537012 289844
rect 537988 289810 538000 289844
rect 537000 289798 538000 289810
rect 538236 289844 539236 289856
rect 538236 289810 538248 289844
rect 539224 289810 539236 289844
rect 538236 289798 539236 289810
rect 539472 289844 540472 289856
rect 539472 289810 539484 289844
rect 540460 289810 540472 289844
rect 539472 289798 540472 289810
rect 540708 289844 541708 289856
rect 540708 289810 540720 289844
rect 541696 289810 541708 289844
rect 540708 289798 541708 289810
rect 541944 289844 542944 289856
rect 541944 289810 541956 289844
rect 542932 289810 542944 289844
rect 541944 289798 542944 289810
rect 543180 289844 544180 289856
rect 543180 289810 543192 289844
rect 544168 289810 544180 289844
rect 543180 289798 544180 289810
rect 544416 289844 545416 289856
rect 544416 289810 544428 289844
rect 545404 289810 545416 289844
rect 544416 289798 545416 289810
rect 545652 289844 546652 289856
rect 545652 289810 545664 289844
rect 546640 289810 546652 289844
rect 545652 289798 546652 289810
rect 534528 289686 535528 289698
rect 534528 289652 534540 289686
rect 535516 289652 535528 289686
rect 534528 289640 535528 289652
rect 535764 289686 536764 289698
rect 535764 289652 535776 289686
rect 536752 289652 536764 289686
rect 535764 289640 536764 289652
rect 537000 289686 538000 289698
rect 537000 289652 537012 289686
rect 537988 289652 538000 289686
rect 537000 289640 538000 289652
rect 538236 289686 539236 289698
rect 538236 289652 538248 289686
rect 539224 289652 539236 289686
rect 538236 289640 539236 289652
rect 539472 289686 540472 289698
rect 539472 289652 539484 289686
rect 540460 289652 540472 289686
rect 539472 289640 540472 289652
rect 540708 289686 541708 289698
rect 540708 289652 540720 289686
rect 541696 289652 541708 289686
rect 540708 289640 541708 289652
rect 541944 289686 542944 289698
rect 541944 289652 541956 289686
rect 542932 289652 542944 289686
rect 541944 289640 542944 289652
rect 543180 289686 544180 289698
rect 543180 289652 543192 289686
rect 544168 289652 544180 289686
rect 543180 289640 544180 289652
rect 544416 289686 545416 289698
rect 544416 289652 544428 289686
rect 545404 289652 545416 289686
rect 544416 289640 545416 289652
rect 545652 289686 546652 289698
rect 545652 289652 545664 289686
rect 546640 289652 546652 289686
rect 545652 289640 546652 289652
rect 537013 285270 538013 285282
rect 537013 285236 537025 285270
rect 538001 285236 538013 285270
rect 537013 285224 538013 285236
rect 538249 285270 539249 285282
rect 538249 285236 538261 285270
rect 539237 285236 539249 285270
rect 538249 285224 539249 285236
rect 539485 285270 540485 285282
rect 539485 285236 539497 285270
rect 540473 285236 540485 285270
rect 539485 285224 540485 285236
rect 540721 285270 541721 285282
rect 540721 285236 540733 285270
rect 541709 285236 541721 285270
rect 540721 285224 541721 285236
rect 541957 285270 542957 285282
rect 541957 285236 541969 285270
rect 542945 285236 542957 285270
rect 541957 285224 542957 285236
rect 543193 285270 544193 285282
rect 543193 285236 543205 285270
rect 544181 285236 544193 285270
rect 543193 285224 544193 285236
rect 537013 285012 538013 285024
rect 537013 284978 537025 285012
rect 538001 284978 538013 285012
rect 537013 284966 538013 284978
rect 538249 285012 539249 285024
rect 538249 284978 538261 285012
rect 539237 284978 539249 285012
rect 538249 284966 539249 284978
rect 539485 285012 540485 285024
rect 539485 284978 539497 285012
rect 540473 284978 540485 285012
rect 539485 284966 540485 284978
rect 540721 285012 541721 285024
rect 540721 284978 540733 285012
rect 541709 284978 541721 285012
rect 540721 284966 541721 284978
rect 541957 285012 542957 285024
rect 541957 284978 541969 285012
rect 542945 284978 542957 285012
rect 541957 284966 542957 284978
rect 543193 285012 544193 285024
rect 543193 284978 543205 285012
rect 544181 284978 544193 285012
rect 543193 284966 544193 284978
rect 537013 284680 538013 284692
rect 537013 284646 537025 284680
rect 538001 284646 538013 284680
rect 537013 284634 538013 284646
rect 538249 284680 539249 284692
rect 538249 284646 538261 284680
rect 539237 284646 539249 284680
rect 538249 284634 539249 284646
rect 539485 284680 540485 284692
rect 539485 284646 539497 284680
rect 540473 284646 540485 284680
rect 539485 284634 540485 284646
rect 540721 284680 541721 284692
rect 540721 284646 540733 284680
rect 541709 284646 541721 284680
rect 540721 284634 541721 284646
rect 541957 284680 542957 284692
rect 541957 284646 541969 284680
rect 542945 284646 542957 284680
rect 541957 284634 542957 284646
rect 543193 284680 544193 284692
rect 543193 284646 543205 284680
rect 544181 284646 544193 284680
rect 543193 284634 544193 284646
rect 537013 284422 538013 284434
rect 537013 284388 537025 284422
rect 538001 284388 538013 284422
rect 537013 284376 538013 284388
rect 538249 284422 539249 284434
rect 538249 284388 538261 284422
rect 539237 284388 539249 284422
rect 538249 284376 539249 284388
rect 539485 284422 540485 284434
rect 539485 284388 539497 284422
rect 540473 284388 540485 284422
rect 539485 284376 540485 284388
rect 540721 284422 541721 284434
rect 540721 284388 540733 284422
rect 541709 284388 541721 284422
rect 540721 284376 541721 284388
rect 541957 284422 542957 284434
rect 541957 284388 541969 284422
rect 542945 284388 542957 284422
rect 541957 284376 542957 284388
rect 543193 284422 544193 284434
rect 543193 284388 543205 284422
rect 544181 284388 544193 284422
rect 543193 284376 544193 284388
rect 12801 275834 13801 275846
rect 12801 275800 12813 275834
rect 13789 275800 13801 275834
rect 12801 275788 13801 275800
rect 12801 275676 13801 275688
rect 12801 275642 12813 275676
rect 13789 275642 13801 275676
rect 12801 275630 13801 275642
rect 12801 275518 13801 275530
rect 12801 275484 12813 275518
rect 13789 275484 13801 275518
rect 12801 275472 13801 275484
rect 12801 275360 13801 275372
rect 12801 275326 12813 275360
rect 13789 275326 13801 275360
rect 12801 275314 13801 275326
rect 12801 275202 13801 275214
rect 12801 275168 12813 275202
rect 13789 275168 13801 275202
rect 12801 275156 13801 275168
rect 12801 275044 13801 275056
rect 12801 275010 12813 275044
rect 13789 275010 13801 275044
rect 12801 274998 13801 275010
rect 12801 274886 13801 274898
rect 12801 274852 12813 274886
rect 13789 274852 13801 274886
rect 12801 274840 13801 274852
rect 12801 274728 13801 274740
rect 12801 274694 12813 274728
rect 13789 274694 13801 274728
rect 12801 274682 13801 274694
rect 12801 274570 13801 274582
rect 12801 274536 12813 274570
rect 13789 274536 13801 274570
rect 12801 274524 13801 274536
rect 12801 274412 13801 274424
rect 12801 274378 12813 274412
rect 13789 274378 13801 274412
rect 12801 274366 13801 274378
rect 12801 274254 13801 274266
rect 12801 274220 12813 274254
rect 13789 274220 13801 274254
rect 12801 274208 13801 274220
rect 12801 274096 13801 274108
rect 12801 274062 12813 274096
rect 13789 274062 13801 274096
rect 12801 274050 13801 274062
rect 12801 273938 13801 273950
rect 12801 273904 12813 273938
rect 13789 273904 13801 273938
rect 12801 273892 13801 273904
rect 12801 273780 13801 273792
rect 12801 273746 12813 273780
rect 13789 273746 13801 273780
rect 12801 273734 13801 273746
rect 12801 273622 13801 273634
rect 12801 273588 12813 273622
rect 13789 273588 13801 273622
rect 12801 273576 13801 273588
rect 12801 273464 13801 273476
rect 12801 273430 12813 273464
rect 13789 273430 13801 273464
rect 12801 273418 13801 273430
rect 12801 273306 13801 273318
rect 12801 273272 12813 273306
rect 13789 273272 13801 273306
rect 12801 273260 13801 273272
rect 12801 273148 13801 273160
rect 12801 273114 12813 273148
rect 13789 273114 13801 273148
rect 12801 273102 13801 273114
rect 12801 272990 13801 273002
rect 12801 272956 12813 272990
rect 13789 272956 13801 272990
rect 12801 272944 13801 272956
rect 12801 272832 13801 272844
rect 12801 272798 12813 272832
rect 13789 272798 13801 272832
rect 12801 272786 13801 272798
rect 12801 272674 13801 272686
rect 12801 272640 12813 272674
rect 13789 272640 13801 272674
rect 12801 272628 13801 272640
rect 12801 272516 13801 272528
rect 12801 272482 12813 272516
rect 13789 272482 13801 272516
rect 12801 272470 13801 272482
rect 12801 272358 13801 272370
rect 12801 272324 12813 272358
rect 13789 272324 13801 272358
rect 12801 272312 13801 272324
rect 12801 272200 13801 272212
rect 12801 272166 12813 272200
rect 13789 272166 13801 272200
rect 12801 272154 13801 272166
rect 12801 272042 13801 272054
rect 12801 272008 12813 272042
rect 13789 272008 13801 272042
rect 12801 271996 13801 272008
rect 12801 271884 13801 271896
rect 12801 271850 12813 271884
rect 13789 271850 13801 271884
rect 12801 271838 13801 271850
rect 12801 271726 13801 271738
rect 12801 271692 12813 271726
rect 13789 271692 13801 271726
rect 12801 271680 13801 271692
rect 12801 271568 13801 271580
rect 12801 271534 12813 271568
rect 13789 271534 13801 271568
rect 12801 271522 13801 271534
rect 12801 271410 13801 271422
rect 12801 271376 12813 271410
rect 13789 271376 13801 271410
rect 12801 271364 13801 271376
rect 12801 271252 13801 271264
rect 12801 271218 12813 271252
rect 13789 271218 13801 271252
rect 12801 271206 13801 271218
rect 12801 271094 13801 271106
rect 12801 271060 12813 271094
rect 13789 271060 13801 271094
rect 12801 271048 13801 271060
rect 12801 270936 13801 270948
rect 12801 270902 12813 270936
rect 13789 270902 13801 270936
rect 12801 270890 13801 270902
rect 12801 270778 13801 270790
rect 12801 270744 12813 270778
rect 13789 270744 13801 270778
rect 12801 270732 13801 270744
rect 12801 270620 13801 270632
rect 12801 270586 12813 270620
rect 13789 270586 13801 270620
rect 12801 270574 13801 270586
rect 12801 270462 13801 270474
rect 12801 270428 12813 270462
rect 13789 270428 13801 270462
rect 12801 270416 13801 270428
rect 12801 270304 13801 270316
rect 12801 270270 12813 270304
rect 13789 270270 13801 270304
rect 12801 270258 13801 270270
rect 12801 270146 13801 270158
rect 12801 270112 12813 270146
rect 13789 270112 13801 270146
rect 12801 270100 13801 270112
rect 12801 269988 13801 270000
rect 12801 269954 12813 269988
rect 13789 269954 13801 269988
rect 12801 269942 13801 269954
rect 12801 269830 13801 269842
rect 12801 269796 12813 269830
rect 13789 269796 13801 269830
rect 12801 269784 13801 269796
rect 12801 269672 13801 269684
rect 12801 269638 12813 269672
rect 13789 269638 13801 269672
rect 12801 269626 13801 269638
rect 12801 269514 13801 269526
rect 12801 269480 12813 269514
rect 13789 269480 13801 269514
rect 12801 269468 13801 269480
rect 14471 274332 15471 274344
rect 14471 274298 14483 274332
rect 15459 274298 15471 274332
rect 14471 274286 15471 274298
rect 14471 274174 15471 274186
rect 14471 274140 14483 274174
rect 15459 274140 15471 274174
rect 14471 274128 15471 274140
rect 14471 274016 15471 274028
rect 14471 273982 14483 274016
rect 15459 273982 15471 274016
rect 14471 273970 15471 273982
rect 14471 273858 15471 273870
rect 14471 273824 14483 273858
rect 15459 273824 15471 273858
rect 14471 273812 15471 273824
rect 14471 273700 15471 273712
rect 14471 273666 14483 273700
rect 15459 273666 15471 273700
rect 14471 273654 15471 273666
rect 14471 273542 15471 273554
rect 14471 273508 14483 273542
rect 15459 273508 15471 273542
rect 14471 273496 15471 273508
rect 14471 273384 15471 273396
rect 14471 273350 14483 273384
rect 15459 273350 15471 273384
rect 14471 273338 15471 273350
rect 14471 273226 15471 273238
rect 14471 273192 14483 273226
rect 15459 273192 15471 273226
rect 14471 273180 15471 273192
rect 14471 273068 15471 273080
rect 14471 273034 14483 273068
rect 15459 273034 15471 273068
rect 14471 273022 15471 273034
rect 14471 272910 15471 272922
rect 14471 272876 14483 272910
rect 15459 272876 15471 272910
rect 14471 272864 15471 272876
rect 14471 272752 15471 272764
rect 14471 272718 14483 272752
rect 15459 272718 15471 272752
rect 14471 272706 15471 272718
rect 14471 272594 15471 272606
rect 14471 272560 14483 272594
rect 15459 272560 15471 272594
rect 14471 272548 15471 272560
rect 14471 272436 15471 272448
rect 14471 272402 14483 272436
rect 15459 272402 15471 272436
rect 14471 272390 15471 272402
rect 14471 272278 15471 272290
rect 14471 272244 14483 272278
rect 15459 272244 15471 272278
rect 14471 272232 15471 272244
rect 14471 272120 15471 272132
rect 14471 272086 14483 272120
rect 15459 272086 15471 272120
rect 14471 272074 15471 272086
rect 14471 271962 15471 271974
rect 14471 271928 14483 271962
rect 15459 271928 15471 271962
rect 14471 271916 15471 271928
rect 14471 271804 15471 271816
rect 14471 271770 14483 271804
rect 15459 271770 15471 271804
rect 14471 271758 15471 271770
rect 14471 271646 15471 271658
rect 14471 271612 14483 271646
rect 15459 271612 15471 271646
rect 14471 271600 15471 271612
rect 14471 271488 15471 271500
rect 14471 271454 14483 271488
rect 15459 271454 15471 271488
rect 14471 271442 15471 271454
rect 14471 271330 15471 271342
rect 14471 271296 14483 271330
rect 15459 271296 15471 271330
rect 14471 271284 15471 271296
rect 14471 271172 15471 271184
rect 14471 271138 14483 271172
rect 15459 271138 15471 271172
rect 14471 271126 15471 271138
rect 14471 271014 15471 271026
rect 14471 270980 14483 271014
rect 15459 270980 15471 271014
rect 14471 270968 15471 270980
rect 16011 274332 17011 274344
rect 16011 274298 16023 274332
rect 16999 274298 17011 274332
rect 16011 274286 17011 274298
rect 16011 274174 17011 274186
rect 16011 274140 16023 274174
rect 16999 274140 17011 274174
rect 16011 274128 17011 274140
rect 16011 274016 17011 274028
rect 16011 273982 16023 274016
rect 16999 273982 17011 274016
rect 16011 273970 17011 273982
rect 16011 273858 17011 273870
rect 16011 273824 16023 273858
rect 16999 273824 17011 273858
rect 16011 273812 17011 273824
rect 16011 273700 17011 273712
rect 16011 273666 16023 273700
rect 16999 273666 17011 273700
rect 16011 273654 17011 273666
rect 16011 273542 17011 273554
rect 16011 273508 16023 273542
rect 16999 273508 17011 273542
rect 16011 273496 17011 273508
rect 16011 273384 17011 273396
rect 16011 273350 16023 273384
rect 16999 273350 17011 273384
rect 16011 273338 17011 273350
rect 16011 273226 17011 273238
rect 16011 273192 16023 273226
rect 16999 273192 17011 273226
rect 16011 273180 17011 273192
rect 16011 273068 17011 273080
rect 16011 273034 16023 273068
rect 16999 273034 17011 273068
rect 16011 273022 17011 273034
rect 16011 272910 17011 272922
rect 16011 272876 16023 272910
rect 16999 272876 17011 272910
rect 16011 272864 17011 272876
rect 16011 272752 17011 272764
rect 16011 272718 16023 272752
rect 16999 272718 17011 272752
rect 16011 272706 17011 272718
rect 16011 272594 17011 272606
rect 16011 272560 16023 272594
rect 16999 272560 17011 272594
rect 16011 272548 17011 272560
rect 16011 272436 17011 272448
rect 16011 272402 16023 272436
rect 16999 272402 17011 272436
rect 16011 272390 17011 272402
rect 16011 272278 17011 272290
rect 16011 272244 16023 272278
rect 16999 272244 17011 272278
rect 16011 272232 17011 272244
rect 16011 272120 17011 272132
rect 16011 272086 16023 272120
rect 16999 272086 17011 272120
rect 16011 272074 17011 272086
rect 16011 271962 17011 271974
rect 16011 271928 16023 271962
rect 16999 271928 17011 271962
rect 16011 271916 17011 271928
rect 16011 271804 17011 271816
rect 16011 271770 16023 271804
rect 16999 271770 17011 271804
rect 16011 271758 17011 271770
rect 16011 271646 17011 271658
rect 16011 271612 16023 271646
rect 16999 271612 17011 271646
rect 16011 271600 17011 271612
rect 16011 271488 17011 271500
rect 16011 271454 16023 271488
rect 16999 271454 17011 271488
rect 16011 271442 17011 271454
rect 16011 271330 17011 271342
rect 16011 271296 16023 271330
rect 16999 271296 17011 271330
rect 16011 271284 17011 271296
rect 16011 271172 17011 271184
rect 16011 271138 16023 271172
rect 16999 271138 17011 271172
rect 16011 271126 17011 271138
rect 16011 271014 17011 271026
rect 16011 270980 16023 271014
rect 16999 270980 17011 271014
rect 16011 270968 17011 270980
rect 24181 273442 25181 273454
rect 24181 273408 24193 273442
rect 25169 273408 25181 273442
rect 24181 273396 25181 273408
rect 24181 273184 25181 273196
rect 24181 273150 24193 273184
rect 25169 273150 25181 273184
rect 24181 273138 25181 273150
rect 24181 272926 25181 272938
rect 24181 272892 24193 272926
rect 25169 272892 25181 272926
rect 24181 272880 25181 272892
rect 24181 272668 25181 272680
rect 24181 272634 24193 272668
rect 25169 272634 25181 272668
rect 24181 272622 25181 272634
rect 24181 272410 25181 272422
rect 24181 272376 24193 272410
rect 25169 272376 25181 272410
rect 24181 272364 25181 272376
rect 24181 272152 25181 272164
rect 24181 272118 24193 272152
rect 25169 272118 25181 272152
rect 24181 272106 25181 272118
rect 24181 271894 25181 271906
rect 24181 271860 24193 271894
rect 25169 271860 25181 271894
rect 24181 271848 25181 271860
rect 25681 273442 26681 273454
rect 25681 273408 25693 273442
rect 26669 273408 26681 273442
rect 25681 273396 26681 273408
rect 25681 273184 26681 273196
rect 25681 273150 25693 273184
rect 26669 273150 26681 273184
rect 25681 273138 26681 273150
rect 25681 272926 26681 272938
rect 25681 272892 25693 272926
rect 26669 272892 26681 272926
rect 25681 272880 26681 272892
rect 25681 272668 26681 272680
rect 25681 272634 25693 272668
rect 26669 272634 26681 272668
rect 25681 272622 26681 272634
rect 25681 272410 26681 272422
rect 25681 272376 25693 272410
rect 26669 272376 26681 272410
rect 25681 272364 26681 272376
rect 25681 272152 26681 272164
rect 25681 272118 25693 272152
rect 26669 272118 26681 272152
rect 25681 272106 26681 272118
rect 25681 271894 26681 271906
rect 25681 271860 25693 271894
rect 26669 271860 26681 271894
rect 25681 271848 26681 271860
<< ndiffc >>
rect 6002 304330 15978 304364
rect 6002 304232 15978 304266
rect 6002 304134 15978 304168
rect 6002 304036 15978 304070
rect 6002 303938 15978 303972
rect 6002 303840 15978 303874
rect 6002 303742 15978 303776
rect 6002 303644 15978 303678
rect 6002 303546 15978 303580
rect 6002 303448 15978 303482
rect 6002 303350 15978 303384
rect 559950 295822 559984 305798
rect 560048 295822 560082 305798
rect 560146 295822 560180 305798
rect 560244 295822 560278 305798
rect 560342 295822 560376 305798
rect 560440 295822 560474 305798
rect 560538 295822 560572 305798
rect 560636 295822 560670 305798
rect 560734 295822 560768 305798
rect 560832 295822 560866 305798
rect 560930 295822 560964 305798
rect 569150 295822 569184 305798
rect 569248 295822 569282 305798
rect 569346 295822 569380 305798
rect 569444 295822 569478 305798
rect 569542 295822 569576 305798
rect 569640 295822 569674 305798
rect 569738 295822 569772 305798
rect 569836 295822 569870 305798
rect 569934 295822 569968 305798
rect 570032 295822 570066 305798
rect 570130 295822 570164 305798
rect 6002 293930 15978 293964
rect 6002 293832 15978 293866
rect 6002 293734 15978 293768
rect 6002 293636 15978 293670
rect 6002 293538 15978 293572
rect 6002 293440 15978 293474
rect 6002 293342 15978 293376
rect 6002 293244 15978 293278
rect 6002 293146 15978 293180
rect 6002 293048 15978 293082
rect 6002 292950 15978 292984
rect 536471 289030 537447 289064
rect 537689 289030 538665 289064
rect 538907 289030 539883 289064
rect 540125 289030 541101 289064
rect 541343 289030 542319 289064
rect 542561 289030 543537 289064
rect 543779 289030 544755 289064
rect 536471 288872 537447 288906
rect 537689 288872 538665 288906
rect 538907 288872 539883 288906
rect 540125 288872 541101 288906
rect 541343 288872 542319 288906
rect 542561 288872 543537 288906
rect 543779 288872 544755 288906
rect 536471 288530 537447 288564
rect 537689 288530 538665 288564
rect 538907 288530 539883 288564
rect 540125 288530 541101 288564
rect 541343 288530 542319 288564
rect 542561 288530 543537 288564
rect 543779 288530 544755 288564
rect 536471 288372 537447 288406
rect 537689 288372 538665 288406
rect 538907 288372 539883 288406
rect 540125 288372 541101 288406
rect 541343 288372 542319 288406
rect 542561 288372 543537 288406
rect 543779 288372 544755 288406
rect 537031 288030 538007 288064
rect 538249 288030 539225 288064
rect 539467 288030 540443 288064
rect 540685 288030 541661 288064
rect 541903 288030 542879 288064
rect 543121 288030 544097 288064
rect 537031 287772 538007 287806
rect 538249 287772 539225 287806
rect 539467 287772 540443 287806
rect 540685 287772 541661 287806
rect 541903 287772 542879 287806
rect 543121 287772 544097 287806
rect 568302 288710 578278 288744
rect 568302 288612 578278 288646
rect 568302 288514 578278 288548
rect 568302 288416 578278 288450
rect 568302 288318 578278 288352
rect 568302 288220 578278 288254
rect 568302 288122 578278 288156
rect 568302 288024 578278 288058
rect 568302 287926 578278 287960
rect 568302 287828 578278 287862
rect 568302 287730 578278 287764
rect 537031 287410 538007 287444
rect 538249 287410 539225 287444
rect 539467 287410 540443 287444
rect 540685 287410 541661 287444
rect 541903 287410 542879 287444
rect 543121 287410 544097 287444
rect 537031 287152 538007 287186
rect 538249 287152 539225 287186
rect 539467 287152 540443 287186
rect 540685 287152 541661 287186
rect 541903 287152 542879 287186
rect 543121 287152 544097 287186
rect 536471 286810 537447 286844
rect 537689 286810 538665 286844
rect 538907 286810 539883 286844
rect 540125 286810 541101 286844
rect 541343 286810 542319 286844
rect 542561 286810 543537 286844
rect 543779 286810 544755 286844
rect 536471 286552 537447 286586
rect 537689 286552 538665 286586
rect 538907 286552 539883 286586
rect 540125 286552 541101 286586
rect 541343 286552 542319 286586
rect 542561 286552 543537 286586
rect 543779 286552 544755 286586
rect 536471 286210 537447 286244
rect 537689 286210 538665 286244
rect 538907 286210 539883 286244
rect 540125 286210 541101 286244
rect 541343 286210 542319 286244
rect 542561 286210 543537 286244
rect 543779 286210 544755 286244
rect 536471 285952 537447 285986
rect 537689 285952 538665 285986
rect 538907 285952 539883 285986
rect 540125 285952 541101 285986
rect 541343 285952 542319 285986
rect 542561 285952 543537 285986
rect 543779 285952 544755 285986
rect 539786 283856 540012 283890
rect 540254 283856 540480 283890
rect 540722 283856 540948 283890
rect 541190 283856 541416 283890
rect 539786 283598 540012 283632
rect 540254 283598 540480 283632
rect 540722 283598 540948 283632
rect 541190 283598 541416 283632
rect 540006 283231 540482 283265
rect 540724 283231 541200 283265
rect 540006 283073 540482 283107
rect 540724 283073 541200 283107
rect 537071 282706 538047 282740
rect 538289 282706 539265 282740
rect 539507 282706 540483 282740
rect 540725 282706 541701 282740
rect 541943 282706 542919 282740
rect 543161 282706 544137 282740
rect 537071 282448 538047 282482
rect 538289 282448 539265 282482
rect 539507 282448 540483 282482
rect 540725 282448 541701 282482
rect 541943 282448 542919 282482
rect 543161 282448 544137 282482
rect 568322 281230 578298 281264
rect 568322 281132 578298 281166
rect 568322 281034 578298 281068
rect 568322 280936 578298 280970
rect 568322 280838 578298 280872
rect 568322 280740 578298 280774
rect 568322 280642 578298 280676
rect 568322 280544 578298 280578
rect 568322 280446 578298 280480
rect 568322 280348 578298 280382
rect 568322 280250 578298 280284
rect 17591 273187 18567 273221
rect 17591 273029 18567 273063
rect 17591 272871 18567 272905
rect 17591 272713 18567 272747
rect 17591 272555 18567 272589
rect 17591 272397 18567 272431
rect 17591 272239 18567 272273
rect 17591 272081 18567 272115
rect 19111 273187 20087 273221
rect 19111 273029 20087 273063
rect 19111 272871 20087 272905
rect 19111 272713 20087 272747
rect 19111 272555 20087 272589
rect 19111 272397 20087 272431
rect 19111 272239 20087 272273
rect 19111 272081 20087 272115
rect 20632 274186 21608 274220
rect 20632 273928 21608 273962
rect 20632 273670 21608 273704
rect 20632 273412 21608 273446
rect 20632 273154 21608 273188
rect 20632 272896 21608 272930
rect 20632 272638 21608 272672
rect 20632 272380 21608 272414
rect 20632 272122 21608 272156
rect 20632 271864 21608 271898
rect 20632 271606 21608 271640
rect 20632 271348 21608 271382
rect 20632 271090 21608 271124
rect 22152 274442 23128 274476
rect 22152 274184 23128 274218
rect 22152 273926 23128 273960
rect 22152 273668 23128 273702
rect 22152 273410 23128 273444
rect 22152 273152 23128 273186
rect 22152 272894 23128 272928
rect 22152 272636 23128 272670
rect 22152 272378 23128 272412
rect 22152 272120 23128 272154
rect 22152 271862 23128 271896
rect 22152 271604 23128 271638
rect 22152 271346 23128 271380
rect 22152 271088 23128 271122
rect 22152 270830 23128 270864
rect 27302 272776 27778 272810
rect 27302 272618 27778 272652
rect 27302 272460 27778 272494
rect 28302 273132 28528 273166
rect 28302 272874 28528 272908
rect 28302 272616 28528 272650
rect 28302 272358 28528 272392
rect 28302 272100 28528 272134
rect 29052 273393 30028 273427
rect 29052 273135 30028 273169
rect 29052 272877 30028 272911
rect 29052 272619 30028 272653
rect 29052 272361 30028 272395
rect 29052 272103 30028 272137
rect 29052 271845 30028 271879
rect 6002 252330 15978 252364
rect 6002 252232 15978 252266
rect 6002 252134 15978 252168
rect 6002 252036 15978 252070
rect 6002 251938 15978 251972
rect 6002 251840 15978 251874
rect 6002 251742 15978 251776
rect 6002 251644 15978 251678
rect 6002 251546 15978 251580
rect 6002 251448 15978 251482
rect 6002 251350 15978 251384
rect 6002 241930 15978 241964
rect 6002 241832 15978 241866
rect 6002 241734 15978 241768
rect 6002 241636 15978 241670
rect 6002 241538 15978 241572
rect 6002 241440 15978 241474
rect 6002 241342 15978 241376
rect 6002 241244 15978 241278
rect 6002 241146 15978 241180
rect 6002 241048 15978 241082
rect 6002 240950 15978 240984
<< pdiffc >>
rect 536380 294750 537356 294784
rect 537616 294750 538592 294784
rect 538852 294750 539828 294784
rect 540088 294750 541064 294784
rect 541324 294750 542300 294784
rect 542560 294750 543536 294784
rect 543796 294750 544772 294784
rect 536380 294592 537356 294626
rect 537616 294592 538592 294626
rect 538852 294592 539828 294626
rect 540088 294592 541064 294626
rect 541324 294592 542300 294626
rect 542560 294592 543536 294626
rect 543796 294592 544772 294626
rect 536380 294210 537356 294244
rect 537616 294210 538592 294244
rect 538852 294210 539828 294244
rect 540088 294210 541064 294244
rect 541324 294210 542300 294244
rect 542560 294210 543536 294244
rect 543796 294210 544772 294244
rect 536380 294052 537356 294086
rect 537616 294052 538592 294086
rect 538852 294052 539828 294086
rect 540088 294052 541064 294086
rect 541324 294052 542300 294086
rect 542560 294052 543536 294086
rect 543796 294052 544772 294086
rect 536380 293670 537356 293704
rect 537616 293670 538592 293704
rect 538852 293670 539828 293704
rect 540088 293670 541064 293704
rect 541324 293670 542300 293704
rect 542560 293670 543536 293704
rect 543796 293670 544772 293704
rect 536380 293512 537356 293546
rect 537616 293512 538592 293546
rect 538852 293512 539828 293546
rect 540088 293512 541064 293546
rect 541324 293512 542300 293546
rect 542560 293512 543536 293546
rect 543796 293512 544772 293546
rect 536380 293130 537356 293164
rect 537616 293130 538592 293164
rect 538852 293130 539828 293164
rect 540088 293130 541064 293164
rect 541324 293130 542300 293164
rect 542560 293130 543536 293164
rect 543796 293130 544772 293164
rect 536380 292972 537356 293006
rect 537616 292972 538592 293006
rect 538852 292972 539828 293006
rect 540088 292972 541064 293006
rect 541324 292972 542300 293006
rect 542560 292972 543536 293006
rect 543796 292972 544772 293006
rect 536380 292550 537356 292584
rect 537616 292550 538592 292584
rect 538852 292550 539828 292584
rect 540088 292550 541064 292584
rect 541324 292550 542300 292584
rect 542560 292550 543536 292584
rect 543796 292550 544772 292584
rect 536380 292392 537356 292426
rect 537616 292392 538592 292426
rect 538852 292392 539828 292426
rect 540088 292392 541064 292426
rect 541324 292392 542300 292426
rect 542560 292392 543536 292426
rect 543796 292392 544772 292426
rect 536380 291970 537356 292004
rect 537616 291970 538592 292004
rect 538852 291970 539828 292004
rect 540088 291970 541064 292004
rect 541324 291970 542300 292004
rect 542560 291970 543536 292004
rect 543796 291970 544772 292004
rect 536380 291812 537356 291846
rect 537616 291812 538592 291846
rect 538852 291812 539828 291846
rect 540088 291812 541064 291846
rect 541324 291812 542300 291846
rect 542560 291812 543536 291846
rect 543796 291812 544772 291846
rect 534540 291430 535516 291464
rect 535776 291430 536752 291464
rect 537012 291430 537988 291464
rect 538248 291430 539224 291464
rect 539484 291430 540460 291464
rect 540720 291430 541696 291464
rect 541956 291430 542932 291464
rect 543192 291430 544168 291464
rect 544428 291430 545404 291464
rect 545664 291430 546640 291464
rect 534540 291272 535516 291306
rect 535776 291272 536752 291306
rect 537012 291272 537988 291306
rect 538248 291272 539224 291306
rect 539484 291272 540460 291306
rect 540720 291272 541696 291306
rect 541956 291272 542932 291306
rect 543192 291272 544168 291306
rect 544428 291272 545404 291306
rect 545664 291272 546640 291306
rect 534540 290890 535516 290924
rect 535776 290890 536752 290924
rect 537012 290890 537988 290924
rect 538248 290890 539224 290924
rect 539484 290890 540460 290924
rect 540720 290890 541696 290924
rect 541956 290890 542932 290924
rect 543192 290890 544168 290924
rect 544428 290890 545404 290924
rect 545664 290890 546640 290924
rect 534540 290732 535516 290766
rect 535776 290732 536752 290766
rect 537012 290732 537988 290766
rect 538248 290732 539224 290766
rect 539484 290732 540460 290766
rect 540720 290732 541696 290766
rect 541956 290732 542932 290766
rect 543192 290732 544168 290766
rect 544428 290732 545404 290766
rect 545664 290732 546640 290766
rect 534540 290350 535516 290384
rect 535776 290350 536752 290384
rect 537012 290350 537988 290384
rect 538248 290350 539224 290384
rect 539484 290350 540460 290384
rect 540720 290350 541696 290384
rect 541956 290350 542932 290384
rect 543192 290350 544168 290384
rect 544428 290350 545404 290384
rect 545664 290350 546640 290384
rect 534540 290192 535516 290226
rect 535776 290192 536752 290226
rect 537012 290192 537988 290226
rect 538248 290192 539224 290226
rect 539484 290192 540460 290226
rect 540720 290192 541696 290226
rect 541956 290192 542932 290226
rect 543192 290192 544168 290226
rect 544428 290192 545404 290226
rect 545664 290192 546640 290226
rect 534540 289810 535516 289844
rect 535776 289810 536752 289844
rect 537012 289810 537988 289844
rect 538248 289810 539224 289844
rect 539484 289810 540460 289844
rect 540720 289810 541696 289844
rect 541956 289810 542932 289844
rect 543192 289810 544168 289844
rect 544428 289810 545404 289844
rect 545664 289810 546640 289844
rect 534540 289652 535516 289686
rect 535776 289652 536752 289686
rect 537012 289652 537988 289686
rect 538248 289652 539224 289686
rect 539484 289652 540460 289686
rect 540720 289652 541696 289686
rect 541956 289652 542932 289686
rect 543192 289652 544168 289686
rect 544428 289652 545404 289686
rect 545664 289652 546640 289686
rect 537025 285236 538001 285270
rect 538261 285236 539237 285270
rect 539497 285236 540473 285270
rect 540733 285236 541709 285270
rect 541969 285236 542945 285270
rect 543205 285236 544181 285270
rect 537025 284978 538001 285012
rect 538261 284978 539237 285012
rect 539497 284978 540473 285012
rect 540733 284978 541709 285012
rect 541969 284978 542945 285012
rect 543205 284978 544181 285012
rect 537025 284646 538001 284680
rect 538261 284646 539237 284680
rect 539497 284646 540473 284680
rect 540733 284646 541709 284680
rect 541969 284646 542945 284680
rect 543205 284646 544181 284680
rect 537025 284388 538001 284422
rect 538261 284388 539237 284422
rect 539497 284388 540473 284422
rect 540733 284388 541709 284422
rect 541969 284388 542945 284422
rect 543205 284388 544181 284422
rect 12813 275800 13789 275834
rect 12813 275642 13789 275676
rect 12813 275484 13789 275518
rect 12813 275326 13789 275360
rect 12813 275168 13789 275202
rect 12813 275010 13789 275044
rect 12813 274852 13789 274886
rect 12813 274694 13789 274728
rect 12813 274536 13789 274570
rect 12813 274378 13789 274412
rect 12813 274220 13789 274254
rect 12813 274062 13789 274096
rect 12813 273904 13789 273938
rect 12813 273746 13789 273780
rect 12813 273588 13789 273622
rect 12813 273430 13789 273464
rect 12813 273272 13789 273306
rect 12813 273114 13789 273148
rect 12813 272956 13789 272990
rect 12813 272798 13789 272832
rect 12813 272640 13789 272674
rect 12813 272482 13789 272516
rect 12813 272324 13789 272358
rect 12813 272166 13789 272200
rect 12813 272008 13789 272042
rect 12813 271850 13789 271884
rect 12813 271692 13789 271726
rect 12813 271534 13789 271568
rect 12813 271376 13789 271410
rect 12813 271218 13789 271252
rect 12813 271060 13789 271094
rect 12813 270902 13789 270936
rect 12813 270744 13789 270778
rect 12813 270586 13789 270620
rect 12813 270428 13789 270462
rect 12813 270270 13789 270304
rect 12813 270112 13789 270146
rect 12813 269954 13789 269988
rect 12813 269796 13789 269830
rect 12813 269638 13789 269672
rect 12813 269480 13789 269514
rect 14483 274298 15459 274332
rect 14483 274140 15459 274174
rect 14483 273982 15459 274016
rect 14483 273824 15459 273858
rect 14483 273666 15459 273700
rect 14483 273508 15459 273542
rect 14483 273350 15459 273384
rect 14483 273192 15459 273226
rect 14483 273034 15459 273068
rect 14483 272876 15459 272910
rect 14483 272718 15459 272752
rect 14483 272560 15459 272594
rect 14483 272402 15459 272436
rect 14483 272244 15459 272278
rect 14483 272086 15459 272120
rect 14483 271928 15459 271962
rect 14483 271770 15459 271804
rect 14483 271612 15459 271646
rect 14483 271454 15459 271488
rect 14483 271296 15459 271330
rect 14483 271138 15459 271172
rect 14483 270980 15459 271014
rect 16023 274298 16999 274332
rect 16023 274140 16999 274174
rect 16023 273982 16999 274016
rect 16023 273824 16999 273858
rect 16023 273666 16999 273700
rect 16023 273508 16999 273542
rect 16023 273350 16999 273384
rect 16023 273192 16999 273226
rect 16023 273034 16999 273068
rect 16023 272876 16999 272910
rect 16023 272718 16999 272752
rect 16023 272560 16999 272594
rect 16023 272402 16999 272436
rect 16023 272244 16999 272278
rect 16023 272086 16999 272120
rect 16023 271928 16999 271962
rect 16023 271770 16999 271804
rect 16023 271612 16999 271646
rect 16023 271454 16999 271488
rect 16023 271296 16999 271330
rect 16023 271138 16999 271172
rect 16023 270980 16999 271014
rect 24193 273408 25169 273442
rect 24193 273150 25169 273184
rect 24193 272892 25169 272926
rect 24193 272634 25169 272668
rect 24193 272376 25169 272410
rect 24193 272118 25169 272152
rect 24193 271860 25169 271894
rect 25693 273408 26669 273442
rect 25693 273150 26669 273184
rect 25693 272892 26669 272926
rect 25693 272634 26669 272668
rect 25693 272376 26669 272410
rect 25693 272118 26669 272152
rect 25693 271860 26669 271894
<< psubdiff >>
rect 559836 305950 561078 305984
rect 559836 305888 559870 305950
rect 5816 304444 5912 304478
rect 16068 304444 16164 304478
rect 5816 303270 5850 304444
rect 16130 304382 16164 304444
rect 16130 303270 16164 303332
rect 5816 303236 5912 303270
rect 16068 303236 16164 303270
rect 561044 305888 561078 305950
rect 559836 295670 559870 295732
rect 561044 295670 561078 295732
rect 559836 295636 559932 295670
rect 560982 295636 561078 295670
rect 569036 305950 570278 305984
rect 569036 305888 569070 305950
rect 570244 305888 570278 305950
rect 569036 295670 569070 295732
rect 570244 295670 570278 295732
rect 569036 295636 569132 295670
rect 570182 295636 570278 295670
rect 5816 294044 5912 294078
rect 16068 294044 16164 294078
rect 5816 292870 5850 294044
rect 16130 293982 16164 294044
rect 16130 292870 16164 292932
rect 5816 292836 5912 292870
rect 16068 292836 16164 292870
rect 530592 292067 530688 292101
rect 533620 292067 533716 292101
rect 530592 292005 530626 292067
rect 533682 292005 533716 292067
rect 530592 290729 530626 290791
rect 547652 292067 547748 292101
rect 550680 292067 550776 292101
rect 547652 292005 547686 292067
rect 533682 290729 533716 290791
rect 530592 290695 530688 290729
rect 533620 290695 533716 290729
rect 550742 292005 550776 292067
rect 547652 290729 547686 290791
rect 550742 290729 550776 290791
rect 547652 290695 547748 290729
rect 550680 290695 550776 290729
rect 530592 290597 530688 290631
rect 533620 290597 533716 290631
rect 530592 290535 530626 290597
rect 533682 290535 533716 290597
rect 530592 289259 530626 289321
rect 547652 290597 547748 290631
rect 550680 290597 550776 290631
rect 547652 290535 547686 290597
rect 533682 289259 533716 289321
rect 530592 289225 530688 289259
rect 533620 289225 533716 289259
rect 550742 290535 550776 290597
rect 547652 289259 547686 289321
rect 550742 289259 550776 289321
rect 547652 289225 547748 289259
rect 550680 289225 550776 289259
rect 536285 289144 536381 289178
rect 544845 289144 544941 289178
rect 536285 289082 536319 289144
rect 544907 289082 544941 289144
rect 536285 288792 536319 288854
rect 544907 288792 544941 288854
rect 536285 288758 536381 288792
rect 544845 288758 544941 288792
rect 568116 288824 568212 288858
rect 578368 288824 578464 288858
rect 568116 288762 568150 288824
rect 536285 288644 536381 288678
rect 544845 288644 544941 288678
rect 536285 288582 536319 288644
rect 544907 288582 544941 288644
rect 536285 288292 536319 288354
rect 544907 288292 544941 288354
rect 536285 288258 536381 288292
rect 544845 288258 544941 288292
rect 536845 288144 536941 288178
rect 544187 288144 544283 288178
rect 536845 288082 536879 288144
rect 544249 288082 544283 288144
rect 536845 287692 536879 287754
rect 544249 287692 544283 287754
rect 536845 287658 536941 287692
rect 544187 287658 544283 287692
rect 568116 287650 568150 287712
rect 578430 287650 578464 288824
rect 568116 287616 568212 287650
rect 578368 287616 578464 287650
rect 536845 287524 536941 287558
rect 544187 287524 544283 287558
rect 536845 287462 536879 287524
rect 544249 287462 544283 287524
rect 536845 287072 536879 287134
rect 544249 287072 544283 287134
rect 536845 287038 536941 287072
rect 544187 287038 544283 287072
rect 536285 286924 536381 286958
rect 544845 286924 544941 286958
rect 536285 286862 536319 286924
rect 544907 286862 544941 286924
rect 536285 286472 536319 286534
rect 544907 286472 544941 286534
rect 536285 286438 536381 286472
rect 544845 286438 544941 286472
rect 536285 286324 536381 286358
rect 544845 286324 544941 286358
rect 536285 286262 536319 286324
rect 544907 286262 544941 286324
rect 536285 285872 536319 285934
rect 544907 285872 544941 285934
rect 536285 285838 536381 285872
rect 544845 285838 544941 285872
rect 539600 283970 539696 284004
rect 541506 283970 541602 284004
rect 539600 283908 539634 283970
rect 541568 283908 541602 283970
rect 539600 283518 539634 283580
rect 541568 283518 541602 283580
rect 539600 283484 539696 283518
rect 541506 283484 541602 283518
rect 539820 283345 539916 283379
rect 541290 283345 541386 283379
rect 539820 283283 539854 283345
rect 541352 283283 541386 283345
rect 539820 282993 539854 283055
rect 541352 282993 541386 283055
rect 539820 282959 539916 282993
rect 541290 282959 541386 282993
rect 536885 282820 536981 282854
rect 544227 282820 544323 282854
rect 536885 282758 536919 282820
rect 544289 282758 544323 282820
rect 536885 282368 536919 282430
rect 544289 282368 544323 282430
rect 536885 282334 536981 282368
rect 544227 282334 544323 282368
rect 568136 281344 568232 281378
rect 578388 281344 578484 281378
rect 568136 281282 568170 281344
rect 537364 281058 537484 281082
rect 537364 280914 537484 280938
rect 543734 281058 543854 281082
rect 543734 280914 543854 280938
rect 568136 280170 568170 280232
rect 578450 280170 578484 281344
rect 568136 280136 568232 280170
rect 578388 280136 578484 280170
rect 11741 279723 11837 279757
rect 13051 279723 13147 279757
rect 11741 279661 11775 279723
rect 13113 279661 13147 279723
rect 11741 276667 11775 276729
rect 13113 276667 13147 276729
rect 11741 276633 11837 276667
rect 13051 276633 13147 276667
rect 13201 279723 13297 279757
rect 14511 279723 14607 279757
rect 13201 279661 13235 279723
rect 14573 279661 14607 279723
rect 13201 276667 13235 276729
rect 537364 278058 537484 278082
rect 537364 277914 537484 277938
rect 543734 278058 543854 278082
rect 543734 277914 543854 277938
rect 14573 276667 14607 276729
rect 13201 276633 13297 276667
rect 14511 276633 14607 276667
rect 30996 275900 31020 276140
rect 31260 275900 31284 276140
rect 32716 275900 32740 276140
rect 32980 275900 33004 276140
rect 34436 275900 34460 276140
rect 34700 275900 34724 276140
rect 35916 275900 35940 276140
rect 36180 275900 36204 276140
rect 37636 275900 37660 276140
rect 37900 275900 37924 276140
rect 39236 275900 39260 276140
rect 39500 275900 39524 276140
rect 40956 275900 40980 276140
rect 41220 275900 41244 276140
rect 42556 275900 42580 276140
rect 42820 275900 42844 276140
rect 44276 275900 44300 276140
rect 44540 275900 44564 276140
rect 537364 275058 537484 275082
rect 537364 274914 537484 274938
rect 543734 275058 543854 275082
rect 543734 274914 543854 274938
rect 21966 274556 22062 274590
rect 23218 274556 23314 274590
rect 21966 274494 22000 274556
rect 20446 274300 20542 274334
rect 21698 274300 21794 274334
rect 20446 274238 20480 274300
rect 17405 273301 17501 273335
rect 18657 273301 18753 273335
rect 17405 273239 17439 273301
rect 18719 273239 18753 273301
rect 17405 272001 17439 272063
rect 18719 272001 18753 272063
rect 17405 271967 17501 272001
rect 18657 271967 18753 272001
rect 18925 273301 19021 273335
rect 20177 273301 20273 273335
rect 18925 273239 18959 273301
rect 20239 273239 20273 273301
rect 18925 272001 18959 272063
rect 20239 272001 20273 272063
rect 18925 271967 19021 272001
rect 20177 271967 20273 272001
rect 21760 274238 21794 274300
rect 20446 271010 20480 271072
rect 21760 271010 21794 271072
rect 20446 270976 20542 271010
rect 21698 270976 21794 271010
rect 23280 274494 23314 274556
rect 21966 270750 22000 270812
rect 28866 273507 28962 273541
rect 30118 273507 30214 273541
rect 28866 273445 28900 273507
rect 28116 273246 28212 273280
rect 28618 273246 28714 273280
rect 28116 273184 28150 273246
rect 27116 272890 27212 272924
rect 27868 272890 27964 272924
rect 27116 272828 27150 272890
rect 27930 272828 27964 272890
rect 27116 272380 27150 272442
rect 27930 272380 27964 272442
rect 27116 272346 27212 272380
rect 27868 272346 27964 272380
rect 28680 273184 28714 273246
rect 28116 272020 28150 272082
rect 28680 272020 28714 272082
rect 28116 271986 28212 272020
rect 28618 271986 28714 272020
rect 30180 273445 30214 273507
rect 28866 271765 28900 271827
rect 537364 272058 537484 272082
rect 537364 271914 537484 271938
rect 543734 272058 543854 272082
rect 543734 271914 543854 271938
rect 30180 271765 30214 271827
rect 28866 271731 28962 271765
rect 30118 271731 30214 271765
rect 23280 270750 23314 270812
rect 21966 270716 22062 270750
rect 23218 270716 23314 270750
rect 30996 269200 31020 269440
rect 31260 269200 31284 269440
rect 32716 269200 32740 269440
rect 32980 269200 33004 269440
rect 34436 269200 34460 269440
rect 34700 269200 34724 269440
rect 35916 269200 35940 269440
rect 36180 269200 36204 269440
rect 37636 269200 37660 269440
rect 37900 269200 37924 269440
rect 39236 269200 39260 269440
rect 39500 269200 39524 269440
rect 40956 269200 40980 269440
rect 41220 269200 41244 269440
rect 42556 269200 42580 269440
rect 42820 269200 42844 269440
rect 44276 269200 44300 269440
rect 44540 269200 44564 269440
rect 537364 269058 537484 269082
rect 537364 268914 537484 268938
rect 543734 269058 543854 269082
rect 543734 268914 543854 268938
rect 11741 268653 11837 268687
rect 13051 268653 13147 268687
rect 11741 268591 11775 268653
rect 13113 268591 13147 268653
rect 11741 265597 11775 265659
rect 13113 265597 13147 265659
rect 11741 265563 11837 265597
rect 13051 265563 13147 265597
rect 13201 268653 13297 268687
rect 14511 268653 14607 268687
rect 13201 268591 13235 268653
rect 14573 268591 14607 268653
rect 13201 265597 13235 265659
rect 14573 265597 14607 265659
rect 13201 265563 13297 265597
rect 14511 265563 14607 265597
rect 5816 252444 5912 252478
rect 16068 252444 16164 252478
rect 5816 251270 5850 252444
rect 16130 252382 16164 252444
rect 16130 251270 16164 251332
rect 5816 251236 5912 251270
rect 16068 251236 16164 251270
rect 5816 242044 5912 242078
rect 16068 242044 16164 242078
rect 5816 240870 5850 242044
rect 16130 241982 16164 242044
rect 16130 240870 16164 240932
rect 5816 240836 5912 240870
rect 16068 240836 16164 240870
<< nsubdiff >>
rect 536185 294864 536281 294898
rect 544871 294864 544967 294898
rect 536185 294802 536219 294864
rect 544933 294802 544967 294864
rect 536185 294512 536219 294574
rect 544933 294512 544967 294574
rect 536185 294478 536281 294512
rect 544871 294478 544967 294512
rect 536185 294324 536281 294358
rect 544871 294324 544967 294358
rect 536185 294262 536219 294324
rect 544933 294262 544967 294324
rect 536185 293972 536219 294034
rect 544933 293972 544967 294034
rect 536185 293938 536281 293972
rect 544871 293938 544967 293972
rect 536185 293784 536281 293818
rect 544871 293784 544967 293818
rect 536185 293722 536219 293784
rect 544933 293722 544967 293784
rect 536185 293432 536219 293494
rect 544933 293432 544967 293494
rect 536185 293398 536281 293432
rect 544871 293398 544967 293432
rect 536185 293244 536281 293278
rect 544871 293244 544967 293278
rect 536185 293182 536219 293244
rect 544933 293182 544967 293244
rect 536185 292892 536219 292954
rect 544933 292892 544967 292954
rect 536185 292858 536281 292892
rect 544871 292858 544967 292892
rect 536185 292664 536281 292698
rect 544871 292664 544967 292698
rect 536185 292602 536219 292664
rect 544933 292602 544967 292664
rect 536185 292312 536219 292374
rect 544933 292312 544967 292374
rect 536185 292278 536281 292312
rect 544871 292278 544967 292312
rect 536185 292084 536281 292118
rect 544871 292084 544967 292118
rect 536185 292022 536219 292084
rect 544933 292022 544967 292084
rect 536185 291732 536219 291794
rect 544933 291732 544967 291794
rect 536185 291698 536281 291732
rect 544871 291698 544967 291732
rect 534345 291544 534441 291578
rect 546739 291544 546835 291578
rect 534345 291482 534379 291544
rect 546801 291482 546835 291544
rect 534345 291192 534379 291254
rect 546801 291192 546835 291254
rect 534345 291158 534441 291192
rect 546739 291158 546835 291192
rect 534345 291004 534441 291038
rect 546739 291004 546835 291038
rect 534345 290942 534379 291004
rect 546801 290942 546835 291004
rect 534345 290652 534379 290714
rect 546801 290652 546835 290714
rect 534345 290618 534441 290652
rect 546739 290618 546835 290652
rect 534345 290464 534441 290498
rect 546739 290464 546835 290498
rect 534345 290402 534379 290464
rect 546801 290402 546835 290464
rect 534345 290112 534379 290174
rect 546801 290112 546835 290174
rect 534345 290078 534441 290112
rect 546739 290078 546835 290112
rect 534345 289924 534441 289958
rect 546739 289924 546835 289958
rect 534345 289862 534379 289924
rect 546801 289862 546835 289924
rect 534345 289572 534379 289634
rect 546801 289572 546835 289634
rect 534345 289538 534441 289572
rect 546739 289538 546835 289572
rect 536830 285350 536926 285384
rect 544280 285350 544376 285384
rect 536830 285288 536864 285350
rect 544342 285288 544376 285350
rect 536830 284898 536864 284960
rect 544342 284898 544376 284960
rect 536830 284864 536926 284898
rect 544280 284864 544376 284898
rect 536830 284760 536926 284794
rect 544280 284760 544376 284794
rect 536830 284698 536864 284760
rect 544342 284698 544376 284760
rect 536830 284308 536864 284370
rect 544342 284308 544376 284370
rect 536830 284274 536926 284308
rect 544280 284274 544376 284308
rect 12618 275914 12714 275948
rect 13888 275914 13984 275948
rect 12618 275852 12652 275914
rect 13950 275852 13984 275914
rect 12618 269400 12652 269462
rect 14288 274412 14384 274446
rect 15558 274412 15654 274446
rect 14288 274350 14322 274412
rect 15620 274350 15654 274412
rect 14288 270900 14322 270962
rect 15620 270900 15654 270962
rect 14288 270866 14384 270900
rect 15558 270866 15654 270900
rect 15828 274412 15924 274446
rect 17098 274412 17194 274446
rect 15828 274350 15862 274412
rect 17160 274350 17194 274412
rect 15828 270900 15862 270962
rect 17160 270900 17194 270962
rect 15828 270866 15924 270900
rect 17098 270866 17194 270900
rect 23998 273522 24094 273556
rect 25268 273522 25364 273556
rect 23998 273460 24032 273522
rect 25330 273460 25364 273522
rect 23998 271780 24032 271842
rect 25330 271780 25364 271842
rect 23998 271746 24094 271780
rect 25268 271746 25364 271780
rect 25498 273522 25594 273556
rect 26768 273522 26864 273556
rect 25498 273460 25532 273522
rect 26830 273460 26864 273522
rect 25498 271780 25532 271842
rect 26830 271780 26864 271842
rect 25498 271746 25594 271780
rect 26768 271746 26864 271780
rect 13950 269400 13984 269462
rect 12618 269366 12714 269400
rect 13888 269366 13984 269400
<< psubdiffcont >>
rect 5912 304444 16068 304478
rect 16130 303332 16164 304382
rect 5912 303236 16068 303270
rect 559836 295732 559870 305888
rect 561044 295732 561078 305888
rect 559932 295636 560982 295670
rect 569036 295732 569070 305888
rect 570244 295732 570278 305888
rect 569132 295636 570182 295670
rect 5912 294044 16068 294078
rect 16130 292932 16164 293982
rect 5912 292836 16068 292870
rect 530688 292067 533620 292101
rect 530592 290791 530626 292005
rect 533682 290791 533716 292005
rect 547748 292067 550680 292101
rect 530688 290695 533620 290729
rect 547652 290791 547686 292005
rect 550742 290791 550776 292005
rect 547748 290695 550680 290729
rect 530688 290597 533620 290631
rect 530592 289321 530626 290535
rect 533682 289321 533716 290535
rect 547748 290597 550680 290631
rect 530688 289225 533620 289259
rect 547652 289321 547686 290535
rect 550742 289321 550776 290535
rect 547748 289225 550680 289259
rect 536381 289144 544845 289178
rect 536285 288854 536319 289082
rect 544907 288854 544941 289082
rect 536381 288758 544845 288792
rect 568212 288824 578368 288858
rect 536381 288644 544845 288678
rect 536285 288354 536319 288582
rect 544907 288354 544941 288582
rect 536381 288258 544845 288292
rect 536941 288144 544187 288178
rect 536845 287754 536879 288082
rect 544249 287754 544283 288082
rect 536941 287658 544187 287692
rect 568116 287712 568150 288762
rect 568212 287616 578368 287650
rect 536941 287524 544187 287558
rect 536845 287134 536879 287462
rect 544249 287134 544283 287462
rect 536941 287038 544187 287072
rect 536381 286924 544845 286958
rect 536285 286534 536319 286862
rect 544907 286534 544941 286862
rect 536381 286438 544845 286472
rect 536381 286324 544845 286358
rect 536285 285934 536319 286262
rect 544907 285934 544941 286262
rect 536381 285838 544845 285872
rect 539696 283970 541506 284004
rect 539600 283580 539634 283908
rect 541568 283580 541602 283908
rect 539696 283484 541506 283518
rect 539916 283345 541290 283379
rect 539820 283055 539854 283283
rect 541352 283055 541386 283283
rect 539916 282959 541290 282993
rect 536981 282820 544227 282854
rect 536885 282430 536919 282758
rect 544289 282430 544323 282758
rect 536981 282334 544227 282368
rect 568232 281344 578388 281378
rect 537364 280938 537484 281058
rect 543734 280938 543854 281058
rect 568136 280232 568170 281282
rect 568232 280136 578388 280170
rect 11837 279723 13051 279757
rect 11741 276729 11775 279661
rect 13113 276729 13147 279661
rect 11837 276633 13051 276667
rect 13297 279723 14511 279757
rect 13201 276729 13235 279661
rect 14573 276729 14607 279661
rect 537364 277938 537484 278058
rect 543734 277938 543854 278058
rect 13297 276633 14511 276667
rect 31020 275900 31260 276140
rect 32740 275900 32980 276140
rect 34460 275900 34700 276140
rect 35940 275900 36180 276140
rect 37660 275900 37900 276140
rect 39260 275900 39500 276140
rect 40980 275900 41220 276140
rect 42580 275900 42820 276140
rect 44300 275900 44540 276140
rect 537364 274938 537484 275058
rect 543734 274938 543854 275058
rect 22062 274556 23218 274590
rect 20542 274300 21698 274334
rect 17501 273301 18657 273335
rect 17405 272063 17439 273239
rect 18719 272063 18753 273239
rect 17501 271967 18657 272001
rect 19021 273301 20177 273335
rect 18925 272063 18959 273239
rect 20239 272063 20273 273239
rect 19021 271967 20177 272001
rect 20446 271072 20480 274238
rect 21760 271072 21794 274238
rect 20542 270976 21698 271010
rect 21966 270812 22000 274494
rect 23280 270812 23314 274494
rect 28962 273507 30118 273541
rect 28212 273246 28618 273280
rect 27212 272890 27868 272924
rect 27116 272442 27150 272828
rect 27930 272442 27964 272828
rect 27212 272346 27868 272380
rect 28116 272082 28150 273184
rect 28680 272082 28714 273184
rect 28212 271986 28618 272020
rect 28866 271827 28900 273445
rect 30180 271827 30214 273445
rect 537364 271938 537484 272058
rect 543734 271938 543854 272058
rect 28962 271731 30118 271765
rect 22062 270716 23218 270750
rect 31020 269200 31260 269440
rect 32740 269200 32980 269440
rect 34460 269200 34700 269440
rect 35940 269200 36180 269440
rect 37660 269200 37900 269440
rect 39260 269200 39500 269440
rect 40980 269200 41220 269440
rect 42580 269200 42820 269440
rect 44300 269200 44540 269440
rect 537364 268938 537484 269058
rect 543734 268938 543854 269058
rect 11837 268653 13051 268687
rect 11741 265659 11775 268591
rect 13113 265659 13147 268591
rect 11837 265563 13051 265597
rect 13297 268653 14511 268687
rect 13201 265659 13235 268591
rect 14573 265659 14607 268591
rect 13297 265563 14511 265597
rect 5912 252444 16068 252478
rect 16130 251332 16164 252382
rect 5912 251236 16068 251270
rect 5912 242044 16068 242078
rect 16130 240932 16164 241982
rect 5912 240836 16068 240870
<< nsubdiffcont >>
rect 536281 294864 544871 294898
rect 536185 294574 536219 294802
rect 544933 294574 544967 294802
rect 536281 294478 544871 294512
rect 536281 294324 544871 294358
rect 536185 294034 536219 294262
rect 544933 294034 544967 294262
rect 536281 293938 544871 293972
rect 536281 293784 544871 293818
rect 536185 293494 536219 293722
rect 544933 293494 544967 293722
rect 536281 293398 544871 293432
rect 536281 293244 544871 293278
rect 536185 292954 536219 293182
rect 544933 292954 544967 293182
rect 536281 292858 544871 292892
rect 536281 292664 544871 292698
rect 536185 292374 536219 292602
rect 544933 292374 544967 292602
rect 536281 292278 544871 292312
rect 536281 292084 544871 292118
rect 536185 291794 536219 292022
rect 544933 291794 544967 292022
rect 536281 291698 544871 291732
rect 534441 291544 546739 291578
rect 534345 291254 534379 291482
rect 546801 291254 546835 291482
rect 534441 291158 546739 291192
rect 534441 291004 546739 291038
rect 534345 290714 534379 290942
rect 546801 290714 546835 290942
rect 534441 290618 546739 290652
rect 534441 290464 546739 290498
rect 534345 290174 534379 290402
rect 546801 290174 546835 290402
rect 534441 290078 546739 290112
rect 534441 289924 546739 289958
rect 534345 289634 534379 289862
rect 546801 289634 546835 289862
rect 534441 289538 546739 289572
rect 536926 285350 544280 285384
rect 536830 284960 536864 285288
rect 544342 284960 544376 285288
rect 536926 284864 544280 284898
rect 536926 284760 544280 284794
rect 536830 284370 536864 284698
rect 544342 284370 544376 284698
rect 536926 284274 544280 284308
rect 12714 275914 13888 275948
rect 12618 269462 12652 275852
rect 13950 269462 13984 275852
rect 14384 274412 15558 274446
rect 14288 270962 14322 274350
rect 15620 270962 15654 274350
rect 14384 270866 15558 270900
rect 15924 274412 17098 274446
rect 15828 270962 15862 274350
rect 17160 270962 17194 274350
rect 15924 270866 17098 270900
rect 24094 273522 25268 273556
rect 23998 271842 24032 273460
rect 25330 271842 25364 273460
rect 24094 271746 25268 271780
rect 25594 273522 26768 273556
rect 25498 271842 25532 273460
rect 26830 271842 26864 273460
rect 25594 271746 26768 271780
rect 12714 269366 13888 269400
<< poly >>
rect 5902 304318 5968 304331
rect 5902 304315 5990 304318
rect 5902 304281 5918 304315
rect 5952 304281 5990 304315
rect 5902 304278 5990 304281
rect 15990 304278 16016 304318
rect 5902 304265 5968 304278
rect 16012 304220 16078 304233
rect 5964 304180 5990 304220
rect 15990 304217 16078 304220
rect 15990 304183 16028 304217
rect 16062 304183 16078 304217
rect 15990 304180 16078 304183
rect 5902 304122 5968 304135
rect 16012 304167 16078 304180
rect 5902 304119 5990 304122
rect 5902 304085 5918 304119
rect 5952 304085 5990 304119
rect 5902 304082 5990 304085
rect 15990 304082 16016 304122
rect 5902 304069 5968 304082
rect 16012 304024 16078 304037
rect 5964 303984 5990 304024
rect 15990 304021 16078 304024
rect 15990 303987 16028 304021
rect 16062 303987 16078 304021
rect 15990 303984 16078 303987
rect 5902 303926 5968 303939
rect 16012 303971 16078 303984
rect 5902 303923 5990 303926
rect 5902 303889 5918 303923
rect 5952 303889 5990 303923
rect 5902 303886 5990 303889
rect 15990 303886 16016 303926
rect 5902 303873 5968 303886
rect 16012 303828 16078 303841
rect 5964 303788 5990 303828
rect 15990 303825 16078 303828
rect 15990 303791 16028 303825
rect 16062 303791 16078 303825
rect 15990 303788 16078 303791
rect 5902 303730 5968 303743
rect 16012 303775 16078 303788
rect 5902 303727 5990 303730
rect 5902 303693 5918 303727
rect 5952 303693 5990 303727
rect 5902 303690 5990 303693
rect 15990 303690 16016 303730
rect 5902 303677 5968 303690
rect 16012 303632 16078 303645
rect 5964 303592 5990 303632
rect 15990 303629 16078 303632
rect 15990 303595 16028 303629
rect 16062 303595 16078 303629
rect 15990 303592 16078 303595
rect 5902 303534 5968 303547
rect 16012 303579 16078 303592
rect 5902 303531 5990 303534
rect 5902 303497 5918 303531
rect 5952 303497 5990 303531
rect 5902 303494 5990 303497
rect 15990 303494 16016 303534
rect 5902 303481 5968 303494
rect 16012 303436 16078 303449
rect 5964 303396 5990 303436
rect 15990 303433 16078 303436
rect 15990 303399 16028 303433
rect 16062 303399 16078 303433
rect 15990 303396 16078 303399
rect 16012 303383 16078 303396
rect 560081 305882 560147 305898
rect 560081 305848 560097 305882
rect 560131 305848 560147 305882
rect 559996 305810 560036 305836
rect 560081 305832 560147 305848
rect 560277 305882 560343 305898
rect 560277 305848 560293 305882
rect 560327 305848 560343 305882
rect 560094 305810 560134 305832
rect 560192 305810 560232 305836
rect 560277 305832 560343 305848
rect 560473 305882 560539 305898
rect 560473 305848 560489 305882
rect 560523 305848 560539 305882
rect 560290 305810 560330 305832
rect 560388 305810 560428 305836
rect 560473 305832 560539 305848
rect 560669 305882 560735 305898
rect 560669 305848 560685 305882
rect 560719 305848 560735 305882
rect 560486 305810 560526 305832
rect 560584 305810 560624 305836
rect 560669 305832 560735 305848
rect 560865 305882 560931 305898
rect 560865 305848 560881 305882
rect 560915 305848 560931 305882
rect 560682 305810 560722 305832
rect 560780 305810 560820 305836
rect 560865 305832 560931 305848
rect 560878 305810 560918 305832
rect 559996 295788 560036 295810
rect 559983 295772 560049 295788
rect 560094 295784 560134 295810
rect 560192 295788 560232 295810
rect 559983 295738 559999 295772
rect 560033 295738 560049 295772
rect 559983 295722 560049 295738
rect 560179 295772 560245 295788
rect 560290 295784 560330 295810
rect 560388 295788 560428 295810
rect 560179 295738 560195 295772
rect 560229 295738 560245 295772
rect 560179 295722 560245 295738
rect 560375 295772 560441 295788
rect 560486 295784 560526 295810
rect 560584 295788 560624 295810
rect 560375 295738 560391 295772
rect 560425 295738 560441 295772
rect 560375 295722 560441 295738
rect 560571 295772 560637 295788
rect 560682 295784 560722 295810
rect 560780 295788 560820 295810
rect 560571 295738 560587 295772
rect 560621 295738 560637 295772
rect 560571 295722 560637 295738
rect 560767 295772 560833 295788
rect 560878 295784 560918 295810
rect 560767 295738 560783 295772
rect 560817 295738 560833 295772
rect 560767 295722 560833 295738
rect 569281 305882 569347 305898
rect 569281 305848 569297 305882
rect 569331 305848 569347 305882
rect 569196 305810 569236 305836
rect 569281 305832 569347 305848
rect 569477 305882 569543 305898
rect 569477 305848 569493 305882
rect 569527 305848 569543 305882
rect 569294 305810 569334 305832
rect 569392 305810 569432 305836
rect 569477 305832 569543 305848
rect 569673 305882 569739 305898
rect 569673 305848 569689 305882
rect 569723 305848 569739 305882
rect 569490 305810 569530 305832
rect 569588 305810 569628 305836
rect 569673 305832 569739 305848
rect 569869 305882 569935 305898
rect 569869 305848 569885 305882
rect 569919 305848 569935 305882
rect 569686 305810 569726 305832
rect 569784 305810 569824 305836
rect 569869 305832 569935 305848
rect 570065 305882 570131 305898
rect 570065 305848 570081 305882
rect 570115 305848 570131 305882
rect 569882 305810 569922 305832
rect 569980 305810 570020 305836
rect 570065 305832 570131 305848
rect 570078 305810 570118 305832
rect 569196 295788 569236 295810
rect 569183 295772 569249 295788
rect 569294 295784 569334 295810
rect 569392 295788 569432 295810
rect 569183 295738 569199 295772
rect 569233 295738 569249 295772
rect 569183 295722 569249 295738
rect 569379 295772 569445 295788
rect 569490 295784 569530 295810
rect 569588 295788 569628 295810
rect 569379 295738 569395 295772
rect 569429 295738 569445 295772
rect 569379 295722 569445 295738
rect 569575 295772 569641 295788
rect 569686 295784 569726 295810
rect 569784 295788 569824 295810
rect 569575 295738 569591 295772
rect 569625 295738 569641 295772
rect 569575 295722 569641 295738
rect 569771 295772 569837 295788
rect 569882 295784 569922 295810
rect 569980 295788 570020 295810
rect 569771 295738 569787 295772
rect 569821 295738 569837 295772
rect 569771 295722 569837 295738
rect 569967 295772 570033 295788
rect 570078 295784 570118 295810
rect 569967 295738 569983 295772
rect 570017 295738 570033 295772
rect 569967 295722 570033 295738
rect 536271 294722 536368 294738
rect 536271 294654 536287 294722
rect 536321 294654 536368 294722
rect 536271 294638 536368 294654
rect 537368 294722 537465 294738
rect 537368 294654 537415 294722
rect 537449 294654 537465 294722
rect 537368 294638 537465 294654
rect 537507 294722 537604 294738
rect 537507 294654 537523 294722
rect 537557 294654 537604 294722
rect 537507 294638 537604 294654
rect 538604 294722 538701 294738
rect 538604 294654 538651 294722
rect 538685 294654 538701 294722
rect 538604 294638 538701 294654
rect 538743 294722 538840 294738
rect 538743 294654 538759 294722
rect 538793 294654 538840 294722
rect 538743 294638 538840 294654
rect 539840 294722 539937 294738
rect 539840 294654 539887 294722
rect 539921 294654 539937 294722
rect 539840 294638 539937 294654
rect 539979 294722 540076 294738
rect 539979 294654 539995 294722
rect 540029 294654 540076 294722
rect 539979 294638 540076 294654
rect 541076 294722 541173 294738
rect 541076 294654 541123 294722
rect 541157 294654 541173 294722
rect 541076 294638 541173 294654
rect 541215 294722 541312 294738
rect 541215 294654 541231 294722
rect 541265 294654 541312 294722
rect 541215 294638 541312 294654
rect 542312 294722 542409 294738
rect 542312 294654 542359 294722
rect 542393 294654 542409 294722
rect 542312 294638 542409 294654
rect 542451 294722 542548 294738
rect 542451 294654 542467 294722
rect 542501 294654 542548 294722
rect 542451 294638 542548 294654
rect 543548 294722 543645 294738
rect 543548 294654 543595 294722
rect 543629 294654 543645 294722
rect 543548 294638 543645 294654
rect 543687 294722 543784 294738
rect 543687 294654 543703 294722
rect 543737 294654 543784 294722
rect 543687 294638 543784 294654
rect 544784 294722 544881 294738
rect 544784 294654 544831 294722
rect 544865 294654 544881 294722
rect 544784 294638 544881 294654
rect 5902 293918 5968 293931
rect 5902 293915 5990 293918
rect 5902 293881 5918 293915
rect 5952 293881 5990 293915
rect 5902 293878 5990 293881
rect 15990 293878 16016 293918
rect 5902 293865 5968 293878
rect 16012 293820 16078 293833
rect 5964 293780 5990 293820
rect 15990 293817 16078 293820
rect 15990 293783 16028 293817
rect 16062 293783 16078 293817
rect 15990 293780 16078 293783
rect 5902 293722 5968 293735
rect 16012 293767 16078 293780
rect 5902 293719 5990 293722
rect 5902 293685 5918 293719
rect 5952 293685 5990 293719
rect 5902 293682 5990 293685
rect 15990 293682 16016 293722
rect 5902 293669 5968 293682
rect 16012 293624 16078 293637
rect 5964 293584 5990 293624
rect 15990 293621 16078 293624
rect 15990 293587 16028 293621
rect 16062 293587 16078 293621
rect 15990 293584 16078 293587
rect 5902 293526 5968 293539
rect 16012 293571 16078 293584
rect 5902 293523 5990 293526
rect 5902 293489 5918 293523
rect 5952 293489 5990 293523
rect 5902 293486 5990 293489
rect 15990 293486 16016 293526
rect 5902 293473 5968 293486
rect 16012 293428 16078 293441
rect 5964 293388 5990 293428
rect 15990 293425 16078 293428
rect 15990 293391 16028 293425
rect 16062 293391 16078 293425
rect 15990 293388 16078 293391
rect 5902 293330 5968 293343
rect 16012 293375 16078 293388
rect 5902 293327 5990 293330
rect 5902 293293 5918 293327
rect 5952 293293 5990 293327
rect 5902 293290 5990 293293
rect 15990 293290 16016 293330
rect 5902 293277 5968 293290
rect 16012 293232 16078 293245
rect 5964 293192 5990 293232
rect 15990 293229 16078 293232
rect 15990 293195 16028 293229
rect 16062 293195 16078 293229
rect 15990 293192 16078 293195
rect 5902 293134 5968 293147
rect 16012 293179 16078 293192
rect 5902 293131 5990 293134
rect 5902 293097 5918 293131
rect 5952 293097 5990 293131
rect 5902 293094 5990 293097
rect 15990 293094 16016 293134
rect 5902 293081 5968 293094
rect 16012 293036 16078 293049
rect 5964 292996 5990 293036
rect 15990 293033 16078 293036
rect 15990 292999 16028 293033
rect 16062 292999 16078 293033
rect 15990 292996 16078 292999
rect 16012 292983 16078 292996
rect 536271 294182 536368 294198
rect 536271 294114 536287 294182
rect 536321 294114 536368 294182
rect 536271 294098 536368 294114
rect 537368 294182 537465 294198
rect 537368 294114 537415 294182
rect 537449 294114 537465 294182
rect 537368 294098 537465 294114
rect 537507 294182 537604 294198
rect 537507 294114 537523 294182
rect 537557 294114 537604 294182
rect 537507 294098 537604 294114
rect 538604 294182 538701 294198
rect 538604 294114 538651 294182
rect 538685 294114 538701 294182
rect 538604 294098 538701 294114
rect 538743 294182 538840 294198
rect 538743 294114 538759 294182
rect 538793 294114 538840 294182
rect 538743 294098 538840 294114
rect 539840 294182 539937 294198
rect 539840 294114 539887 294182
rect 539921 294114 539937 294182
rect 539840 294098 539937 294114
rect 539979 294182 540076 294198
rect 539979 294114 539995 294182
rect 540029 294114 540076 294182
rect 539979 294098 540076 294114
rect 541076 294182 541173 294198
rect 541076 294114 541123 294182
rect 541157 294114 541173 294182
rect 541076 294098 541173 294114
rect 541215 294182 541312 294198
rect 541215 294114 541231 294182
rect 541265 294114 541312 294182
rect 541215 294098 541312 294114
rect 542312 294182 542409 294198
rect 542312 294114 542359 294182
rect 542393 294114 542409 294182
rect 542312 294098 542409 294114
rect 542451 294182 542548 294198
rect 542451 294114 542467 294182
rect 542501 294114 542548 294182
rect 542451 294098 542548 294114
rect 543548 294182 543645 294198
rect 543548 294114 543595 294182
rect 543629 294114 543645 294182
rect 543548 294098 543645 294114
rect 543687 294182 543784 294198
rect 543687 294114 543703 294182
rect 543737 294114 543784 294182
rect 543687 294098 543784 294114
rect 544784 294182 544881 294198
rect 544784 294114 544831 294182
rect 544865 294114 544881 294182
rect 544784 294098 544881 294114
rect 536271 293642 536368 293658
rect 536271 293574 536287 293642
rect 536321 293574 536368 293642
rect 536271 293558 536368 293574
rect 537368 293642 537465 293658
rect 537368 293574 537415 293642
rect 537449 293574 537465 293642
rect 537368 293558 537465 293574
rect 537507 293642 537604 293658
rect 537507 293574 537523 293642
rect 537557 293574 537604 293642
rect 537507 293558 537604 293574
rect 538604 293642 538701 293658
rect 538604 293574 538651 293642
rect 538685 293574 538701 293642
rect 538604 293558 538701 293574
rect 538743 293642 538840 293658
rect 538743 293574 538759 293642
rect 538793 293574 538840 293642
rect 538743 293558 538840 293574
rect 539840 293642 539937 293658
rect 539840 293574 539887 293642
rect 539921 293574 539937 293642
rect 539840 293558 539937 293574
rect 539979 293642 540076 293658
rect 539979 293574 539995 293642
rect 540029 293574 540076 293642
rect 539979 293558 540076 293574
rect 541076 293642 541173 293658
rect 541076 293574 541123 293642
rect 541157 293574 541173 293642
rect 541076 293558 541173 293574
rect 541215 293642 541312 293658
rect 541215 293574 541231 293642
rect 541265 293574 541312 293642
rect 541215 293558 541312 293574
rect 542312 293642 542409 293658
rect 542312 293574 542359 293642
rect 542393 293574 542409 293642
rect 542312 293558 542409 293574
rect 542451 293642 542548 293658
rect 542451 293574 542467 293642
rect 542501 293574 542548 293642
rect 542451 293558 542548 293574
rect 543548 293642 543645 293658
rect 543548 293574 543595 293642
rect 543629 293574 543645 293642
rect 543548 293558 543645 293574
rect 543687 293642 543784 293658
rect 543687 293574 543703 293642
rect 543737 293574 543784 293642
rect 543687 293558 543784 293574
rect 544784 293642 544881 293658
rect 544784 293574 544831 293642
rect 544865 293574 544881 293642
rect 544784 293558 544881 293574
rect 536271 293102 536368 293118
rect 536271 293034 536287 293102
rect 536321 293034 536368 293102
rect 536271 293018 536368 293034
rect 537368 293102 537465 293118
rect 537368 293034 537415 293102
rect 537449 293034 537465 293102
rect 537368 293018 537465 293034
rect 537507 293102 537604 293118
rect 537507 293034 537523 293102
rect 537557 293034 537604 293102
rect 537507 293018 537604 293034
rect 538604 293102 538701 293118
rect 538604 293034 538651 293102
rect 538685 293034 538701 293102
rect 538604 293018 538701 293034
rect 538743 293102 538840 293118
rect 538743 293034 538759 293102
rect 538793 293034 538840 293102
rect 538743 293018 538840 293034
rect 539840 293102 539937 293118
rect 539840 293034 539887 293102
rect 539921 293034 539937 293102
rect 539840 293018 539937 293034
rect 539979 293102 540076 293118
rect 539979 293034 539995 293102
rect 540029 293034 540076 293102
rect 539979 293018 540076 293034
rect 541076 293102 541173 293118
rect 541076 293034 541123 293102
rect 541157 293034 541173 293102
rect 541076 293018 541173 293034
rect 541215 293102 541312 293118
rect 541215 293034 541231 293102
rect 541265 293034 541312 293102
rect 541215 293018 541312 293034
rect 542312 293102 542409 293118
rect 542312 293034 542359 293102
rect 542393 293034 542409 293102
rect 542312 293018 542409 293034
rect 542451 293102 542548 293118
rect 542451 293034 542467 293102
rect 542501 293034 542548 293102
rect 542451 293018 542548 293034
rect 543548 293102 543645 293118
rect 543548 293034 543595 293102
rect 543629 293034 543645 293102
rect 543548 293018 543645 293034
rect 543687 293102 543784 293118
rect 543687 293034 543703 293102
rect 543737 293034 543784 293102
rect 543687 293018 543784 293034
rect 544784 293102 544881 293118
rect 544784 293034 544831 293102
rect 544865 293034 544881 293102
rect 544784 293018 544881 293034
rect 536271 292522 536368 292538
rect 536271 292454 536287 292522
rect 536321 292454 536368 292522
rect 536271 292438 536368 292454
rect 537368 292522 537465 292538
rect 537368 292454 537415 292522
rect 537449 292454 537465 292522
rect 537368 292438 537465 292454
rect 537507 292522 537604 292538
rect 537507 292454 537523 292522
rect 537557 292454 537604 292522
rect 537507 292438 537604 292454
rect 538604 292522 538701 292538
rect 538604 292454 538651 292522
rect 538685 292454 538701 292522
rect 538604 292438 538701 292454
rect 538743 292522 538840 292538
rect 538743 292454 538759 292522
rect 538793 292454 538840 292522
rect 538743 292438 538840 292454
rect 539840 292522 539937 292538
rect 539840 292454 539887 292522
rect 539921 292454 539937 292522
rect 539840 292438 539937 292454
rect 539979 292522 540076 292538
rect 539979 292454 539995 292522
rect 540029 292454 540076 292522
rect 539979 292438 540076 292454
rect 541076 292522 541173 292538
rect 541076 292454 541123 292522
rect 541157 292454 541173 292522
rect 541076 292438 541173 292454
rect 541215 292522 541312 292538
rect 541215 292454 541231 292522
rect 541265 292454 541312 292522
rect 541215 292438 541312 292454
rect 542312 292522 542409 292538
rect 542312 292454 542359 292522
rect 542393 292454 542409 292522
rect 542312 292438 542409 292454
rect 542451 292522 542548 292538
rect 542451 292454 542467 292522
rect 542501 292454 542548 292522
rect 542451 292438 542548 292454
rect 543548 292522 543645 292538
rect 543548 292454 543595 292522
rect 543629 292454 543645 292522
rect 543548 292438 543645 292454
rect 543687 292522 543784 292538
rect 543687 292454 543703 292522
rect 543737 292454 543784 292522
rect 543687 292438 543784 292454
rect 544784 292522 544881 292538
rect 544784 292454 544831 292522
rect 544865 292454 544881 292522
rect 544784 292438 544881 292454
rect 536271 291942 536368 291958
rect 536271 291874 536287 291942
rect 536321 291874 536368 291942
rect 536271 291858 536368 291874
rect 537368 291942 537465 291958
rect 537368 291874 537415 291942
rect 537449 291874 537465 291942
rect 537368 291858 537465 291874
rect 537507 291942 537604 291958
rect 537507 291874 537523 291942
rect 537557 291874 537604 291942
rect 537507 291858 537604 291874
rect 538604 291942 538701 291958
rect 538604 291874 538651 291942
rect 538685 291874 538701 291942
rect 538604 291858 538701 291874
rect 538743 291942 538840 291958
rect 538743 291874 538759 291942
rect 538793 291874 538840 291942
rect 538743 291858 538840 291874
rect 539840 291942 539937 291958
rect 539840 291874 539887 291942
rect 539921 291874 539937 291942
rect 539840 291858 539937 291874
rect 539979 291942 540076 291958
rect 539979 291874 539995 291942
rect 540029 291874 540076 291942
rect 539979 291858 540076 291874
rect 541076 291942 541173 291958
rect 541076 291874 541123 291942
rect 541157 291874 541173 291942
rect 541076 291858 541173 291874
rect 541215 291942 541312 291958
rect 541215 291874 541231 291942
rect 541265 291874 541312 291942
rect 541215 291858 541312 291874
rect 542312 291942 542409 291958
rect 542312 291874 542359 291942
rect 542393 291874 542409 291942
rect 542312 291858 542409 291874
rect 542451 291942 542548 291958
rect 542451 291874 542467 291942
rect 542501 291874 542548 291942
rect 542451 291858 542548 291874
rect 543548 291942 543645 291958
rect 543548 291874 543595 291942
rect 543629 291874 543645 291942
rect 543548 291858 543645 291874
rect 543687 291942 543784 291958
rect 543687 291874 543703 291942
rect 543737 291874 543784 291942
rect 543687 291858 543784 291874
rect 544784 291942 544881 291958
rect 544784 291874 544831 291942
rect 544865 291874 544881 291942
rect 544784 291858 544881 291874
rect 534431 291402 534528 291418
rect 534431 291334 534447 291402
rect 534481 291334 534528 291402
rect 534431 291318 534528 291334
rect 535528 291402 535625 291418
rect 535528 291334 535575 291402
rect 535609 291334 535625 291402
rect 535528 291318 535625 291334
rect 535667 291402 535764 291418
rect 535667 291334 535683 291402
rect 535717 291334 535764 291402
rect 535667 291318 535764 291334
rect 536764 291402 536861 291418
rect 536764 291334 536811 291402
rect 536845 291334 536861 291402
rect 536764 291318 536861 291334
rect 536903 291402 537000 291418
rect 536903 291334 536919 291402
rect 536953 291334 537000 291402
rect 536903 291318 537000 291334
rect 538000 291402 538097 291418
rect 538000 291334 538047 291402
rect 538081 291334 538097 291402
rect 538000 291318 538097 291334
rect 538139 291402 538236 291418
rect 538139 291334 538155 291402
rect 538189 291334 538236 291402
rect 538139 291318 538236 291334
rect 539236 291402 539333 291418
rect 539236 291334 539283 291402
rect 539317 291334 539333 291402
rect 539236 291318 539333 291334
rect 539375 291402 539472 291418
rect 539375 291334 539391 291402
rect 539425 291334 539472 291402
rect 539375 291318 539472 291334
rect 540472 291402 540569 291418
rect 540472 291334 540519 291402
rect 540553 291334 540569 291402
rect 540472 291318 540569 291334
rect 540611 291402 540708 291418
rect 540611 291334 540627 291402
rect 540661 291334 540708 291402
rect 540611 291318 540708 291334
rect 541708 291402 541805 291418
rect 541708 291334 541755 291402
rect 541789 291334 541805 291402
rect 541708 291318 541805 291334
rect 541847 291402 541944 291418
rect 541847 291334 541863 291402
rect 541897 291334 541944 291402
rect 541847 291318 541944 291334
rect 542944 291402 543041 291418
rect 542944 291334 542991 291402
rect 543025 291334 543041 291402
rect 542944 291318 543041 291334
rect 543083 291402 543180 291418
rect 543083 291334 543099 291402
rect 543133 291334 543180 291402
rect 543083 291318 543180 291334
rect 544180 291402 544277 291418
rect 544180 291334 544227 291402
rect 544261 291334 544277 291402
rect 544180 291318 544277 291334
rect 544319 291402 544416 291418
rect 544319 291334 544335 291402
rect 544369 291334 544416 291402
rect 544319 291318 544416 291334
rect 545416 291402 545513 291418
rect 545416 291334 545463 291402
rect 545497 291334 545513 291402
rect 545416 291318 545513 291334
rect 545555 291402 545652 291418
rect 545555 291334 545571 291402
rect 545605 291334 545652 291402
rect 545555 291318 545652 291334
rect 546652 291402 546749 291418
rect 546652 291334 546699 291402
rect 546733 291334 546749 291402
rect 546652 291318 546749 291334
rect 534431 290862 534528 290878
rect 534431 290794 534447 290862
rect 534481 290794 534528 290862
rect 534431 290778 534528 290794
rect 535528 290862 535625 290878
rect 535528 290794 535575 290862
rect 535609 290794 535625 290862
rect 535528 290778 535625 290794
rect 535667 290862 535764 290878
rect 535667 290794 535683 290862
rect 535717 290794 535764 290862
rect 535667 290778 535764 290794
rect 536764 290862 536861 290878
rect 536764 290794 536811 290862
rect 536845 290794 536861 290862
rect 536764 290778 536861 290794
rect 536903 290862 537000 290878
rect 536903 290794 536919 290862
rect 536953 290794 537000 290862
rect 536903 290778 537000 290794
rect 538000 290862 538097 290878
rect 538000 290794 538047 290862
rect 538081 290794 538097 290862
rect 538000 290778 538097 290794
rect 538139 290862 538236 290878
rect 538139 290794 538155 290862
rect 538189 290794 538236 290862
rect 538139 290778 538236 290794
rect 539236 290862 539333 290878
rect 539236 290794 539283 290862
rect 539317 290794 539333 290862
rect 539236 290778 539333 290794
rect 539375 290862 539472 290878
rect 539375 290794 539391 290862
rect 539425 290794 539472 290862
rect 539375 290778 539472 290794
rect 540472 290862 540569 290878
rect 540472 290794 540519 290862
rect 540553 290794 540569 290862
rect 540472 290778 540569 290794
rect 540611 290862 540708 290878
rect 540611 290794 540627 290862
rect 540661 290794 540708 290862
rect 540611 290778 540708 290794
rect 541708 290862 541805 290878
rect 541708 290794 541755 290862
rect 541789 290794 541805 290862
rect 541708 290778 541805 290794
rect 541847 290862 541944 290878
rect 541847 290794 541863 290862
rect 541897 290794 541944 290862
rect 541847 290778 541944 290794
rect 542944 290862 543041 290878
rect 542944 290794 542991 290862
rect 543025 290794 543041 290862
rect 542944 290778 543041 290794
rect 543083 290862 543180 290878
rect 543083 290794 543099 290862
rect 543133 290794 543180 290862
rect 543083 290778 543180 290794
rect 544180 290862 544277 290878
rect 544180 290794 544227 290862
rect 544261 290794 544277 290862
rect 544180 290778 544277 290794
rect 544319 290862 544416 290878
rect 544319 290794 544335 290862
rect 544369 290794 544416 290862
rect 544319 290778 544416 290794
rect 545416 290862 545513 290878
rect 545416 290794 545463 290862
rect 545497 290794 545513 290862
rect 545416 290778 545513 290794
rect 545555 290862 545652 290878
rect 545555 290794 545571 290862
rect 545605 290794 545652 290862
rect 545555 290778 545652 290794
rect 546652 290862 546749 290878
rect 546652 290794 546699 290862
rect 546733 290794 546749 290862
rect 546652 290778 546749 290794
rect 534431 290322 534528 290338
rect 534431 290254 534447 290322
rect 534481 290254 534528 290322
rect 534431 290238 534528 290254
rect 535528 290322 535625 290338
rect 535528 290254 535575 290322
rect 535609 290254 535625 290322
rect 535528 290238 535625 290254
rect 535667 290322 535764 290338
rect 535667 290254 535683 290322
rect 535717 290254 535764 290322
rect 535667 290238 535764 290254
rect 536764 290322 536861 290338
rect 536764 290254 536811 290322
rect 536845 290254 536861 290322
rect 536764 290238 536861 290254
rect 536903 290322 537000 290338
rect 536903 290254 536919 290322
rect 536953 290254 537000 290322
rect 536903 290238 537000 290254
rect 538000 290322 538097 290338
rect 538000 290254 538047 290322
rect 538081 290254 538097 290322
rect 538000 290238 538097 290254
rect 538139 290322 538236 290338
rect 538139 290254 538155 290322
rect 538189 290254 538236 290322
rect 538139 290238 538236 290254
rect 539236 290322 539333 290338
rect 539236 290254 539283 290322
rect 539317 290254 539333 290322
rect 539236 290238 539333 290254
rect 539375 290322 539472 290338
rect 539375 290254 539391 290322
rect 539425 290254 539472 290322
rect 539375 290238 539472 290254
rect 540472 290322 540569 290338
rect 540472 290254 540519 290322
rect 540553 290254 540569 290322
rect 540472 290238 540569 290254
rect 540611 290322 540708 290338
rect 540611 290254 540627 290322
rect 540661 290254 540708 290322
rect 540611 290238 540708 290254
rect 541708 290322 541805 290338
rect 541708 290254 541755 290322
rect 541789 290254 541805 290322
rect 541708 290238 541805 290254
rect 541847 290322 541944 290338
rect 541847 290254 541863 290322
rect 541897 290254 541944 290322
rect 541847 290238 541944 290254
rect 542944 290322 543041 290338
rect 542944 290254 542991 290322
rect 543025 290254 543041 290322
rect 542944 290238 543041 290254
rect 543083 290322 543180 290338
rect 543083 290254 543099 290322
rect 543133 290254 543180 290322
rect 543083 290238 543180 290254
rect 544180 290322 544277 290338
rect 544180 290254 544227 290322
rect 544261 290254 544277 290322
rect 544180 290238 544277 290254
rect 544319 290322 544416 290338
rect 544319 290254 544335 290322
rect 544369 290254 544416 290322
rect 544319 290238 544416 290254
rect 545416 290322 545513 290338
rect 545416 290254 545463 290322
rect 545497 290254 545513 290322
rect 545416 290238 545513 290254
rect 545555 290322 545652 290338
rect 545555 290254 545571 290322
rect 545605 290254 545652 290322
rect 545555 290238 545652 290254
rect 546652 290322 546749 290338
rect 546652 290254 546699 290322
rect 546733 290254 546749 290322
rect 546652 290238 546749 290254
rect 534431 289782 534528 289798
rect 534431 289714 534447 289782
rect 534481 289714 534528 289782
rect 534431 289698 534528 289714
rect 535528 289782 535625 289798
rect 535528 289714 535575 289782
rect 535609 289714 535625 289782
rect 535528 289698 535625 289714
rect 535667 289782 535764 289798
rect 535667 289714 535683 289782
rect 535717 289714 535764 289782
rect 535667 289698 535764 289714
rect 536764 289782 536861 289798
rect 536764 289714 536811 289782
rect 536845 289714 536861 289782
rect 536764 289698 536861 289714
rect 536903 289782 537000 289798
rect 536903 289714 536919 289782
rect 536953 289714 537000 289782
rect 536903 289698 537000 289714
rect 538000 289782 538097 289798
rect 538000 289714 538047 289782
rect 538081 289714 538097 289782
rect 538000 289698 538097 289714
rect 538139 289782 538236 289798
rect 538139 289714 538155 289782
rect 538189 289714 538236 289782
rect 538139 289698 538236 289714
rect 539236 289782 539333 289798
rect 539236 289714 539283 289782
rect 539317 289714 539333 289782
rect 539236 289698 539333 289714
rect 539375 289782 539472 289798
rect 539375 289714 539391 289782
rect 539425 289714 539472 289782
rect 539375 289698 539472 289714
rect 540472 289782 540569 289798
rect 540472 289714 540519 289782
rect 540553 289714 540569 289782
rect 540472 289698 540569 289714
rect 540611 289782 540708 289798
rect 540611 289714 540627 289782
rect 540661 289714 540708 289782
rect 540611 289698 540708 289714
rect 541708 289782 541805 289798
rect 541708 289714 541755 289782
rect 541789 289714 541805 289782
rect 541708 289698 541805 289714
rect 541847 289782 541944 289798
rect 541847 289714 541863 289782
rect 541897 289714 541944 289782
rect 541847 289698 541944 289714
rect 542944 289782 543041 289798
rect 542944 289714 542991 289782
rect 543025 289714 543041 289782
rect 542944 289698 543041 289714
rect 543083 289782 543180 289798
rect 543083 289714 543099 289782
rect 543133 289714 543180 289782
rect 543083 289698 543180 289714
rect 544180 289782 544277 289798
rect 544180 289714 544227 289782
rect 544261 289714 544277 289782
rect 544180 289698 544277 289714
rect 544319 289782 544416 289798
rect 544319 289714 544335 289782
rect 544369 289714 544416 289782
rect 544319 289698 544416 289714
rect 545416 289782 545513 289798
rect 545416 289714 545463 289782
rect 545497 289714 545513 289782
rect 545416 289698 545513 289714
rect 545555 289782 545652 289798
rect 545555 289714 545571 289782
rect 545605 289714 545652 289782
rect 545555 289698 545652 289714
rect 546652 289782 546749 289798
rect 546652 289714 546699 289782
rect 546733 289714 546749 289782
rect 546652 289698 546749 289714
rect 536371 289002 536459 289018
rect 536371 288934 536387 289002
rect 536421 288934 536459 289002
rect 536371 288918 536459 288934
rect 537459 289002 537547 289018
rect 537459 288934 537497 289002
rect 537531 288934 537547 289002
rect 537459 288918 537547 288934
rect 537589 289002 537677 289018
rect 537589 288934 537605 289002
rect 537639 288934 537677 289002
rect 537589 288918 537677 288934
rect 538677 289002 538765 289018
rect 538677 288934 538715 289002
rect 538749 288934 538765 289002
rect 538677 288918 538765 288934
rect 538807 289002 538895 289018
rect 538807 288934 538823 289002
rect 538857 288934 538895 289002
rect 538807 288918 538895 288934
rect 539895 289002 539983 289018
rect 539895 288934 539933 289002
rect 539967 288934 539983 289002
rect 539895 288918 539983 288934
rect 540025 289002 540113 289018
rect 540025 288934 540041 289002
rect 540075 288934 540113 289002
rect 540025 288918 540113 288934
rect 541113 289002 541201 289018
rect 541113 288934 541151 289002
rect 541185 288934 541201 289002
rect 541113 288918 541201 288934
rect 541243 289002 541331 289018
rect 541243 288934 541259 289002
rect 541293 288934 541331 289002
rect 541243 288918 541331 288934
rect 542331 289002 542419 289018
rect 542331 288934 542369 289002
rect 542403 288934 542419 289002
rect 542331 288918 542419 288934
rect 542461 289002 542549 289018
rect 542461 288934 542477 289002
rect 542511 288934 542549 289002
rect 542461 288918 542549 288934
rect 543549 289002 543637 289018
rect 543549 288934 543587 289002
rect 543621 288934 543637 289002
rect 543549 288918 543637 288934
rect 543679 289002 543767 289018
rect 543679 288934 543695 289002
rect 543729 288934 543767 289002
rect 543679 288918 543767 288934
rect 544767 289002 544855 289018
rect 544767 288934 544805 289002
rect 544839 288934 544855 289002
rect 544767 288918 544855 288934
rect 536371 288502 536459 288518
rect 536371 288434 536387 288502
rect 536421 288434 536459 288502
rect 536371 288418 536459 288434
rect 537459 288502 537547 288518
rect 537459 288434 537497 288502
rect 537531 288434 537547 288502
rect 537459 288418 537547 288434
rect 537589 288502 537677 288518
rect 537589 288434 537605 288502
rect 537639 288434 537677 288502
rect 537589 288418 537677 288434
rect 538677 288502 538765 288518
rect 538677 288434 538715 288502
rect 538749 288434 538765 288502
rect 538677 288418 538765 288434
rect 538807 288502 538895 288518
rect 538807 288434 538823 288502
rect 538857 288434 538895 288502
rect 538807 288418 538895 288434
rect 539895 288502 539983 288518
rect 539895 288434 539933 288502
rect 539967 288434 539983 288502
rect 539895 288418 539983 288434
rect 540025 288502 540113 288518
rect 540025 288434 540041 288502
rect 540075 288434 540113 288502
rect 540025 288418 540113 288434
rect 541113 288502 541201 288518
rect 541113 288434 541151 288502
rect 541185 288434 541201 288502
rect 541113 288418 541201 288434
rect 541243 288502 541331 288518
rect 541243 288434 541259 288502
rect 541293 288434 541331 288502
rect 541243 288418 541331 288434
rect 542331 288502 542419 288518
rect 542331 288434 542369 288502
rect 542403 288434 542419 288502
rect 542331 288418 542419 288434
rect 542461 288502 542549 288518
rect 542461 288434 542477 288502
rect 542511 288434 542549 288502
rect 542461 288418 542549 288434
rect 543549 288502 543637 288518
rect 543549 288434 543587 288502
rect 543621 288434 543637 288502
rect 543549 288418 543637 288434
rect 543679 288502 543767 288518
rect 543679 288434 543695 288502
rect 543729 288434 543767 288502
rect 543679 288418 543767 288434
rect 544767 288502 544855 288518
rect 544767 288434 544805 288502
rect 544839 288434 544855 288502
rect 544767 288418 544855 288434
rect 536931 288002 537019 288018
rect 536931 287834 536947 288002
rect 536981 287834 537019 288002
rect 536931 287818 537019 287834
rect 538019 288002 538107 288018
rect 538019 287834 538057 288002
rect 538091 287834 538107 288002
rect 538019 287818 538107 287834
rect 538149 288002 538237 288018
rect 538149 287834 538165 288002
rect 538199 287834 538237 288002
rect 538149 287818 538237 287834
rect 539237 288002 539325 288018
rect 539237 287834 539275 288002
rect 539309 287834 539325 288002
rect 539237 287818 539325 287834
rect 539367 288002 539455 288018
rect 539367 287834 539383 288002
rect 539417 287834 539455 288002
rect 539367 287818 539455 287834
rect 540455 288002 540543 288018
rect 540455 287834 540493 288002
rect 540527 287834 540543 288002
rect 540455 287818 540543 287834
rect 540585 288002 540673 288018
rect 540585 287834 540601 288002
rect 540635 287834 540673 288002
rect 540585 287818 540673 287834
rect 541673 288002 541761 288018
rect 541673 287834 541711 288002
rect 541745 287834 541761 288002
rect 541673 287818 541761 287834
rect 541803 288002 541891 288018
rect 541803 287834 541819 288002
rect 541853 287834 541891 288002
rect 541803 287818 541891 287834
rect 542891 288002 542979 288018
rect 542891 287834 542929 288002
rect 542963 287834 542979 288002
rect 542891 287818 542979 287834
rect 543021 288002 543109 288018
rect 543021 287834 543037 288002
rect 543071 287834 543109 288002
rect 543021 287818 543109 287834
rect 544109 288002 544197 288018
rect 544109 287834 544147 288002
rect 544181 287834 544197 288002
rect 544109 287818 544197 287834
rect 568202 288698 568268 288711
rect 568202 288695 568290 288698
rect 568202 288661 568218 288695
rect 568252 288661 568290 288695
rect 568202 288658 568290 288661
rect 578290 288658 578316 288698
rect 568202 288645 568268 288658
rect 578312 288600 578378 288613
rect 568264 288560 568290 288600
rect 578290 288597 578378 288600
rect 578290 288563 578328 288597
rect 578362 288563 578378 288597
rect 578290 288560 578378 288563
rect 568202 288502 568268 288515
rect 578312 288547 578378 288560
rect 568202 288499 568290 288502
rect 568202 288465 568218 288499
rect 568252 288465 568290 288499
rect 568202 288462 568290 288465
rect 578290 288462 578316 288502
rect 568202 288449 568268 288462
rect 578312 288404 578378 288417
rect 568264 288364 568290 288404
rect 578290 288401 578378 288404
rect 578290 288367 578328 288401
rect 578362 288367 578378 288401
rect 578290 288364 578378 288367
rect 568202 288306 568268 288319
rect 578312 288351 578378 288364
rect 568202 288303 568290 288306
rect 568202 288269 568218 288303
rect 568252 288269 568290 288303
rect 568202 288266 568290 288269
rect 578290 288266 578316 288306
rect 568202 288253 568268 288266
rect 578312 288208 578378 288221
rect 568264 288168 568290 288208
rect 578290 288205 578378 288208
rect 578290 288171 578328 288205
rect 578362 288171 578378 288205
rect 578290 288168 578378 288171
rect 568202 288110 568268 288123
rect 578312 288155 578378 288168
rect 568202 288107 568290 288110
rect 568202 288073 568218 288107
rect 568252 288073 568290 288107
rect 568202 288070 568290 288073
rect 578290 288070 578316 288110
rect 568202 288057 568268 288070
rect 578312 288012 578378 288025
rect 568264 287972 568290 288012
rect 578290 288009 578378 288012
rect 578290 287975 578328 288009
rect 578362 287975 578378 288009
rect 578290 287972 578378 287975
rect 568202 287914 568268 287927
rect 578312 287959 578378 287972
rect 568202 287911 568290 287914
rect 568202 287877 568218 287911
rect 568252 287877 568290 287911
rect 568202 287874 568290 287877
rect 578290 287874 578316 287914
rect 568202 287861 568268 287874
rect 578312 287816 578378 287829
rect 568264 287776 568290 287816
rect 578290 287813 578378 287816
rect 578290 287779 578328 287813
rect 578362 287779 578378 287813
rect 578290 287776 578378 287779
rect 578312 287763 578378 287776
rect 536931 287382 537019 287398
rect 536931 287214 536947 287382
rect 536981 287214 537019 287382
rect 536931 287198 537019 287214
rect 538019 287382 538107 287398
rect 538019 287214 538057 287382
rect 538091 287214 538107 287382
rect 538019 287198 538107 287214
rect 538149 287382 538237 287398
rect 538149 287214 538165 287382
rect 538199 287214 538237 287382
rect 538149 287198 538237 287214
rect 539237 287382 539325 287398
rect 539237 287214 539275 287382
rect 539309 287214 539325 287382
rect 539237 287198 539325 287214
rect 539367 287382 539455 287398
rect 539367 287214 539383 287382
rect 539417 287214 539455 287382
rect 539367 287198 539455 287214
rect 540455 287382 540543 287398
rect 540455 287214 540493 287382
rect 540527 287214 540543 287382
rect 540455 287198 540543 287214
rect 540585 287382 540673 287398
rect 540585 287214 540601 287382
rect 540635 287214 540673 287382
rect 540585 287198 540673 287214
rect 541673 287382 541761 287398
rect 541673 287214 541711 287382
rect 541745 287214 541761 287382
rect 541673 287198 541761 287214
rect 541803 287382 541891 287398
rect 541803 287214 541819 287382
rect 541853 287214 541891 287382
rect 541803 287198 541891 287214
rect 542891 287382 542979 287398
rect 542891 287214 542929 287382
rect 542963 287214 542979 287382
rect 542891 287198 542979 287214
rect 543021 287382 543109 287398
rect 543021 287214 543037 287382
rect 543071 287214 543109 287382
rect 543021 287198 543109 287214
rect 544109 287382 544197 287398
rect 544109 287214 544147 287382
rect 544181 287214 544197 287382
rect 544109 287198 544197 287214
rect 536371 286782 536459 286798
rect 536371 286614 536387 286782
rect 536421 286614 536459 286782
rect 536371 286598 536459 286614
rect 537459 286782 537547 286798
rect 537459 286614 537497 286782
rect 537531 286614 537547 286782
rect 537459 286598 537547 286614
rect 537589 286782 537677 286798
rect 537589 286614 537605 286782
rect 537639 286614 537677 286782
rect 537589 286598 537677 286614
rect 538677 286782 538765 286798
rect 538677 286614 538715 286782
rect 538749 286614 538765 286782
rect 538677 286598 538765 286614
rect 538807 286782 538895 286798
rect 538807 286614 538823 286782
rect 538857 286614 538895 286782
rect 538807 286598 538895 286614
rect 539895 286782 539983 286798
rect 539895 286614 539933 286782
rect 539967 286614 539983 286782
rect 539895 286598 539983 286614
rect 540025 286782 540113 286798
rect 540025 286614 540041 286782
rect 540075 286614 540113 286782
rect 540025 286598 540113 286614
rect 541113 286782 541201 286798
rect 541113 286614 541151 286782
rect 541185 286614 541201 286782
rect 541113 286598 541201 286614
rect 541243 286782 541331 286798
rect 541243 286614 541259 286782
rect 541293 286614 541331 286782
rect 541243 286598 541331 286614
rect 542331 286782 542419 286798
rect 542331 286614 542369 286782
rect 542403 286614 542419 286782
rect 542331 286598 542419 286614
rect 542461 286782 542549 286798
rect 542461 286614 542477 286782
rect 542511 286614 542549 286782
rect 542461 286598 542549 286614
rect 543549 286782 543637 286798
rect 543549 286614 543587 286782
rect 543621 286614 543637 286782
rect 543549 286598 543637 286614
rect 543679 286782 543767 286798
rect 543679 286614 543695 286782
rect 543729 286614 543767 286782
rect 543679 286598 543767 286614
rect 544767 286782 544855 286798
rect 544767 286614 544805 286782
rect 544839 286614 544855 286782
rect 544767 286598 544855 286614
rect 536371 286182 536459 286198
rect 536371 286014 536387 286182
rect 536421 286014 536459 286182
rect 536371 285998 536459 286014
rect 537459 286182 537547 286198
rect 537459 286014 537497 286182
rect 537531 286014 537547 286182
rect 537459 285998 537547 286014
rect 537589 286182 537677 286198
rect 537589 286014 537605 286182
rect 537639 286014 537677 286182
rect 537589 285998 537677 286014
rect 538677 286182 538765 286198
rect 538677 286014 538715 286182
rect 538749 286014 538765 286182
rect 538677 285998 538765 286014
rect 538807 286182 538895 286198
rect 538807 286014 538823 286182
rect 538857 286014 538895 286182
rect 538807 285998 538895 286014
rect 539895 286182 539983 286198
rect 539895 286014 539933 286182
rect 539967 286014 539983 286182
rect 539895 285998 539983 286014
rect 540025 286182 540113 286198
rect 540025 286014 540041 286182
rect 540075 286014 540113 286182
rect 540025 285998 540113 286014
rect 541113 286182 541201 286198
rect 541113 286014 541151 286182
rect 541185 286014 541201 286182
rect 541113 285998 541201 286014
rect 541243 286182 541331 286198
rect 541243 286014 541259 286182
rect 541293 286014 541331 286182
rect 541243 285998 541331 286014
rect 542331 286182 542419 286198
rect 542331 286014 542369 286182
rect 542403 286014 542419 286182
rect 542331 285998 542419 286014
rect 542461 286182 542549 286198
rect 542461 286014 542477 286182
rect 542511 286014 542549 286182
rect 542461 285998 542549 286014
rect 543549 286182 543637 286198
rect 543549 286014 543587 286182
rect 543621 286014 543637 286182
rect 543549 285998 543637 286014
rect 543679 286182 543767 286198
rect 543679 286014 543695 286182
rect 543729 286014 543767 286182
rect 543679 285998 543767 286014
rect 544767 286182 544855 286198
rect 544767 286014 544805 286182
rect 544839 286014 544855 286182
rect 544767 285998 544855 286014
rect 536916 285208 537013 285224
rect 536916 285040 536932 285208
rect 536966 285040 537013 285208
rect 536916 285024 537013 285040
rect 538013 285208 538110 285224
rect 538013 285040 538060 285208
rect 538094 285040 538110 285208
rect 538013 285024 538110 285040
rect 538152 285208 538249 285224
rect 538152 285040 538168 285208
rect 538202 285040 538249 285208
rect 538152 285024 538249 285040
rect 539249 285208 539346 285224
rect 539249 285040 539296 285208
rect 539330 285040 539346 285208
rect 539249 285024 539346 285040
rect 539388 285208 539485 285224
rect 539388 285040 539404 285208
rect 539438 285040 539485 285208
rect 539388 285024 539485 285040
rect 540485 285208 540582 285224
rect 540485 285040 540532 285208
rect 540566 285040 540582 285208
rect 540485 285024 540582 285040
rect 540624 285208 540721 285224
rect 540624 285040 540640 285208
rect 540674 285040 540721 285208
rect 540624 285024 540721 285040
rect 541721 285208 541818 285224
rect 541721 285040 541768 285208
rect 541802 285040 541818 285208
rect 541721 285024 541818 285040
rect 541860 285208 541957 285224
rect 541860 285040 541876 285208
rect 541910 285040 541957 285208
rect 541860 285024 541957 285040
rect 542957 285208 543054 285224
rect 542957 285040 543004 285208
rect 543038 285040 543054 285208
rect 542957 285024 543054 285040
rect 543096 285208 543193 285224
rect 543096 285040 543112 285208
rect 543146 285040 543193 285208
rect 543096 285024 543193 285040
rect 544193 285208 544290 285224
rect 544193 285040 544240 285208
rect 544274 285040 544290 285208
rect 544193 285024 544290 285040
rect 536916 284618 537013 284634
rect 536916 284450 536932 284618
rect 536966 284450 537013 284618
rect 536916 284434 537013 284450
rect 538013 284618 538110 284634
rect 538013 284450 538060 284618
rect 538094 284450 538110 284618
rect 538013 284434 538110 284450
rect 538152 284618 538249 284634
rect 538152 284450 538168 284618
rect 538202 284450 538249 284618
rect 538152 284434 538249 284450
rect 539249 284618 539346 284634
rect 539249 284450 539296 284618
rect 539330 284450 539346 284618
rect 539249 284434 539346 284450
rect 539388 284618 539485 284634
rect 539388 284450 539404 284618
rect 539438 284450 539485 284618
rect 539388 284434 539485 284450
rect 540485 284618 540582 284634
rect 540485 284450 540532 284618
rect 540566 284450 540582 284618
rect 540485 284434 540582 284450
rect 540624 284618 540721 284634
rect 540624 284450 540640 284618
rect 540674 284450 540721 284618
rect 540624 284434 540721 284450
rect 541721 284618 541818 284634
rect 541721 284450 541768 284618
rect 541802 284450 541818 284618
rect 541721 284434 541818 284450
rect 541860 284618 541957 284634
rect 541860 284450 541876 284618
rect 541910 284450 541957 284618
rect 541860 284434 541957 284450
rect 542957 284618 543054 284634
rect 542957 284450 543004 284618
rect 543038 284450 543054 284618
rect 542957 284434 543054 284450
rect 543096 284618 543193 284634
rect 543096 284450 543112 284618
rect 543146 284450 543193 284618
rect 543096 284434 543193 284450
rect 544193 284618 544290 284634
rect 544193 284450 544240 284618
rect 544274 284450 544290 284618
rect 544193 284434 544290 284450
rect 539686 283828 539774 283844
rect 539686 283660 539702 283828
rect 539736 283660 539774 283828
rect 539686 283644 539774 283660
rect 540024 283828 540112 283844
rect 540024 283660 540062 283828
rect 540096 283660 540112 283828
rect 540024 283644 540112 283660
rect 540154 283828 540242 283844
rect 540154 283660 540170 283828
rect 540204 283660 540242 283828
rect 540154 283644 540242 283660
rect 540492 283828 540580 283844
rect 540492 283660 540530 283828
rect 540564 283660 540580 283828
rect 540492 283644 540580 283660
rect 540622 283828 540710 283844
rect 540622 283660 540638 283828
rect 540672 283660 540710 283828
rect 540622 283644 540710 283660
rect 540960 283828 541048 283844
rect 540960 283660 540998 283828
rect 541032 283660 541048 283828
rect 540960 283644 541048 283660
rect 541090 283828 541178 283844
rect 541090 283660 541106 283828
rect 541140 283660 541178 283828
rect 541090 283644 541178 283660
rect 541428 283828 541516 283844
rect 541428 283660 541466 283828
rect 541500 283660 541516 283828
rect 541428 283644 541516 283660
rect 539906 283203 539994 283219
rect 539906 283135 539922 283203
rect 539956 283135 539994 283203
rect 539906 283119 539994 283135
rect 540494 283203 540582 283219
rect 540494 283135 540532 283203
rect 540566 283135 540582 283203
rect 540494 283119 540582 283135
rect 540624 283203 540712 283219
rect 540624 283135 540640 283203
rect 540674 283135 540712 283203
rect 540624 283119 540712 283135
rect 541212 283203 541300 283219
rect 541212 283135 541250 283203
rect 541284 283135 541300 283203
rect 541212 283119 541300 283135
rect 536971 282678 537059 282694
rect 536971 282510 536987 282678
rect 537021 282510 537059 282678
rect 536971 282494 537059 282510
rect 538059 282678 538147 282694
rect 538059 282510 538097 282678
rect 538131 282510 538147 282678
rect 538059 282494 538147 282510
rect 538189 282678 538277 282694
rect 538189 282510 538205 282678
rect 538239 282510 538277 282678
rect 538189 282494 538277 282510
rect 539277 282678 539365 282694
rect 539277 282510 539315 282678
rect 539349 282510 539365 282678
rect 539277 282494 539365 282510
rect 539407 282678 539495 282694
rect 539407 282510 539423 282678
rect 539457 282510 539495 282678
rect 539407 282494 539495 282510
rect 540495 282678 540583 282694
rect 540495 282510 540533 282678
rect 540567 282510 540583 282678
rect 540495 282494 540583 282510
rect 540625 282678 540713 282694
rect 540625 282510 540641 282678
rect 540675 282510 540713 282678
rect 540625 282494 540713 282510
rect 541713 282678 541801 282694
rect 541713 282510 541751 282678
rect 541785 282510 541801 282678
rect 541713 282494 541801 282510
rect 541843 282678 541931 282694
rect 541843 282510 541859 282678
rect 541893 282510 541931 282678
rect 541843 282494 541931 282510
rect 542931 282678 543019 282694
rect 542931 282510 542969 282678
rect 543003 282510 543019 282678
rect 542931 282494 543019 282510
rect 543061 282678 543149 282694
rect 543061 282510 543077 282678
rect 543111 282510 543149 282678
rect 543061 282494 543149 282510
rect 544149 282678 544237 282694
rect 544149 282510 544187 282678
rect 544221 282510 544237 282678
rect 544149 282494 544237 282510
rect 568222 281218 568288 281231
rect 568222 281215 568310 281218
rect 568222 281181 568238 281215
rect 568272 281181 568310 281215
rect 568222 281178 568310 281181
rect 578310 281178 578336 281218
rect 568222 281165 568288 281178
rect 578332 281120 578398 281133
rect 568284 281080 568310 281120
rect 578310 281117 578398 281120
rect 578310 281083 578348 281117
rect 578382 281083 578398 281117
rect 578310 281080 578398 281083
rect 568222 281022 568288 281035
rect 578332 281067 578398 281080
rect 568222 281019 568310 281022
rect 568222 280985 568238 281019
rect 568272 280985 568310 281019
rect 568222 280982 568310 280985
rect 578310 280982 578336 281022
rect 568222 280969 568288 280982
rect 578332 280924 578398 280937
rect 568284 280884 568310 280924
rect 578310 280921 578398 280924
rect 578310 280887 578348 280921
rect 578382 280887 578398 280921
rect 578310 280884 578398 280887
rect 568222 280826 568288 280839
rect 578332 280871 578398 280884
rect 568222 280823 568310 280826
rect 568222 280789 568238 280823
rect 568272 280789 568310 280823
rect 568222 280786 568310 280789
rect 578310 280786 578336 280826
rect 568222 280773 568288 280786
rect 578332 280728 578398 280741
rect 568284 280688 568310 280728
rect 578310 280725 578398 280728
rect 578310 280691 578348 280725
rect 578382 280691 578398 280725
rect 578310 280688 578398 280691
rect 568222 280630 568288 280643
rect 578332 280675 578398 280688
rect 568222 280627 568310 280630
rect 568222 280593 568238 280627
rect 568272 280593 568310 280627
rect 568222 280590 568310 280593
rect 578310 280590 578336 280630
rect 568222 280577 568288 280590
rect 578332 280532 578398 280545
rect 568284 280492 568310 280532
rect 578310 280529 578398 280532
rect 578310 280495 578348 280529
rect 578382 280495 578398 280529
rect 578310 280492 578398 280495
rect 568222 280434 568288 280447
rect 578332 280479 578398 280492
rect 568222 280431 568310 280434
rect 568222 280397 568238 280431
rect 568272 280397 568310 280431
rect 568222 280394 568310 280397
rect 578310 280394 578336 280434
rect 568222 280381 568288 280394
rect 578332 280336 578398 280349
rect 568284 280296 568310 280336
rect 578310 280333 578398 280336
rect 578310 280299 578348 280333
rect 578382 280299 578398 280333
rect 578310 280296 578398 280299
rect 578332 280283 578398 280296
rect 12704 275772 12801 275788
rect 12704 275704 12720 275772
rect 12754 275704 12801 275772
rect 12704 275688 12801 275704
rect 13801 275772 13898 275788
rect 13801 275704 13848 275772
rect 13882 275704 13898 275772
rect 13801 275688 13898 275704
rect 12704 275614 12801 275630
rect 12704 275546 12720 275614
rect 12754 275546 12801 275614
rect 12704 275530 12801 275546
rect 13801 275614 13898 275630
rect 13801 275546 13848 275614
rect 13882 275546 13898 275614
rect 13801 275530 13898 275546
rect 12704 275456 12801 275472
rect 12704 275388 12720 275456
rect 12754 275388 12801 275456
rect 12704 275372 12801 275388
rect 13801 275456 13898 275472
rect 13801 275388 13848 275456
rect 13882 275388 13898 275456
rect 13801 275372 13898 275388
rect 12704 275298 12801 275314
rect 12704 275230 12720 275298
rect 12754 275230 12801 275298
rect 12704 275214 12801 275230
rect 13801 275298 13898 275314
rect 13801 275230 13848 275298
rect 13882 275230 13898 275298
rect 13801 275214 13898 275230
rect 12704 275140 12801 275156
rect 12704 275072 12720 275140
rect 12754 275072 12801 275140
rect 12704 275056 12801 275072
rect 13801 275140 13898 275156
rect 13801 275072 13848 275140
rect 13882 275072 13898 275140
rect 13801 275056 13898 275072
rect 12704 274982 12801 274998
rect 12704 274914 12720 274982
rect 12754 274914 12801 274982
rect 12704 274898 12801 274914
rect 13801 274982 13898 274998
rect 13801 274914 13848 274982
rect 13882 274914 13898 274982
rect 13801 274898 13898 274914
rect 12704 274824 12801 274840
rect 12704 274756 12720 274824
rect 12754 274756 12801 274824
rect 12704 274740 12801 274756
rect 13801 274824 13898 274840
rect 13801 274756 13848 274824
rect 13882 274756 13898 274824
rect 13801 274740 13898 274756
rect 12704 274666 12801 274682
rect 12704 274598 12720 274666
rect 12754 274598 12801 274666
rect 12704 274582 12801 274598
rect 13801 274666 13898 274682
rect 13801 274598 13848 274666
rect 13882 274598 13898 274666
rect 13801 274582 13898 274598
rect 12704 274508 12801 274524
rect 12704 274440 12720 274508
rect 12754 274440 12801 274508
rect 12704 274424 12801 274440
rect 13801 274508 13898 274524
rect 13801 274440 13848 274508
rect 13882 274440 13898 274508
rect 13801 274424 13898 274440
rect 12704 274350 12801 274366
rect 12704 274282 12720 274350
rect 12754 274282 12801 274350
rect 12704 274266 12801 274282
rect 13801 274350 13898 274366
rect 13801 274282 13848 274350
rect 13882 274282 13898 274350
rect 13801 274266 13898 274282
rect 12704 274192 12801 274208
rect 12704 274124 12720 274192
rect 12754 274124 12801 274192
rect 12704 274108 12801 274124
rect 13801 274192 13898 274208
rect 13801 274124 13848 274192
rect 13882 274124 13898 274192
rect 13801 274108 13898 274124
rect 12704 274034 12801 274050
rect 12704 273966 12720 274034
rect 12754 273966 12801 274034
rect 12704 273950 12801 273966
rect 13801 274034 13898 274050
rect 13801 273966 13848 274034
rect 13882 273966 13898 274034
rect 13801 273950 13898 273966
rect 12704 273876 12801 273892
rect 12704 273808 12720 273876
rect 12754 273808 12801 273876
rect 12704 273792 12801 273808
rect 13801 273876 13898 273892
rect 13801 273808 13848 273876
rect 13882 273808 13898 273876
rect 13801 273792 13898 273808
rect 12704 273718 12801 273734
rect 12704 273650 12720 273718
rect 12754 273650 12801 273718
rect 12704 273634 12801 273650
rect 13801 273718 13898 273734
rect 13801 273650 13848 273718
rect 13882 273650 13898 273718
rect 13801 273634 13898 273650
rect 12704 273560 12801 273576
rect 12704 273492 12720 273560
rect 12754 273492 12801 273560
rect 12704 273476 12801 273492
rect 13801 273560 13898 273576
rect 13801 273492 13848 273560
rect 13882 273492 13898 273560
rect 13801 273476 13898 273492
rect 12704 273402 12801 273418
rect 12704 273334 12720 273402
rect 12754 273334 12801 273402
rect 12704 273318 12801 273334
rect 13801 273402 13898 273418
rect 13801 273334 13848 273402
rect 13882 273334 13898 273402
rect 13801 273318 13898 273334
rect 12704 273244 12801 273260
rect 12704 273176 12720 273244
rect 12754 273176 12801 273244
rect 12704 273160 12801 273176
rect 13801 273244 13898 273260
rect 13801 273176 13848 273244
rect 13882 273176 13898 273244
rect 13801 273160 13898 273176
rect 12704 273086 12801 273102
rect 12704 273018 12720 273086
rect 12754 273018 12801 273086
rect 12704 273002 12801 273018
rect 13801 273086 13898 273102
rect 13801 273018 13848 273086
rect 13882 273018 13898 273086
rect 13801 273002 13898 273018
rect 12704 272928 12801 272944
rect 12704 272860 12720 272928
rect 12754 272860 12801 272928
rect 12704 272844 12801 272860
rect 13801 272928 13898 272944
rect 13801 272860 13848 272928
rect 13882 272860 13898 272928
rect 13801 272844 13898 272860
rect 12704 272770 12801 272786
rect 12704 272702 12720 272770
rect 12754 272702 12801 272770
rect 12704 272686 12801 272702
rect 13801 272770 13898 272786
rect 13801 272702 13848 272770
rect 13882 272702 13898 272770
rect 13801 272686 13898 272702
rect 12704 272612 12801 272628
rect 12704 272544 12720 272612
rect 12754 272544 12801 272612
rect 12704 272528 12801 272544
rect 13801 272612 13898 272628
rect 13801 272544 13848 272612
rect 13882 272544 13898 272612
rect 13801 272528 13898 272544
rect 12704 272454 12801 272470
rect 12704 272386 12720 272454
rect 12754 272386 12801 272454
rect 12704 272370 12801 272386
rect 13801 272454 13898 272470
rect 13801 272386 13848 272454
rect 13882 272386 13898 272454
rect 13801 272370 13898 272386
rect 12704 272296 12801 272312
rect 12704 272228 12720 272296
rect 12754 272228 12801 272296
rect 12704 272212 12801 272228
rect 13801 272296 13898 272312
rect 13801 272228 13848 272296
rect 13882 272228 13898 272296
rect 13801 272212 13898 272228
rect 12704 272138 12801 272154
rect 12704 272070 12720 272138
rect 12754 272070 12801 272138
rect 12704 272054 12801 272070
rect 13801 272138 13898 272154
rect 13801 272070 13848 272138
rect 13882 272070 13898 272138
rect 13801 272054 13898 272070
rect 12704 271980 12801 271996
rect 12704 271912 12720 271980
rect 12754 271912 12801 271980
rect 12704 271896 12801 271912
rect 13801 271980 13898 271996
rect 13801 271912 13848 271980
rect 13882 271912 13898 271980
rect 13801 271896 13898 271912
rect 12704 271822 12801 271838
rect 12704 271754 12720 271822
rect 12754 271754 12801 271822
rect 12704 271738 12801 271754
rect 13801 271822 13898 271838
rect 13801 271754 13848 271822
rect 13882 271754 13898 271822
rect 13801 271738 13898 271754
rect 12704 271664 12801 271680
rect 12704 271596 12720 271664
rect 12754 271596 12801 271664
rect 12704 271580 12801 271596
rect 13801 271664 13898 271680
rect 13801 271596 13848 271664
rect 13882 271596 13898 271664
rect 13801 271580 13898 271596
rect 12704 271506 12801 271522
rect 12704 271438 12720 271506
rect 12754 271438 12801 271506
rect 12704 271422 12801 271438
rect 13801 271506 13898 271522
rect 13801 271438 13848 271506
rect 13882 271438 13898 271506
rect 13801 271422 13898 271438
rect 12704 271348 12801 271364
rect 12704 271280 12720 271348
rect 12754 271280 12801 271348
rect 12704 271264 12801 271280
rect 13801 271348 13898 271364
rect 13801 271280 13848 271348
rect 13882 271280 13898 271348
rect 13801 271264 13898 271280
rect 12704 271190 12801 271206
rect 12704 271122 12720 271190
rect 12754 271122 12801 271190
rect 12704 271106 12801 271122
rect 13801 271190 13898 271206
rect 13801 271122 13848 271190
rect 13882 271122 13898 271190
rect 13801 271106 13898 271122
rect 12704 271032 12801 271048
rect 12704 270964 12720 271032
rect 12754 270964 12801 271032
rect 12704 270948 12801 270964
rect 13801 271032 13898 271048
rect 13801 270964 13848 271032
rect 13882 270964 13898 271032
rect 13801 270948 13898 270964
rect 12704 270874 12801 270890
rect 12704 270806 12720 270874
rect 12754 270806 12801 270874
rect 12704 270790 12801 270806
rect 13801 270874 13898 270890
rect 13801 270806 13848 270874
rect 13882 270806 13898 270874
rect 13801 270790 13898 270806
rect 12704 270716 12801 270732
rect 12704 270648 12720 270716
rect 12754 270648 12801 270716
rect 12704 270632 12801 270648
rect 13801 270716 13898 270732
rect 13801 270648 13848 270716
rect 13882 270648 13898 270716
rect 13801 270632 13898 270648
rect 12704 270558 12801 270574
rect 12704 270490 12720 270558
rect 12754 270490 12801 270558
rect 12704 270474 12801 270490
rect 13801 270558 13898 270574
rect 13801 270490 13848 270558
rect 13882 270490 13898 270558
rect 13801 270474 13898 270490
rect 12704 270400 12801 270416
rect 12704 270332 12720 270400
rect 12754 270332 12801 270400
rect 12704 270316 12801 270332
rect 13801 270400 13898 270416
rect 13801 270332 13848 270400
rect 13882 270332 13898 270400
rect 13801 270316 13898 270332
rect 12704 270242 12801 270258
rect 12704 270174 12720 270242
rect 12754 270174 12801 270242
rect 12704 270158 12801 270174
rect 13801 270242 13898 270258
rect 13801 270174 13848 270242
rect 13882 270174 13898 270242
rect 13801 270158 13898 270174
rect 12704 270084 12801 270100
rect 12704 270016 12720 270084
rect 12754 270016 12801 270084
rect 12704 270000 12801 270016
rect 13801 270084 13898 270100
rect 13801 270016 13848 270084
rect 13882 270016 13898 270084
rect 13801 270000 13898 270016
rect 12704 269926 12801 269942
rect 12704 269858 12720 269926
rect 12754 269858 12801 269926
rect 12704 269842 12801 269858
rect 13801 269926 13898 269942
rect 13801 269858 13848 269926
rect 13882 269858 13898 269926
rect 13801 269842 13898 269858
rect 12704 269768 12801 269784
rect 12704 269700 12720 269768
rect 12754 269700 12801 269768
rect 12704 269684 12801 269700
rect 13801 269768 13898 269784
rect 13801 269700 13848 269768
rect 13882 269700 13898 269768
rect 13801 269684 13898 269700
rect 12704 269610 12801 269626
rect 12704 269542 12720 269610
rect 12754 269542 12801 269610
rect 12704 269526 12801 269542
rect 13801 269610 13898 269626
rect 13801 269542 13848 269610
rect 13882 269542 13898 269610
rect 13801 269526 13898 269542
rect 14374 274270 14471 274286
rect 14374 274202 14390 274270
rect 14424 274202 14471 274270
rect 14374 274186 14471 274202
rect 15471 274270 15568 274286
rect 15471 274202 15518 274270
rect 15552 274202 15568 274270
rect 15471 274186 15568 274202
rect 14374 274112 14471 274128
rect 14374 274044 14390 274112
rect 14424 274044 14471 274112
rect 14374 274028 14471 274044
rect 15471 274112 15568 274128
rect 15471 274044 15518 274112
rect 15552 274044 15568 274112
rect 15471 274028 15568 274044
rect 14374 273954 14471 273970
rect 14374 273886 14390 273954
rect 14424 273886 14471 273954
rect 14374 273870 14471 273886
rect 15471 273954 15568 273970
rect 15471 273886 15518 273954
rect 15552 273886 15568 273954
rect 15471 273870 15568 273886
rect 14374 273796 14471 273812
rect 14374 273728 14390 273796
rect 14424 273728 14471 273796
rect 14374 273712 14471 273728
rect 15471 273796 15568 273812
rect 15471 273728 15518 273796
rect 15552 273728 15568 273796
rect 15471 273712 15568 273728
rect 14374 273638 14471 273654
rect 14374 273570 14390 273638
rect 14424 273570 14471 273638
rect 14374 273554 14471 273570
rect 15471 273638 15568 273654
rect 15471 273570 15518 273638
rect 15552 273570 15568 273638
rect 15471 273554 15568 273570
rect 14374 273480 14471 273496
rect 14374 273412 14390 273480
rect 14424 273412 14471 273480
rect 14374 273396 14471 273412
rect 15471 273480 15568 273496
rect 15471 273412 15518 273480
rect 15552 273412 15568 273480
rect 15471 273396 15568 273412
rect 14374 273322 14471 273338
rect 14374 273254 14390 273322
rect 14424 273254 14471 273322
rect 14374 273238 14471 273254
rect 15471 273322 15568 273338
rect 15471 273254 15518 273322
rect 15552 273254 15568 273322
rect 15471 273238 15568 273254
rect 14374 273164 14471 273180
rect 14374 273096 14390 273164
rect 14424 273096 14471 273164
rect 14374 273080 14471 273096
rect 15471 273164 15568 273180
rect 15471 273096 15518 273164
rect 15552 273096 15568 273164
rect 15471 273080 15568 273096
rect 14374 273006 14471 273022
rect 14374 272938 14390 273006
rect 14424 272938 14471 273006
rect 14374 272922 14471 272938
rect 15471 273006 15568 273022
rect 15471 272938 15518 273006
rect 15552 272938 15568 273006
rect 15471 272922 15568 272938
rect 14374 272848 14471 272864
rect 14374 272780 14390 272848
rect 14424 272780 14471 272848
rect 14374 272764 14471 272780
rect 15471 272848 15568 272864
rect 15471 272780 15518 272848
rect 15552 272780 15568 272848
rect 15471 272764 15568 272780
rect 14374 272690 14471 272706
rect 14374 272622 14390 272690
rect 14424 272622 14471 272690
rect 14374 272606 14471 272622
rect 15471 272690 15568 272706
rect 15471 272622 15518 272690
rect 15552 272622 15568 272690
rect 15471 272606 15568 272622
rect 14374 272532 14471 272548
rect 14374 272464 14390 272532
rect 14424 272464 14471 272532
rect 14374 272448 14471 272464
rect 15471 272532 15568 272548
rect 15471 272464 15518 272532
rect 15552 272464 15568 272532
rect 15471 272448 15568 272464
rect 14374 272374 14471 272390
rect 14374 272306 14390 272374
rect 14424 272306 14471 272374
rect 14374 272290 14471 272306
rect 15471 272374 15568 272390
rect 15471 272306 15518 272374
rect 15552 272306 15568 272374
rect 15471 272290 15568 272306
rect 14374 272216 14471 272232
rect 14374 272148 14390 272216
rect 14424 272148 14471 272216
rect 14374 272132 14471 272148
rect 15471 272216 15568 272232
rect 15471 272148 15518 272216
rect 15552 272148 15568 272216
rect 15471 272132 15568 272148
rect 14374 272058 14471 272074
rect 14374 271990 14390 272058
rect 14424 271990 14471 272058
rect 14374 271974 14471 271990
rect 15471 272058 15568 272074
rect 15471 271990 15518 272058
rect 15552 271990 15568 272058
rect 15471 271974 15568 271990
rect 14374 271900 14471 271916
rect 14374 271832 14390 271900
rect 14424 271832 14471 271900
rect 14374 271816 14471 271832
rect 15471 271900 15568 271916
rect 15471 271832 15518 271900
rect 15552 271832 15568 271900
rect 15471 271816 15568 271832
rect 14374 271742 14471 271758
rect 14374 271674 14390 271742
rect 14424 271674 14471 271742
rect 14374 271658 14471 271674
rect 15471 271742 15568 271758
rect 15471 271674 15518 271742
rect 15552 271674 15568 271742
rect 15471 271658 15568 271674
rect 14374 271584 14471 271600
rect 14374 271516 14390 271584
rect 14424 271516 14471 271584
rect 14374 271500 14471 271516
rect 15471 271584 15568 271600
rect 15471 271516 15518 271584
rect 15552 271516 15568 271584
rect 15471 271500 15568 271516
rect 14374 271426 14471 271442
rect 14374 271358 14390 271426
rect 14424 271358 14471 271426
rect 14374 271342 14471 271358
rect 15471 271426 15568 271442
rect 15471 271358 15518 271426
rect 15552 271358 15568 271426
rect 15471 271342 15568 271358
rect 14374 271268 14471 271284
rect 14374 271200 14390 271268
rect 14424 271200 14471 271268
rect 14374 271184 14471 271200
rect 15471 271268 15568 271284
rect 15471 271200 15518 271268
rect 15552 271200 15568 271268
rect 15471 271184 15568 271200
rect 14374 271110 14471 271126
rect 14374 271042 14390 271110
rect 14424 271042 14471 271110
rect 14374 271026 14471 271042
rect 15471 271110 15568 271126
rect 15471 271042 15518 271110
rect 15552 271042 15568 271110
rect 15471 271026 15568 271042
rect 15914 274270 16011 274286
rect 15914 274202 15930 274270
rect 15964 274202 16011 274270
rect 15914 274186 16011 274202
rect 17011 274270 17108 274286
rect 17011 274202 17058 274270
rect 17092 274202 17108 274270
rect 17011 274186 17108 274202
rect 15914 274112 16011 274128
rect 15914 274044 15930 274112
rect 15964 274044 16011 274112
rect 15914 274028 16011 274044
rect 17011 274112 17108 274128
rect 17011 274044 17058 274112
rect 17092 274044 17108 274112
rect 17011 274028 17108 274044
rect 15914 273954 16011 273970
rect 15914 273886 15930 273954
rect 15964 273886 16011 273954
rect 15914 273870 16011 273886
rect 17011 273954 17108 273970
rect 17011 273886 17058 273954
rect 17092 273886 17108 273954
rect 17011 273870 17108 273886
rect 15914 273796 16011 273812
rect 15914 273728 15930 273796
rect 15964 273728 16011 273796
rect 15914 273712 16011 273728
rect 17011 273796 17108 273812
rect 17011 273728 17058 273796
rect 17092 273728 17108 273796
rect 17011 273712 17108 273728
rect 15914 273638 16011 273654
rect 15914 273570 15930 273638
rect 15964 273570 16011 273638
rect 15914 273554 16011 273570
rect 17011 273638 17108 273654
rect 17011 273570 17058 273638
rect 17092 273570 17108 273638
rect 17011 273554 17108 273570
rect 15914 273480 16011 273496
rect 15914 273412 15930 273480
rect 15964 273412 16011 273480
rect 15914 273396 16011 273412
rect 17011 273480 17108 273496
rect 17011 273412 17058 273480
rect 17092 273412 17108 273480
rect 17011 273396 17108 273412
rect 15914 273322 16011 273338
rect 15914 273254 15930 273322
rect 15964 273254 16011 273322
rect 15914 273238 16011 273254
rect 17011 273322 17108 273338
rect 17011 273254 17058 273322
rect 17092 273254 17108 273322
rect 17011 273238 17108 273254
rect 15914 273164 16011 273180
rect 15914 273096 15930 273164
rect 15964 273096 16011 273164
rect 15914 273080 16011 273096
rect 17011 273164 17108 273180
rect 17011 273096 17058 273164
rect 17092 273096 17108 273164
rect 17011 273080 17108 273096
rect 15914 273006 16011 273022
rect 15914 272938 15930 273006
rect 15964 272938 16011 273006
rect 15914 272922 16011 272938
rect 17011 273006 17108 273022
rect 17011 272938 17058 273006
rect 17092 272938 17108 273006
rect 17011 272922 17108 272938
rect 15914 272848 16011 272864
rect 15914 272780 15930 272848
rect 15964 272780 16011 272848
rect 15914 272764 16011 272780
rect 17011 272848 17108 272864
rect 17011 272780 17058 272848
rect 17092 272780 17108 272848
rect 17011 272764 17108 272780
rect 15914 272690 16011 272706
rect 15914 272622 15930 272690
rect 15964 272622 16011 272690
rect 15914 272606 16011 272622
rect 17011 272690 17108 272706
rect 17011 272622 17058 272690
rect 17092 272622 17108 272690
rect 17011 272606 17108 272622
rect 15914 272532 16011 272548
rect 15914 272464 15930 272532
rect 15964 272464 16011 272532
rect 15914 272448 16011 272464
rect 17011 272532 17108 272548
rect 17011 272464 17058 272532
rect 17092 272464 17108 272532
rect 17011 272448 17108 272464
rect 15914 272374 16011 272390
rect 15914 272306 15930 272374
rect 15964 272306 16011 272374
rect 15914 272290 16011 272306
rect 17011 272374 17108 272390
rect 17011 272306 17058 272374
rect 17092 272306 17108 272374
rect 17011 272290 17108 272306
rect 15914 272216 16011 272232
rect 15914 272148 15930 272216
rect 15964 272148 16011 272216
rect 15914 272132 16011 272148
rect 17011 272216 17108 272232
rect 17011 272148 17058 272216
rect 17092 272148 17108 272216
rect 17011 272132 17108 272148
rect 15914 272058 16011 272074
rect 15914 271990 15930 272058
rect 15964 271990 16011 272058
rect 15914 271974 16011 271990
rect 17011 272058 17108 272074
rect 17011 271990 17058 272058
rect 17092 271990 17108 272058
rect 17011 271974 17108 271990
rect 15914 271900 16011 271916
rect 15914 271832 15930 271900
rect 15964 271832 16011 271900
rect 15914 271816 16011 271832
rect 17011 271900 17108 271916
rect 17011 271832 17058 271900
rect 17092 271832 17108 271900
rect 17011 271816 17108 271832
rect 15914 271742 16011 271758
rect 15914 271674 15930 271742
rect 15964 271674 16011 271742
rect 15914 271658 16011 271674
rect 17011 271742 17108 271758
rect 17011 271674 17058 271742
rect 17092 271674 17108 271742
rect 17011 271658 17108 271674
rect 15914 271584 16011 271600
rect 15914 271516 15930 271584
rect 15964 271516 16011 271584
rect 15914 271500 16011 271516
rect 17011 271584 17108 271600
rect 17011 271516 17058 271584
rect 17092 271516 17108 271584
rect 17011 271500 17108 271516
rect 15914 271426 16011 271442
rect 15914 271358 15930 271426
rect 15964 271358 16011 271426
rect 15914 271342 16011 271358
rect 17011 271426 17108 271442
rect 17011 271358 17058 271426
rect 17092 271358 17108 271426
rect 17011 271342 17108 271358
rect 15914 271268 16011 271284
rect 15914 271200 15930 271268
rect 15964 271200 16011 271268
rect 15914 271184 16011 271200
rect 17011 271268 17108 271284
rect 17011 271200 17058 271268
rect 17092 271200 17108 271268
rect 17011 271184 17108 271200
rect 15914 271110 16011 271126
rect 15914 271042 15930 271110
rect 15964 271042 16011 271110
rect 15914 271026 16011 271042
rect 17011 271110 17108 271126
rect 17011 271042 17058 271110
rect 17092 271042 17108 271110
rect 17011 271026 17108 271042
rect 17491 273159 17579 273175
rect 17491 273091 17507 273159
rect 17541 273091 17579 273159
rect 17491 273075 17579 273091
rect 18579 273159 18667 273175
rect 18579 273091 18617 273159
rect 18651 273091 18667 273159
rect 18579 273075 18667 273091
rect 17491 273001 17579 273017
rect 17491 272933 17507 273001
rect 17541 272933 17579 273001
rect 17491 272917 17579 272933
rect 18579 273001 18667 273017
rect 18579 272933 18617 273001
rect 18651 272933 18667 273001
rect 18579 272917 18667 272933
rect 17491 272843 17579 272859
rect 17491 272775 17507 272843
rect 17541 272775 17579 272843
rect 17491 272759 17579 272775
rect 18579 272843 18667 272859
rect 18579 272775 18617 272843
rect 18651 272775 18667 272843
rect 18579 272759 18667 272775
rect 17491 272685 17579 272701
rect 17491 272617 17507 272685
rect 17541 272617 17579 272685
rect 17491 272601 17579 272617
rect 18579 272685 18667 272701
rect 18579 272617 18617 272685
rect 18651 272617 18667 272685
rect 18579 272601 18667 272617
rect 17491 272527 17579 272543
rect 17491 272459 17507 272527
rect 17541 272459 17579 272527
rect 17491 272443 17579 272459
rect 18579 272527 18667 272543
rect 18579 272459 18617 272527
rect 18651 272459 18667 272527
rect 18579 272443 18667 272459
rect 17491 272369 17579 272385
rect 17491 272301 17507 272369
rect 17541 272301 17579 272369
rect 17491 272285 17579 272301
rect 18579 272369 18667 272385
rect 18579 272301 18617 272369
rect 18651 272301 18667 272369
rect 18579 272285 18667 272301
rect 17491 272211 17579 272227
rect 17491 272143 17507 272211
rect 17541 272143 17579 272211
rect 17491 272127 17579 272143
rect 18579 272211 18667 272227
rect 18579 272143 18617 272211
rect 18651 272143 18667 272211
rect 18579 272127 18667 272143
rect 19011 273159 19099 273175
rect 19011 273091 19027 273159
rect 19061 273091 19099 273159
rect 19011 273075 19099 273091
rect 20099 273159 20187 273175
rect 20099 273091 20137 273159
rect 20171 273091 20187 273159
rect 20099 273075 20187 273091
rect 19011 273001 19099 273017
rect 19011 272933 19027 273001
rect 19061 272933 19099 273001
rect 19011 272917 19099 272933
rect 20099 273001 20187 273017
rect 20099 272933 20137 273001
rect 20171 272933 20187 273001
rect 20099 272917 20187 272933
rect 19011 272843 19099 272859
rect 19011 272775 19027 272843
rect 19061 272775 19099 272843
rect 19011 272759 19099 272775
rect 20099 272843 20187 272859
rect 20099 272775 20137 272843
rect 20171 272775 20187 272843
rect 20099 272759 20187 272775
rect 19011 272685 19099 272701
rect 19011 272617 19027 272685
rect 19061 272617 19099 272685
rect 19011 272601 19099 272617
rect 20099 272685 20187 272701
rect 20099 272617 20137 272685
rect 20171 272617 20187 272685
rect 20099 272601 20187 272617
rect 19011 272527 19099 272543
rect 19011 272459 19027 272527
rect 19061 272459 19099 272527
rect 19011 272443 19099 272459
rect 20099 272527 20187 272543
rect 20099 272459 20137 272527
rect 20171 272459 20187 272527
rect 20099 272443 20187 272459
rect 19011 272369 19099 272385
rect 19011 272301 19027 272369
rect 19061 272301 19099 272369
rect 19011 272285 19099 272301
rect 20099 272369 20187 272385
rect 20099 272301 20137 272369
rect 20171 272301 20187 272369
rect 20099 272285 20187 272301
rect 19011 272211 19099 272227
rect 19011 272143 19027 272211
rect 19061 272143 19099 272211
rect 19011 272127 19099 272143
rect 20099 272211 20187 272227
rect 20099 272143 20137 272211
rect 20171 272143 20187 272211
rect 20099 272127 20187 272143
rect 20532 274158 20620 274174
rect 20532 273990 20548 274158
rect 20582 273990 20620 274158
rect 20532 273974 20620 273990
rect 21620 274158 21708 274174
rect 21620 273990 21658 274158
rect 21692 273990 21708 274158
rect 21620 273974 21708 273990
rect 20532 273900 20620 273916
rect 20532 273732 20548 273900
rect 20582 273732 20620 273900
rect 20532 273716 20620 273732
rect 21620 273900 21708 273916
rect 21620 273732 21658 273900
rect 21692 273732 21708 273900
rect 21620 273716 21708 273732
rect 20532 273642 20620 273658
rect 20532 273474 20548 273642
rect 20582 273474 20620 273642
rect 20532 273458 20620 273474
rect 21620 273642 21708 273658
rect 21620 273474 21658 273642
rect 21692 273474 21708 273642
rect 21620 273458 21708 273474
rect 20532 273384 20620 273400
rect 20532 273216 20548 273384
rect 20582 273216 20620 273384
rect 20532 273200 20620 273216
rect 21620 273384 21708 273400
rect 21620 273216 21658 273384
rect 21692 273216 21708 273384
rect 21620 273200 21708 273216
rect 20532 273126 20620 273142
rect 20532 272958 20548 273126
rect 20582 272958 20620 273126
rect 20532 272942 20620 272958
rect 21620 273126 21708 273142
rect 21620 272958 21658 273126
rect 21692 272958 21708 273126
rect 21620 272942 21708 272958
rect 20532 272868 20620 272884
rect 20532 272700 20548 272868
rect 20582 272700 20620 272868
rect 20532 272684 20620 272700
rect 21620 272868 21708 272884
rect 21620 272700 21658 272868
rect 21692 272700 21708 272868
rect 21620 272684 21708 272700
rect 20532 272610 20620 272626
rect 20532 272442 20548 272610
rect 20582 272442 20620 272610
rect 20532 272426 20620 272442
rect 21620 272610 21708 272626
rect 21620 272442 21658 272610
rect 21692 272442 21708 272610
rect 21620 272426 21708 272442
rect 20532 272352 20620 272368
rect 20532 272184 20548 272352
rect 20582 272184 20620 272352
rect 20532 272168 20620 272184
rect 21620 272352 21708 272368
rect 21620 272184 21658 272352
rect 21692 272184 21708 272352
rect 21620 272168 21708 272184
rect 20532 272094 20620 272110
rect 20532 271926 20548 272094
rect 20582 271926 20620 272094
rect 20532 271910 20620 271926
rect 21620 272094 21708 272110
rect 21620 271926 21658 272094
rect 21692 271926 21708 272094
rect 21620 271910 21708 271926
rect 20532 271836 20620 271852
rect 20532 271668 20548 271836
rect 20582 271668 20620 271836
rect 20532 271652 20620 271668
rect 21620 271836 21708 271852
rect 21620 271668 21658 271836
rect 21692 271668 21708 271836
rect 21620 271652 21708 271668
rect 20532 271578 20620 271594
rect 20532 271410 20548 271578
rect 20582 271410 20620 271578
rect 20532 271394 20620 271410
rect 21620 271578 21708 271594
rect 21620 271410 21658 271578
rect 21692 271410 21708 271578
rect 21620 271394 21708 271410
rect 20532 271320 20620 271336
rect 20532 271152 20548 271320
rect 20582 271152 20620 271320
rect 20532 271136 20620 271152
rect 21620 271320 21708 271336
rect 21620 271152 21658 271320
rect 21692 271152 21708 271320
rect 21620 271136 21708 271152
rect 22052 274414 22140 274430
rect 22052 274246 22068 274414
rect 22102 274246 22140 274414
rect 22052 274230 22140 274246
rect 23140 274414 23228 274430
rect 23140 274246 23178 274414
rect 23212 274246 23228 274414
rect 23140 274230 23228 274246
rect 22052 274156 22140 274172
rect 22052 273988 22068 274156
rect 22102 273988 22140 274156
rect 22052 273972 22140 273988
rect 23140 274156 23228 274172
rect 23140 273988 23178 274156
rect 23212 273988 23228 274156
rect 23140 273972 23228 273988
rect 22052 273898 22140 273914
rect 22052 273730 22068 273898
rect 22102 273730 22140 273898
rect 22052 273714 22140 273730
rect 23140 273898 23228 273914
rect 23140 273730 23178 273898
rect 23212 273730 23228 273898
rect 23140 273714 23228 273730
rect 22052 273640 22140 273656
rect 22052 273472 22068 273640
rect 22102 273472 22140 273640
rect 22052 273456 22140 273472
rect 23140 273640 23228 273656
rect 23140 273472 23178 273640
rect 23212 273472 23228 273640
rect 23140 273456 23228 273472
rect 22052 273382 22140 273398
rect 22052 273214 22068 273382
rect 22102 273214 22140 273382
rect 22052 273198 22140 273214
rect 23140 273382 23228 273398
rect 23140 273214 23178 273382
rect 23212 273214 23228 273382
rect 23140 273198 23228 273214
rect 22052 273124 22140 273140
rect 22052 272956 22068 273124
rect 22102 272956 22140 273124
rect 22052 272940 22140 272956
rect 23140 273124 23228 273140
rect 23140 272956 23178 273124
rect 23212 272956 23228 273124
rect 23140 272940 23228 272956
rect 22052 272866 22140 272882
rect 22052 272698 22068 272866
rect 22102 272698 22140 272866
rect 22052 272682 22140 272698
rect 23140 272866 23228 272882
rect 23140 272698 23178 272866
rect 23212 272698 23228 272866
rect 23140 272682 23228 272698
rect 22052 272608 22140 272624
rect 22052 272440 22068 272608
rect 22102 272440 22140 272608
rect 22052 272424 22140 272440
rect 23140 272608 23228 272624
rect 23140 272440 23178 272608
rect 23212 272440 23228 272608
rect 23140 272424 23228 272440
rect 22052 272350 22140 272366
rect 22052 272182 22068 272350
rect 22102 272182 22140 272350
rect 22052 272166 22140 272182
rect 23140 272350 23228 272366
rect 23140 272182 23178 272350
rect 23212 272182 23228 272350
rect 23140 272166 23228 272182
rect 22052 272092 22140 272108
rect 22052 271924 22068 272092
rect 22102 271924 22140 272092
rect 22052 271908 22140 271924
rect 23140 272092 23228 272108
rect 23140 271924 23178 272092
rect 23212 271924 23228 272092
rect 23140 271908 23228 271924
rect 22052 271834 22140 271850
rect 22052 271666 22068 271834
rect 22102 271666 22140 271834
rect 22052 271650 22140 271666
rect 23140 271834 23228 271850
rect 23140 271666 23178 271834
rect 23212 271666 23228 271834
rect 23140 271650 23228 271666
rect 22052 271576 22140 271592
rect 22052 271408 22068 271576
rect 22102 271408 22140 271576
rect 22052 271392 22140 271408
rect 23140 271576 23228 271592
rect 23140 271408 23178 271576
rect 23212 271408 23228 271576
rect 23140 271392 23228 271408
rect 22052 271318 22140 271334
rect 22052 271150 22068 271318
rect 22102 271150 22140 271318
rect 22052 271134 22140 271150
rect 23140 271318 23228 271334
rect 23140 271150 23178 271318
rect 23212 271150 23228 271318
rect 23140 271134 23228 271150
rect 22052 271060 22140 271076
rect 22052 270892 22068 271060
rect 22102 270892 22140 271060
rect 22052 270876 22140 270892
rect 23140 271060 23228 271076
rect 23140 270892 23178 271060
rect 23212 270892 23228 271060
rect 23140 270876 23228 270892
rect 24084 273380 24181 273396
rect 24084 273212 24100 273380
rect 24134 273212 24181 273380
rect 24084 273196 24181 273212
rect 25181 273380 25278 273396
rect 25181 273212 25228 273380
rect 25262 273212 25278 273380
rect 25181 273196 25278 273212
rect 24084 273122 24181 273138
rect 24084 272954 24100 273122
rect 24134 272954 24181 273122
rect 24084 272938 24181 272954
rect 25181 273122 25278 273138
rect 25181 272954 25228 273122
rect 25262 272954 25278 273122
rect 25181 272938 25278 272954
rect 24084 272864 24181 272880
rect 24084 272696 24100 272864
rect 24134 272696 24181 272864
rect 24084 272680 24181 272696
rect 25181 272864 25278 272880
rect 25181 272696 25228 272864
rect 25262 272696 25278 272864
rect 25181 272680 25278 272696
rect 24084 272606 24181 272622
rect 24084 272438 24100 272606
rect 24134 272438 24181 272606
rect 24084 272422 24181 272438
rect 25181 272606 25278 272622
rect 25181 272438 25228 272606
rect 25262 272438 25278 272606
rect 25181 272422 25278 272438
rect 24084 272348 24181 272364
rect 24084 272180 24100 272348
rect 24134 272180 24181 272348
rect 24084 272164 24181 272180
rect 25181 272348 25278 272364
rect 25181 272180 25228 272348
rect 25262 272180 25278 272348
rect 25181 272164 25278 272180
rect 24084 272090 24181 272106
rect 24084 271922 24100 272090
rect 24134 271922 24181 272090
rect 24084 271906 24181 271922
rect 25181 272090 25278 272106
rect 25181 271922 25228 272090
rect 25262 271922 25278 272090
rect 25181 271906 25278 271922
rect 25584 273380 25681 273396
rect 25584 273212 25600 273380
rect 25634 273212 25681 273380
rect 25584 273196 25681 273212
rect 26681 273380 26778 273396
rect 26681 273212 26728 273380
rect 26762 273212 26778 273380
rect 26681 273196 26778 273212
rect 25584 273122 25681 273138
rect 25584 272954 25600 273122
rect 25634 272954 25681 273122
rect 25584 272938 25681 272954
rect 26681 273122 26778 273138
rect 26681 272954 26728 273122
rect 26762 272954 26778 273122
rect 26681 272938 26778 272954
rect 25584 272864 25681 272880
rect 25584 272696 25600 272864
rect 25634 272696 25681 272864
rect 25584 272680 25681 272696
rect 26681 272864 26778 272880
rect 26681 272696 26728 272864
rect 26762 272696 26778 272864
rect 26681 272680 26778 272696
rect 25584 272606 25681 272622
rect 25584 272438 25600 272606
rect 25634 272438 25681 272606
rect 25584 272422 25681 272438
rect 26681 272606 26778 272622
rect 26681 272438 26728 272606
rect 26762 272438 26778 272606
rect 26681 272422 26778 272438
rect 25584 272348 25681 272364
rect 25584 272180 25600 272348
rect 25634 272180 25681 272348
rect 25584 272164 25681 272180
rect 26681 272348 26778 272364
rect 26681 272180 26728 272348
rect 26762 272180 26778 272348
rect 26681 272164 26778 272180
rect 25584 272090 25681 272106
rect 25584 271922 25600 272090
rect 25634 271922 25681 272090
rect 25584 271906 25681 271922
rect 26681 272090 26778 272106
rect 26681 271922 26728 272090
rect 26762 271922 26778 272090
rect 26681 271906 26778 271922
rect 27202 272748 27290 272764
rect 27202 272680 27218 272748
rect 27252 272680 27290 272748
rect 27202 272664 27290 272680
rect 27790 272748 27878 272764
rect 27790 272680 27828 272748
rect 27862 272680 27878 272748
rect 27790 272664 27878 272680
rect 27202 272590 27290 272606
rect 27202 272522 27218 272590
rect 27252 272522 27290 272590
rect 27202 272506 27290 272522
rect 27790 272590 27878 272606
rect 27790 272522 27828 272590
rect 27862 272522 27878 272590
rect 27790 272506 27878 272522
rect 28202 273104 28290 273120
rect 28202 272936 28218 273104
rect 28252 272936 28290 273104
rect 28202 272920 28290 272936
rect 28540 273104 28628 273120
rect 28540 272936 28578 273104
rect 28612 272936 28628 273104
rect 28540 272920 28628 272936
rect 28202 272846 28290 272862
rect 28202 272678 28218 272846
rect 28252 272678 28290 272846
rect 28202 272662 28290 272678
rect 28540 272846 28628 272862
rect 28540 272678 28578 272846
rect 28612 272678 28628 272846
rect 28540 272662 28628 272678
rect 28202 272588 28290 272604
rect 28202 272420 28218 272588
rect 28252 272420 28290 272588
rect 28202 272404 28290 272420
rect 28540 272588 28628 272604
rect 28540 272420 28578 272588
rect 28612 272420 28628 272588
rect 28540 272404 28628 272420
rect 28202 272330 28290 272346
rect 28202 272162 28218 272330
rect 28252 272162 28290 272330
rect 28202 272146 28290 272162
rect 28540 272330 28628 272346
rect 28540 272162 28578 272330
rect 28612 272162 28628 272330
rect 28540 272146 28628 272162
rect 28952 273365 29040 273381
rect 28952 273197 28968 273365
rect 29002 273197 29040 273365
rect 28952 273181 29040 273197
rect 30040 273365 30128 273381
rect 30040 273197 30078 273365
rect 30112 273197 30128 273365
rect 30040 273181 30128 273197
rect 28952 273107 29040 273123
rect 28952 272939 28968 273107
rect 29002 272939 29040 273107
rect 28952 272923 29040 272939
rect 30040 273107 30128 273123
rect 30040 272939 30078 273107
rect 30112 272939 30128 273107
rect 30040 272923 30128 272939
rect 28952 272849 29040 272865
rect 28952 272681 28968 272849
rect 29002 272681 29040 272849
rect 28952 272665 29040 272681
rect 30040 272849 30128 272865
rect 30040 272681 30078 272849
rect 30112 272681 30128 272849
rect 30040 272665 30128 272681
rect 28952 272591 29040 272607
rect 28952 272423 28968 272591
rect 29002 272423 29040 272591
rect 28952 272407 29040 272423
rect 30040 272591 30128 272607
rect 30040 272423 30078 272591
rect 30112 272423 30128 272591
rect 30040 272407 30128 272423
rect 28952 272333 29040 272349
rect 28952 272165 28968 272333
rect 29002 272165 29040 272333
rect 28952 272149 29040 272165
rect 30040 272333 30128 272349
rect 30040 272165 30078 272333
rect 30112 272165 30128 272333
rect 30040 272149 30128 272165
rect 28952 272075 29040 272091
rect 28952 271907 28968 272075
rect 29002 271907 29040 272075
rect 28952 271891 29040 271907
rect 30040 272075 30128 272091
rect 30040 271907 30078 272075
rect 30112 271907 30128 272075
rect 30040 271891 30128 271907
rect 5902 252318 5968 252331
rect 5902 252315 5990 252318
rect 5902 252281 5918 252315
rect 5952 252281 5990 252315
rect 5902 252278 5990 252281
rect 15990 252278 16016 252318
rect 5902 252265 5968 252278
rect 16012 252220 16078 252233
rect 5964 252180 5990 252220
rect 15990 252217 16078 252220
rect 15990 252183 16028 252217
rect 16062 252183 16078 252217
rect 15990 252180 16078 252183
rect 5902 252122 5968 252135
rect 16012 252167 16078 252180
rect 5902 252119 5990 252122
rect 5902 252085 5918 252119
rect 5952 252085 5990 252119
rect 5902 252082 5990 252085
rect 15990 252082 16016 252122
rect 5902 252069 5968 252082
rect 16012 252024 16078 252037
rect 5964 251984 5990 252024
rect 15990 252021 16078 252024
rect 15990 251987 16028 252021
rect 16062 251987 16078 252021
rect 15990 251984 16078 251987
rect 5902 251926 5968 251939
rect 16012 251971 16078 251984
rect 5902 251923 5990 251926
rect 5902 251889 5918 251923
rect 5952 251889 5990 251923
rect 5902 251886 5990 251889
rect 15990 251886 16016 251926
rect 5902 251873 5968 251886
rect 16012 251828 16078 251841
rect 5964 251788 5990 251828
rect 15990 251825 16078 251828
rect 15990 251791 16028 251825
rect 16062 251791 16078 251825
rect 15990 251788 16078 251791
rect 5902 251730 5968 251743
rect 16012 251775 16078 251788
rect 5902 251727 5990 251730
rect 5902 251693 5918 251727
rect 5952 251693 5990 251727
rect 5902 251690 5990 251693
rect 15990 251690 16016 251730
rect 5902 251677 5968 251690
rect 16012 251632 16078 251645
rect 5964 251592 5990 251632
rect 15990 251629 16078 251632
rect 15990 251595 16028 251629
rect 16062 251595 16078 251629
rect 15990 251592 16078 251595
rect 5902 251534 5968 251547
rect 16012 251579 16078 251592
rect 5902 251531 5990 251534
rect 5902 251497 5918 251531
rect 5952 251497 5990 251531
rect 5902 251494 5990 251497
rect 15990 251494 16016 251534
rect 5902 251481 5968 251494
rect 16012 251436 16078 251449
rect 5964 251396 5990 251436
rect 15990 251433 16078 251436
rect 15990 251399 16028 251433
rect 16062 251399 16078 251433
rect 15990 251396 16078 251399
rect 16012 251383 16078 251396
rect 5902 241918 5968 241931
rect 5902 241915 5990 241918
rect 5902 241881 5918 241915
rect 5952 241881 5990 241915
rect 5902 241878 5990 241881
rect 15990 241878 16016 241918
rect 5902 241865 5968 241878
rect 16012 241820 16078 241833
rect 5964 241780 5990 241820
rect 15990 241817 16078 241820
rect 15990 241783 16028 241817
rect 16062 241783 16078 241817
rect 15990 241780 16078 241783
rect 5902 241722 5968 241735
rect 16012 241767 16078 241780
rect 5902 241719 5990 241722
rect 5902 241685 5918 241719
rect 5952 241685 5990 241719
rect 5902 241682 5990 241685
rect 15990 241682 16016 241722
rect 5902 241669 5968 241682
rect 16012 241624 16078 241637
rect 5964 241584 5990 241624
rect 15990 241621 16078 241624
rect 15990 241587 16028 241621
rect 16062 241587 16078 241621
rect 15990 241584 16078 241587
rect 5902 241526 5968 241539
rect 16012 241571 16078 241584
rect 5902 241523 5990 241526
rect 5902 241489 5918 241523
rect 5952 241489 5990 241523
rect 5902 241486 5990 241489
rect 15990 241486 16016 241526
rect 5902 241473 5968 241486
rect 16012 241428 16078 241441
rect 5964 241388 5990 241428
rect 15990 241425 16078 241428
rect 15990 241391 16028 241425
rect 16062 241391 16078 241425
rect 15990 241388 16078 241391
rect 5902 241330 5968 241343
rect 16012 241375 16078 241388
rect 5902 241327 5990 241330
rect 5902 241293 5918 241327
rect 5952 241293 5990 241327
rect 5902 241290 5990 241293
rect 15990 241290 16016 241330
rect 5902 241277 5968 241290
rect 16012 241232 16078 241245
rect 5964 241192 5990 241232
rect 15990 241229 16078 241232
rect 15990 241195 16028 241229
rect 16062 241195 16078 241229
rect 15990 241192 16078 241195
rect 5902 241134 5968 241147
rect 16012 241179 16078 241192
rect 5902 241131 5990 241134
rect 5902 241097 5918 241131
rect 5952 241097 5990 241131
rect 5902 241094 5990 241097
rect 15990 241094 16016 241134
rect 5902 241081 5968 241094
rect 16012 241036 16078 241049
rect 5964 240996 5990 241036
rect 15990 241033 16078 241036
rect 15990 240999 16028 241033
rect 16062 240999 16078 241033
rect 15990 240996 16078 240999
rect 16012 240983 16078 240996
<< polycont >>
rect 5918 304281 5952 304315
rect 16028 304183 16062 304217
rect 5918 304085 5952 304119
rect 16028 303987 16062 304021
rect 5918 303889 5952 303923
rect 16028 303791 16062 303825
rect 5918 303693 5952 303727
rect 16028 303595 16062 303629
rect 5918 303497 5952 303531
rect 16028 303399 16062 303433
rect 560097 305848 560131 305882
rect 560293 305848 560327 305882
rect 560489 305848 560523 305882
rect 560685 305848 560719 305882
rect 560881 305848 560915 305882
rect 559999 295738 560033 295772
rect 560195 295738 560229 295772
rect 560391 295738 560425 295772
rect 560587 295738 560621 295772
rect 560783 295738 560817 295772
rect 569297 305848 569331 305882
rect 569493 305848 569527 305882
rect 569689 305848 569723 305882
rect 569885 305848 569919 305882
rect 570081 305848 570115 305882
rect 569199 295738 569233 295772
rect 569395 295738 569429 295772
rect 569591 295738 569625 295772
rect 569787 295738 569821 295772
rect 569983 295738 570017 295772
rect 536287 294654 536321 294722
rect 537415 294654 537449 294722
rect 537523 294654 537557 294722
rect 538651 294654 538685 294722
rect 538759 294654 538793 294722
rect 539887 294654 539921 294722
rect 539995 294654 540029 294722
rect 541123 294654 541157 294722
rect 541231 294654 541265 294722
rect 542359 294654 542393 294722
rect 542467 294654 542501 294722
rect 543595 294654 543629 294722
rect 543703 294654 543737 294722
rect 544831 294654 544865 294722
rect 5918 293881 5952 293915
rect 16028 293783 16062 293817
rect 5918 293685 5952 293719
rect 16028 293587 16062 293621
rect 5918 293489 5952 293523
rect 16028 293391 16062 293425
rect 5918 293293 5952 293327
rect 16028 293195 16062 293229
rect 5918 293097 5952 293131
rect 16028 292999 16062 293033
rect 536287 294114 536321 294182
rect 537415 294114 537449 294182
rect 537523 294114 537557 294182
rect 538651 294114 538685 294182
rect 538759 294114 538793 294182
rect 539887 294114 539921 294182
rect 539995 294114 540029 294182
rect 541123 294114 541157 294182
rect 541231 294114 541265 294182
rect 542359 294114 542393 294182
rect 542467 294114 542501 294182
rect 543595 294114 543629 294182
rect 543703 294114 543737 294182
rect 544831 294114 544865 294182
rect 536287 293574 536321 293642
rect 537415 293574 537449 293642
rect 537523 293574 537557 293642
rect 538651 293574 538685 293642
rect 538759 293574 538793 293642
rect 539887 293574 539921 293642
rect 539995 293574 540029 293642
rect 541123 293574 541157 293642
rect 541231 293574 541265 293642
rect 542359 293574 542393 293642
rect 542467 293574 542501 293642
rect 543595 293574 543629 293642
rect 543703 293574 543737 293642
rect 544831 293574 544865 293642
rect 536287 293034 536321 293102
rect 537415 293034 537449 293102
rect 537523 293034 537557 293102
rect 538651 293034 538685 293102
rect 538759 293034 538793 293102
rect 539887 293034 539921 293102
rect 539995 293034 540029 293102
rect 541123 293034 541157 293102
rect 541231 293034 541265 293102
rect 542359 293034 542393 293102
rect 542467 293034 542501 293102
rect 543595 293034 543629 293102
rect 543703 293034 543737 293102
rect 544831 293034 544865 293102
rect 536287 292454 536321 292522
rect 537415 292454 537449 292522
rect 537523 292454 537557 292522
rect 538651 292454 538685 292522
rect 538759 292454 538793 292522
rect 539887 292454 539921 292522
rect 539995 292454 540029 292522
rect 541123 292454 541157 292522
rect 541231 292454 541265 292522
rect 542359 292454 542393 292522
rect 542467 292454 542501 292522
rect 543595 292454 543629 292522
rect 543703 292454 543737 292522
rect 544831 292454 544865 292522
rect 536287 291874 536321 291942
rect 537415 291874 537449 291942
rect 537523 291874 537557 291942
rect 538651 291874 538685 291942
rect 538759 291874 538793 291942
rect 539887 291874 539921 291942
rect 539995 291874 540029 291942
rect 541123 291874 541157 291942
rect 541231 291874 541265 291942
rect 542359 291874 542393 291942
rect 542467 291874 542501 291942
rect 543595 291874 543629 291942
rect 543703 291874 543737 291942
rect 544831 291874 544865 291942
rect 534447 291334 534481 291402
rect 535575 291334 535609 291402
rect 535683 291334 535717 291402
rect 536811 291334 536845 291402
rect 536919 291334 536953 291402
rect 538047 291334 538081 291402
rect 538155 291334 538189 291402
rect 539283 291334 539317 291402
rect 539391 291334 539425 291402
rect 540519 291334 540553 291402
rect 540627 291334 540661 291402
rect 541755 291334 541789 291402
rect 541863 291334 541897 291402
rect 542991 291334 543025 291402
rect 543099 291334 543133 291402
rect 544227 291334 544261 291402
rect 544335 291334 544369 291402
rect 545463 291334 545497 291402
rect 545571 291334 545605 291402
rect 546699 291334 546733 291402
rect 534447 290794 534481 290862
rect 535575 290794 535609 290862
rect 535683 290794 535717 290862
rect 536811 290794 536845 290862
rect 536919 290794 536953 290862
rect 538047 290794 538081 290862
rect 538155 290794 538189 290862
rect 539283 290794 539317 290862
rect 539391 290794 539425 290862
rect 540519 290794 540553 290862
rect 540627 290794 540661 290862
rect 541755 290794 541789 290862
rect 541863 290794 541897 290862
rect 542991 290794 543025 290862
rect 543099 290794 543133 290862
rect 544227 290794 544261 290862
rect 544335 290794 544369 290862
rect 545463 290794 545497 290862
rect 545571 290794 545605 290862
rect 546699 290794 546733 290862
rect 534447 290254 534481 290322
rect 535575 290254 535609 290322
rect 535683 290254 535717 290322
rect 536811 290254 536845 290322
rect 536919 290254 536953 290322
rect 538047 290254 538081 290322
rect 538155 290254 538189 290322
rect 539283 290254 539317 290322
rect 539391 290254 539425 290322
rect 540519 290254 540553 290322
rect 540627 290254 540661 290322
rect 541755 290254 541789 290322
rect 541863 290254 541897 290322
rect 542991 290254 543025 290322
rect 543099 290254 543133 290322
rect 544227 290254 544261 290322
rect 544335 290254 544369 290322
rect 545463 290254 545497 290322
rect 545571 290254 545605 290322
rect 546699 290254 546733 290322
rect 534447 289714 534481 289782
rect 535575 289714 535609 289782
rect 535683 289714 535717 289782
rect 536811 289714 536845 289782
rect 536919 289714 536953 289782
rect 538047 289714 538081 289782
rect 538155 289714 538189 289782
rect 539283 289714 539317 289782
rect 539391 289714 539425 289782
rect 540519 289714 540553 289782
rect 540627 289714 540661 289782
rect 541755 289714 541789 289782
rect 541863 289714 541897 289782
rect 542991 289714 543025 289782
rect 543099 289714 543133 289782
rect 544227 289714 544261 289782
rect 544335 289714 544369 289782
rect 545463 289714 545497 289782
rect 545571 289714 545605 289782
rect 546699 289714 546733 289782
rect 536387 288934 536421 289002
rect 537497 288934 537531 289002
rect 537605 288934 537639 289002
rect 538715 288934 538749 289002
rect 538823 288934 538857 289002
rect 539933 288934 539967 289002
rect 540041 288934 540075 289002
rect 541151 288934 541185 289002
rect 541259 288934 541293 289002
rect 542369 288934 542403 289002
rect 542477 288934 542511 289002
rect 543587 288934 543621 289002
rect 543695 288934 543729 289002
rect 544805 288934 544839 289002
rect 536387 288434 536421 288502
rect 537497 288434 537531 288502
rect 537605 288434 537639 288502
rect 538715 288434 538749 288502
rect 538823 288434 538857 288502
rect 539933 288434 539967 288502
rect 540041 288434 540075 288502
rect 541151 288434 541185 288502
rect 541259 288434 541293 288502
rect 542369 288434 542403 288502
rect 542477 288434 542511 288502
rect 543587 288434 543621 288502
rect 543695 288434 543729 288502
rect 544805 288434 544839 288502
rect 536947 287834 536981 288002
rect 538057 287834 538091 288002
rect 538165 287834 538199 288002
rect 539275 287834 539309 288002
rect 539383 287834 539417 288002
rect 540493 287834 540527 288002
rect 540601 287834 540635 288002
rect 541711 287834 541745 288002
rect 541819 287834 541853 288002
rect 542929 287834 542963 288002
rect 543037 287834 543071 288002
rect 544147 287834 544181 288002
rect 568218 288661 568252 288695
rect 578328 288563 578362 288597
rect 568218 288465 568252 288499
rect 578328 288367 578362 288401
rect 568218 288269 568252 288303
rect 578328 288171 578362 288205
rect 568218 288073 568252 288107
rect 578328 287975 578362 288009
rect 568218 287877 568252 287911
rect 578328 287779 578362 287813
rect 536947 287214 536981 287382
rect 538057 287214 538091 287382
rect 538165 287214 538199 287382
rect 539275 287214 539309 287382
rect 539383 287214 539417 287382
rect 540493 287214 540527 287382
rect 540601 287214 540635 287382
rect 541711 287214 541745 287382
rect 541819 287214 541853 287382
rect 542929 287214 542963 287382
rect 543037 287214 543071 287382
rect 544147 287214 544181 287382
rect 536387 286614 536421 286782
rect 537497 286614 537531 286782
rect 537605 286614 537639 286782
rect 538715 286614 538749 286782
rect 538823 286614 538857 286782
rect 539933 286614 539967 286782
rect 540041 286614 540075 286782
rect 541151 286614 541185 286782
rect 541259 286614 541293 286782
rect 542369 286614 542403 286782
rect 542477 286614 542511 286782
rect 543587 286614 543621 286782
rect 543695 286614 543729 286782
rect 544805 286614 544839 286782
rect 536387 286014 536421 286182
rect 537497 286014 537531 286182
rect 537605 286014 537639 286182
rect 538715 286014 538749 286182
rect 538823 286014 538857 286182
rect 539933 286014 539967 286182
rect 540041 286014 540075 286182
rect 541151 286014 541185 286182
rect 541259 286014 541293 286182
rect 542369 286014 542403 286182
rect 542477 286014 542511 286182
rect 543587 286014 543621 286182
rect 543695 286014 543729 286182
rect 544805 286014 544839 286182
rect 536932 285040 536966 285208
rect 538060 285040 538094 285208
rect 538168 285040 538202 285208
rect 539296 285040 539330 285208
rect 539404 285040 539438 285208
rect 540532 285040 540566 285208
rect 540640 285040 540674 285208
rect 541768 285040 541802 285208
rect 541876 285040 541910 285208
rect 543004 285040 543038 285208
rect 543112 285040 543146 285208
rect 544240 285040 544274 285208
rect 536932 284450 536966 284618
rect 538060 284450 538094 284618
rect 538168 284450 538202 284618
rect 539296 284450 539330 284618
rect 539404 284450 539438 284618
rect 540532 284450 540566 284618
rect 540640 284450 540674 284618
rect 541768 284450 541802 284618
rect 541876 284450 541910 284618
rect 543004 284450 543038 284618
rect 543112 284450 543146 284618
rect 544240 284450 544274 284618
rect 539702 283660 539736 283828
rect 540062 283660 540096 283828
rect 540170 283660 540204 283828
rect 540530 283660 540564 283828
rect 540638 283660 540672 283828
rect 540998 283660 541032 283828
rect 541106 283660 541140 283828
rect 541466 283660 541500 283828
rect 539922 283135 539956 283203
rect 540532 283135 540566 283203
rect 540640 283135 540674 283203
rect 541250 283135 541284 283203
rect 536987 282510 537021 282678
rect 538097 282510 538131 282678
rect 538205 282510 538239 282678
rect 539315 282510 539349 282678
rect 539423 282510 539457 282678
rect 540533 282510 540567 282678
rect 540641 282510 540675 282678
rect 541751 282510 541785 282678
rect 541859 282510 541893 282678
rect 542969 282510 543003 282678
rect 543077 282510 543111 282678
rect 544187 282510 544221 282678
rect 568238 281181 568272 281215
rect 578348 281083 578382 281117
rect 568238 280985 568272 281019
rect 578348 280887 578382 280921
rect 568238 280789 568272 280823
rect 578348 280691 578382 280725
rect 568238 280593 568272 280627
rect 578348 280495 578382 280529
rect 568238 280397 568272 280431
rect 578348 280299 578382 280333
rect 12720 275704 12754 275772
rect 13848 275704 13882 275772
rect 12720 275546 12754 275614
rect 13848 275546 13882 275614
rect 12720 275388 12754 275456
rect 13848 275388 13882 275456
rect 12720 275230 12754 275298
rect 13848 275230 13882 275298
rect 12720 275072 12754 275140
rect 13848 275072 13882 275140
rect 12720 274914 12754 274982
rect 13848 274914 13882 274982
rect 12720 274756 12754 274824
rect 13848 274756 13882 274824
rect 12720 274598 12754 274666
rect 13848 274598 13882 274666
rect 12720 274440 12754 274508
rect 13848 274440 13882 274508
rect 12720 274282 12754 274350
rect 13848 274282 13882 274350
rect 12720 274124 12754 274192
rect 13848 274124 13882 274192
rect 12720 273966 12754 274034
rect 13848 273966 13882 274034
rect 12720 273808 12754 273876
rect 13848 273808 13882 273876
rect 12720 273650 12754 273718
rect 13848 273650 13882 273718
rect 12720 273492 12754 273560
rect 13848 273492 13882 273560
rect 12720 273334 12754 273402
rect 13848 273334 13882 273402
rect 12720 273176 12754 273244
rect 13848 273176 13882 273244
rect 12720 273018 12754 273086
rect 13848 273018 13882 273086
rect 12720 272860 12754 272928
rect 13848 272860 13882 272928
rect 12720 272702 12754 272770
rect 13848 272702 13882 272770
rect 12720 272544 12754 272612
rect 13848 272544 13882 272612
rect 12720 272386 12754 272454
rect 13848 272386 13882 272454
rect 12720 272228 12754 272296
rect 13848 272228 13882 272296
rect 12720 272070 12754 272138
rect 13848 272070 13882 272138
rect 12720 271912 12754 271980
rect 13848 271912 13882 271980
rect 12720 271754 12754 271822
rect 13848 271754 13882 271822
rect 12720 271596 12754 271664
rect 13848 271596 13882 271664
rect 12720 271438 12754 271506
rect 13848 271438 13882 271506
rect 12720 271280 12754 271348
rect 13848 271280 13882 271348
rect 12720 271122 12754 271190
rect 13848 271122 13882 271190
rect 12720 270964 12754 271032
rect 13848 270964 13882 271032
rect 12720 270806 12754 270874
rect 13848 270806 13882 270874
rect 12720 270648 12754 270716
rect 13848 270648 13882 270716
rect 12720 270490 12754 270558
rect 13848 270490 13882 270558
rect 12720 270332 12754 270400
rect 13848 270332 13882 270400
rect 12720 270174 12754 270242
rect 13848 270174 13882 270242
rect 12720 270016 12754 270084
rect 13848 270016 13882 270084
rect 12720 269858 12754 269926
rect 13848 269858 13882 269926
rect 12720 269700 12754 269768
rect 13848 269700 13882 269768
rect 12720 269542 12754 269610
rect 13848 269542 13882 269610
rect 14390 274202 14424 274270
rect 15518 274202 15552 274270
rect 14390 274044 14424 274112
rect 15518 274044 15552 274112
rect 14390 273886 14424 273954
rect 15518 273886 15552 273954
rect 14390 273728 14424 273796
rect 15518 273728 15552 273796
rect 14390 273570 14424 273638
rect 15518 273570 15552 273638
rect 14390 273412 14424 273480
rect 15518 273412 15552 273480
rect 14390 273254 14424 273322
rect 15518 273254 15552 273322
rect 14390 273096 14424 273164
rect 15518 273096 15552 273164
rect 14390 272938 14424 273006
rect 15518 272938 15552 273006
rect 14390 272780 14424 272848
rect 15518 272780 15552 272848
rect 14390 272622 14424 272690
rect 15518 272622 15552 272690
rect 14390 272464 14424 272532
rect 15518 272464 15552 272532
rect 14390 272306 14424 272374
rect 15518 272306 15552 272374
rect 14390 272148 14424 272216
rect 15518 272148 15552 272216
rect 14390 271990 14424 272058
rect 15518 271990 15552 272058
rect 14390 271832 14424 271900
rect 15518 271832 15552 271900
rect 14390 271674 14424 271742
rect 15518 271674 15552 271742
rect 14390 271516 14424 271584
rect 15518 271516 15552 271584
rect 14390 271358 14424 271426
rect 15518 271358 15552 271426
rect 14390 271200 14424 271268
rect 15518 271200 15552 271268
rect 14390 271042 14424 271110
rect 15518 271042 15552 271110
rect 15930 274202 15964 274270
rect 17058 274202 17092 274270
rect 15930 274044 15964 274112
rect 17058 274044 17092 274112
rect 15930 273886 15964 273954
rect 17058 273886 17092 273954
rect 15930 273728 15964 273796
rect 17058 273728 17092 273796
rect 15930 273570 15964 273638
rect 17058 273570 17092 273638
rect 15930 273412 15964 273480
rect 17058 273412 17092 273480
rect 15930 273254 15964 273322
rect 17058 273254 17092 273322
rect 15930 273096 15964 273164
rect 17058 273096 17092 273164
rect 15930 272938 15964 273006
rect 17058 272938 17092 273006
rect 15930 272780 15964 272848
rect 17058 272780 17092 272848
rect 15930 272622 15964 272690
rect 17058 272622 17092 272690
rect 15930 272464 15964 272532
rect 17058 272464 17092 272532
rect 15930 272306 15964 272374
rect 17058 272306 17092 272374
rect 15930 272148 15964 272216
rect 17058 272148 17092 272216
rect 15930 271990 15964 272058
rect 17058 271990 17092 272058
rect 15930 271832 15964 271900
rect 17058 271832 17092 271900
rect 15930 271674 15964 271742
rect 17058 271674 17092 271742
rect 15930 271516 15964 271584
rect 17058 271516 17092 271584
rect 15930 271358 15964 271426
rect 17058 271358 17092 271426
rect 15930 271200 15964 271268
rect 17058 271200 17092 271268
rect 15930 271042 15964 271110
rect 17058 271042 17092 271110
rect 17507 273091 17541 273159
rect 18617 273091 18651 273159
rect 17507 272933 17541 273001
rect 18617 272933 18651 273001
rect 17507 272775 17541 272843
rect 18617 272775 18651 272843
rect 17507 272617 17541 272685
rect 18617 272617 18651 272685
rect 17507 272459 17541 272527
rect 18617 272459 18651 272527
rect 17507 272301 17541 272369
rect 18617 272301 18651 272369
rect 17507 272143 17541 272211
rect 18617 272143 18651 272211
rect 19027 273091 19061 273159
rect 20137 273091 20171 273159
rect 19027 272933 19061 273001
rect 20137 272933 20171 273001
rect 19027 272775 19061 272843
rect 20137 272775 20171 272843
rect 19027 272617 19061 272685
rect 20137 272617 20171 272685
rect 19027 272459 19061 272527
rect 20137 272459 20171 272527
rect 19027 272301 19061 272369
rect 20137 272301 20171 272369
rect 19027 272143 19061 272211
rect 20137 272143 20171 272211
rect 20548 273990 20582 274158
rect 21658 273990 21692 274158
rect 20548 273732 20582 273900
rect 21658 273732 21692 273900
rect 20548 273474 20582 273642
rect 21658 273474 21692 273642
rect 20548 273216 20582 273384
rect 21658 273216 21692 273384
rect 20548 272958 20582 273126
rect 21658 272958 21692 273126
rect 20548 272700 20582 272868
rect 21658 272700 21692 272868
rect 20548 272442 20582 272610
rect 21658 272442 21692 272610
rect 20548 272184 20582 272352
rect 21658 272184 21692 272352
rect 20548 271926 20582 272094
rect 21658 271926 21692 272094
rect 20548 271668 20582 271836
rect 21658 271668 21692 271836
rect 20548 271410 20582 271578
rect 21658 271410 21692 271578
rect 20548 271152 20582 271320
rect 21658 271152 21692 271320
rect 22068 274246 22102 274414
rect 23178 274246 23212 274414
rect 22068 273988 22102 274156
rect 23178 273988 23212 274156
rect 22068 273730 22102 273898
rect 23178 273730 23212 273898
rect 22068 273472 22102 273640
rect 23178 273472 23212 273640
rect 22068 273214 22102 273382
rect 23178 273214 23212 273382
rect 22068 272956 22102 273124
rect 23178 272956 23212 273124
rect 22068 272698 22102 272866
rect 23178 272698 23212 272866
rect 22068 272440 22102 272608
rect 23178 272440 23212 272608
rect 22068 272182 22102 272350
rect 23178 272182 23212 272350
rect 22068 271924 22102 272092
rect 23178 271924 23212 272092
rect 22068 271666 22102 271834
rect 23178 271666 23212 271834
rect 22068 271408 22102 271576
rect 23178 271408 23212 271576
rect 22068 271150 22102 271318
rect 23178 271150 23212 271318
rect 22068 270892 22102 271060
rect 23178 270892 23212 271060
rect 24100 273212 24134 273380
rect 25228 273212 25262 273380
rect 24100 272954 24134 273122
rect 25228 272954 25262 273122
rect 24100 272696 24134 272864
rect 25228 272696 25262 272864
rect 24100 272438 24134 272606
rect 25228 272438 25262 272606
rect 24100 272180 24134 272348
rect 25228 272180 25262 272348
rect 24100 271922 24134 272090
rect 25228 271922 25262 272090
rect 25600 273212 25634 273380
rect 26728 273212 26762 273380
rect 25600 272954 25634 273122
rect 26728 272954 26762 273122
rect 25600 272696 25634 272864
rect 26728 272696 26762 272864
rect 25600 272438 25634 272606
rect 26728 272438 26762 272606
rect 25600 272180 25634 272348
rect 26728 272180 26762 272348
rect 25600 271922 25634 272090
rect 26728 271922 26762 272090
rect 27218 272680 27252 272748
rect 27828 272680 27862 272748
rect 27218 272522 27252 272590
rect 27828 272522 27862 272590
rect 28218 272936 28252 273104
rect 28578 272936 28612 273104
rect 28218 272678 28252 272846
rect 28578 272678 28612 272846
rect 28218 272420 28252 272588
rect 28578 272420 28612 272588
rect 28218 272162 28252 272330
rect 28578 272162 28612 272330
rect 28968 273197 29002 273365
rect 30078 273197 30112 273365
rect 28968 272939 29002 273107
rect 30078 272939 30112 273107
rect 28968 272681 29002 272849
rect 30078 272681 30112 272849
rect 28968 272423 29002 272591
rect 30078 272423 30112 272591
rect 28968 272165 29002 272333
rect 30078 272165 30112 272333
rect 28968 271907 29002 272075
rect 30078 271907 30112 272075
rect 5918 252281 5952 252315
rect 16028 252183 16062 252217
rect 5918 252085 5952 252119
rect 16028 251987 16062 252021
rect 5918 251889 5952 251923
rect 16028 251791 16062 251825
rect 5918 251693 5952 251727
rect 16028 251595 16062 251629
rect 5918 251497 5952 251531
rect 16028 251399 16062 251433
rect 5918 241881 5952 241915
rect 16028 241783 16062 241817
rect 5918 241685 5952 241719
rect 16028 241587 16062 241621
rect 5918 241489 5952 241523
rect 16028 241391 16062 241425
rect 5918 241293 5952 241327
rect 16028 241195 16062 241229
rect 5918 241097 5952 241131
rect 16028 240999 16062 241033
<< xpolycontact >>
rect 530722 290825 531154 291971
rect 533154 290825 533586 291971
rect 547782 290825 548214 291971
rect 550214 290825 550646 291971
rect 530722 289355 531154 290501
rect 533154 289355 533586 290501
rect 547782 289355 548214 290501
rect 550214 289355 550646 290501
rect 537761 281570 538907 282002
rect 539281 281570 540427 282002
rect 540791 281576 541937 282008
rect 542301 281576 543447 282008
rect 11871 279195 13017 279627
rect 11871 276763 13017 277195
rect 13331 279195 14477 279627
rect 13331 276763 14477 277195
rect 11871 268125 13017 268557
rect 11871 265693 13017 266125
rect 13331 268125 14477 268557
rect 13331 265693 14477 266125
rect 537761 267338 538907 267770
rect 539281 267338 540427 267770
rect 540791 267344 541937 267776
rect 542301 267344 543447 267776
<< locali >>
rect 559836 305950 561078 305984
rect 559836 305888 559870 305950
rect 5816 304444 5912 304478
rect 16068 304444 16164 304478
rect 5816 303270 5850 304444
rect 16130 304382 16164 304444
rect 5918 304315 5952 304331
rect 5986 304330 6002 304364
rect 15978 304330 15994 304364
rect 5918 304265 5952 304281
rect 5986 304232 6002 304266
rect 15978 304232 15994 304266
rect 16028 304217 16062 304233
rect 5918 304119 5952 304135
rect 5986 304134 6002 304168
rect 15978 304134 15994 304168
rect 16028 304167 16062 304183
rect 5918 304069 5952 304085
rect 5986 304036 6002 304070
rect 15978 304036 15994 304070
rect 16028 304021 16062 304037
rect 5918 303923 5952 303939
rect 5986 303938 6002 303972
rect 15978 303938 15994 303972
rect 16028 303971 16062 303987
rect 5918 303873 5952 303889
rect 5986 303840 6002 303874
rect 15978 303840 15994 303874
rect 16028 303825 16062 303841
rect 5918 303727 5952 303743
rect 5986 303742 6002 303776
rect 15978 303742 15994 303776
rect 16028 303775 16062 303791
rect 5918 303677 5952 303693
rect 5986 303644 6002 303678
rect 15978 303644 15994 303678
rect 16028 303629 16062 303645
rect 5918 303531 5952 303547
rect 5986 303546 6002 303580
rect 15978 303546 15994 303580
rect 16028 303579 16062 303595
rect 5918 303481 5952 303497
rect 5986 303448 6002 303482
rect 15978 303448 15994 303482
rect 16028 303433 16062 303449
rect 5986 303350 6002 303384
rect 15978 303350 15994 303384
rect 16028 303383 16062 303399
rect 16130 303270 16164 303332
rect 5816 303236 5912 303270
rect 16068 303236 16164 303270
rect 561044 305888 561078 305950
rect 560081 305848 560097 305882
rect 560131 305848 560147 305882
rect 560277 305848 560293 305882
rect 560327 305848 560343 305882
rect 560473 305848 560489 305882
rect 560523 305848 560539 305882
rect 560669 305848 560685 305882
rect 560719 305848 560735 305882
rect 560865 305848 560881 305882
rect 560915 305848 560931 305882
rect 559950 305798 559984 305814
rect 559950 295806 559984 295822
rect 560048 305798 560082 305814
rect 560048 295806 560082 295822
rect 560146 305798 560180 305814
rect 560146 295806 560180 295822
rect 560244 305798 560278 305814
rect 560244 295806 560278 295822
rect 560342 305798 560376 305814
rect 560342 295806 560376 295822
rect 560440 305798 560474 305814
rect 560440 295806 560474 295822
rect 560538 305798 560572 305814
rect 560538 295806 560572 295822
rect 560636 305798 560670 305814
rect 560636 295806 560670 295822
rect 560734 305798 560768 305814
rect 560734 295806 560768 295822
rect 560832 305798 560866 305814
rect 560832 295806 560866 295822
rect 560930 305798 560964 305814
rect 560930 295806 560964 295822
rect 559983 295738 559999 295772
rect 560033 295738 560049 295772
rect 560179 295738 560195 295772
rect 560229 295738 560245 295772
rect 560375 295738 560391 295772
rect 560425 295738 560441 295772
rect 560571 295738 560587 295772
rect 560621 295738 560637 295772
rect 560767 295738 560783 295772
rect 560817 295738 560833 295772
rect 559836 295670 559870 295732
rect 561044 295670 561078 295732
rect 559836 295636 559932 295670
rect 560982 295636 561078 295670
rect 569036 305950 570278 305984
rect 569036 305888 569070 305950
rect 570244 305888 570278 305950
rect 569281 305848 569297 305882
rect 569331 305848 569347 305882
rect 569477 305848 569493 305882
rect 569527 305848 569543 305882
rect 569673 305848 569689 305882
rect 569723 305848 569739 305882
rect 569869 305848 569885 305882
rect 569919 305848 569935 305882
rect 570065 305848 570081 305882
rect 570115 305848 570131 305882
rect 569150 305798 569184 305814
rect 569150 295806 569184 295822
rect 569248 305798 569282 305814
rect 569248 295806 569282 295822
rect 569346 305798 569380 305814
rect 569346 295806 569380 295822
rect 569444 305798 569478 305814
rect 569444 295806 569478 295822
rect 569542 305798 569576 305814
rect 569542 295806 569576 295822
rect 569640 305798 569674 305814
rect 569640 295806 569674 295822
rect 569738 305798 569772 305814
rect 569738 295806 569772 295822
rect 569836 305798 569870 305814
rect 569836 295806 569870 295822
rect 569934 305798 569968 305814
rect 569934 295806 569968 295822
rect 570032 305798 570066 305814
rect 570032 295806 570066 295822
rect 570130 305798 570164 305814
rect 570130 295806 570164 295822
rect 569183 295738 569199 295772
rect 569233 295738 569249 295772
rect 569379 295738 569395 295772
rect 569429 295738 569445 295772
rect 569575 295738 569591 295772
rect 569625 295738 569641 295772
rect 569771 295738 569787 295772
rect 569821 295738 569837 295772
rect 569967 295738 569983 295772
rect 570017 295738 570033 295772
rect 569036 295670 569070 295732
rect 570244 295670 570278 295732
rect 569036 295636 569132 295670
rect 570182 295636 570278 295670
rect 536185 294864 536281 294898
rect 544871 294864 544967 294898
rect 536185 294802 536219 294864
rect 544933 294802 544967 294864
rect 536364 294750 536380 294784
rect 537356 294750 537372 294784
rect 537600 294750 537616 294784
rect 538592 294750 538608 294784
rect 538836 294750 538852 294784
rect 539828 294750 539844 294784
rect 540072 294750 540088 294784
rect 541064 294750 541080 294784
rect 541308 294750 541324 294784
rect 542300 294750 542316 294784
rect 542544 294750 542560 294784
rect 543536 294750 543552 294784
rect 543780 294750 543796 294784
rect 544772 294750 544788 294784
rect 536287 294722 536321 294738
rect 536287 294638 536321 294654
rect 537415 294722 537449 294738
rect 537415 294638 537449 294654
rect 537523 294722 537557 294738
rect 537523 294638 537557 294654
rect 538651 294722 538685 294738
rect 538651 294638 538685 294654
rect 538759 294722 538793 294738
rect 538759 294638 538793 294654
rect 539887 294722 539921 294738
rect 539887 294638 539921 294654
rect 539995 294722 540029 294738
rect 539995 294638 540029 294654
rect 541123 294722 541157 294738
rect 541123 294638 541157 294654
rect 541231 294722 541265 294738
rect 541231 294638 541265 294654
rect 542359 294722 542393 294738
rect 542359 294638 542393 294654
rect 542467 294722 542501 294738
rect 542467 294638 542501 294654
rect 543595 294722 543629 294738
rect 543595 294638 543629 294654
rect 543703 294722 543737 294738
rect 543703 294638 543737 294654
rect 544831 294722 544865 294738
rect 544831 294638 544865 294654
rect 536364 294592 536380 294626
rect 537356 294592 537372 294626
rect 537600 294592 537616 294626
rect 538592 294592 538608 294626
rect 538836 294592 538852 294626
rect 539828 294592 539844 294626
rect 540072 294592 540088 294626
rect 541064 294592 541080 294626
rect 541308 294592 541324 294626
rect 542300 294592 542316 294626
rect 542544 294592 542560 294626
rect 543536 294592 543552 294626
rect 543780 294592 543796 294626
rect 544772 294592 544788 294626
rect 536185 294512 536219 294574
rect 544933 294512 544967 294574
rect 536185 294478 536281 294512
rect 544871 294478 544967 294512
rect 536185 294324 536281 294358
rect 544871 294324 544967 294358
rect 536185 294262 536219 294324
rect 5816 294044 5912 294078
rect 16068 294044 16164 294078
rect 5816 292870 5850 294044
rect 16130 293982 16164 294044
rect 5918 293915 5952 293931
rect 5986 293930 6002 293964
rect 15978 293930 15994 293964
rect 5918 293865 5952 293881
rect 5986 293832 6002 293866
rect 15978 293832 15994 293866
rect 16028 293817 16062 293833
rect 5918 293719 5952 293735
rect 5986 293734 6002 293768
rect 15978 293734 15994 293768
rect 16028 293767 16062 293783
rect 544933 294262 544967 294324
rect 536364 294210 536380 294244
rect 537356 294210 537372 294244
rect 537600 294210 537616 294244
rect 538592 294210 538608 294244
rect 538836 294210 538852 294244
rect 539828 294210 539844 294244
rect 540072 294210 540088 294244
rect 541064 294210 541080 294244
rect 541308 294210 541324 294244
rect 542300 294210 542316 294244
rect 542544 294210 542560 294244
rect 543536 294210 543552 294244
rect 543780 294210 543796 294244
rect 544772 294210 544788 294244
rect 536287 294182 536321 294198
rect 536287 294098 536321 294114
rect 537415 294182 537449 294198
rect 537415 294098 537449 294114
rect 537523 294182 537557 294198
rect 537523 294098 537557 294114
rect 538651 294182 538685 294198
rect 538651 294098 538685 294114
rect 538759 294182 538793 294198
rect 538759 294098 538793 294114
rect 539887 294182 539921 294198
rect 539887 294098 539921 294114
rect 539995 294182 540029 294198
rect 539995 294098 540029 294114
rect 541123 294182 541157 294198
rect 541123 294098 541157 294114
rect 541231 294182 541265 294198
rect 541231 294098 541265 294114
rect 542359 294182 542393 294198
rect 542359 294098 542393 294114
rect 542467 294182 542501 294198
rect 542467 294098 542501 294114
rect 543595 294182 543629 294198
rect 543595 294098 543629 294114
rect 543703 294182 543737 294198
rect 543703 294098 543737 294114
rect 544831 294182 544865 294198
rect 544831 294098 544865 294114
rect 536364 294052 536380 294086
rect 537356 294052 537372 294086
rect 537600 294052 537616 294086
rect 538592 294052 538608 294086
rect 538836 294052 538852 294086
rect 539828 294052 539844 294086
rect 540072 294052 540088 294086
rect 541064 294052 541080 294086
rect 541308 294052 541324 294086
rect 542300 294052 542316 294086
rect 542544 294052 542560 294086
rect 543536 294052 543552 294086
rect 543780 294052 543796 294086
rect 544772 294052 544788 294086
rect 536185 293972 536219 294034
rect 544933 293972 544967 294034
rect 536185 293938 536281 293972
rect 544871 293938 544967 293972
rect 537969 293912 538229 293938
rect 537969 293842 537979 293912
rect 538069 293842 538119 293912
rect 538209 293842 538229 293912
rect 537969 293818 538229 293842
rect 540439 293922 540729 293938
rect 540439 293912 540619 293922
rect 540439 293842 540459 293912
rect 540549 293852 540619 293912
rect 540709 293852 540729 293922
rect 540549 293842 540729 293852
rect 540439 293818 540729 293842
rect 542899 293922 543189 293938
rect 542899 293852 542919 293922
rect 542999 293852 543089 293922
rect 543169 293852 543189 293922
rect 542899 293818 543189 293852
rect 5918 293669 5952 293685
rect 5986 293636 6002 293670
rect 15978 293636 15994 293670
rect 16028 293621 16062 293637
rect 5918 293523 5952 293539
rect 5986 293538 6002 293572
rect 15978 293538 15994 293572
rect 16028 293571 16062 293587
rect 5918 293473 5952 293489
rect 5986 293440 6002 293474
rect 15978 293440 15994 293474
rect 16028 293425 16062 293441
rect 5918 293327 5952 293343
rect 5986 293342 6002 293376
rect 15978 293342 15994 293376
rect 16028 293375 16062 293391
rect 5918 293277 5952 293293
rect 5986 293244 6002 293278
rect 15978 293244 15994 293278
rect 16028 293229 16062 293245
rect 5918 293131 5952 293147
rect 5986 293146 6002 293180
rect 15978 293146 15994 293180
rect 16028 293179 16062 293195
rect 536185 293784 536281 293818
rect 544871 293784 544967 293818
rect 536185 293722 536219 293784
rect 544933 293722 544967 293784
rect 536364 293670 536380 293704
rect 537356 293670 537372 293704
rect 537600 293670 537616 293704
rect 538592 293670 538608 293704
rect 538836 293670 538852 293704
rect 539828 293670 539844 293704
rect 540072 293670 540088 293704
rect 541064 293670 541080 293704
rect 541308 293670 541324 293704
rect 542300 293670 542316 293704
rect 542544 293670 542560 293704
rect 543536 293670 543552 293704
rect 543780 293670 543796 293704
rect 544772 293670 544788 293704
rect 536287 293642 536321 293658
rect 536287 293558 536321 293574
rect 537415 293642 537449 293658
rect 537415 293558 537449 293574
rect 537523 293642 537557 293658
rect 537523 293558 537557 293574
rect 538651 293642 538685 293658
rect 538651 293558 538685 293574
rect 538759 293642 538793 293658
rect 538759 293558 538793 293574
rect 539887 293642 539921 293658
rect 539887 293558 539921 293574
rect 539995 293642 540029 293658
rect 539995 293558 540029 293574
rect 541123 293642 541157 293658
rect 541123 293558 541157 293574
rect 541231 293642 541265 293658
rect 541231 293558 541265 293574
rect 542359 293642 542393 293658
rect 542359 293558 542393 293574
rect 542467 293642 542501 293658
rect 542467 293558 542501 293574
rect 543595 293642 543629 293658
rect 543595 293558 543629 293574
rect 543703 293642 543737 293658
rect 543703 293558 543737 293574
rect 544831 293642 544865 293658
rect 544831 293558 544865 293574
rect 536364 293512 536380 293546
rect 537356 293512 537372 293546
rect 537600 293512 537616 293546
rect 538592 293512 538608 293546
rect 538836 293512 538852 293546
rect 539828 293512 539844 293546
rect 540072 293512 540088 293546
rect 541064 293512 541080 293546
rect 541308 293512 541324 293546
rect 542300 293512 542316 293546
rect 542544 293512 542560 293546
rect 543536 293512 543552 293546
rect 543780 293512 543796 293546
rect 544772 293512 544788 293546
rect 536185 293432 536219 293494
rect 544933 293432 544967 293494
rect 536185 293398 536281 293432
rect 544871 293398 544967 293432
rect 537959 293382 538249 293398
rect 537959 293302 537979 293382
rect 538059 293302 538149 293382
rect 538229 293302 538249 293382
rect 537959 293278 538249 293302
rect 540439 293382 540729 293398
rect 540439 293302 540459 293382
rect 540539 293302 540629 293382
rect 540709 293302 540729 293382
rect 540439 293278 540729 293302
rect 542899 293382 543189 293398
rect 542899 293302 542919 293382
rect 542999 293302 543089 293382
rect 543169 293302 543189 293382
rect 542899 293278 543189 293302
rect 5918 293081 5952 293097
rect 5986 293048 6002 293082
rect 15978 293048 15994 293082
rect 16028 293033 16062 293049
rect 5986 292950 6002 292984
rect 15978 292950 15994 292984
rect 16028 292983 16062 292999
rect 16130 292870 16164 292932
rect 5816 292836 5912 292870
rect 16068 292836 16164 292870
rect 536185 293244 536281 293278
rect 544871 293244 544967 293278
rect 536185 293182 536219 293244
rect 544933 293182 544967 293244
rect 536364 293130 536380 293164
rect 537356 293130 537372 293164
rect 537600 293130 537616 293164
rect 538592 293130 538608 293164
rect 538836 293130 538852 293164
rect 539828 293130 539844 293164
rect 540072 293130 540088 293164
rect 541064 293130 541080 293164
rect 541308 293130 541324 293164
rect 542300 293130 542316 293164
rect 542544 293130 542560 293164
rect 543536 293130 543552 293164
rect 543780 293130 543796 293164
rect 544772 293130 544788 293164
rect 536287 293102 536321 293118
rect 536287 293018 536321 293034
rect 537415 293102 537449 293118
rect 537415 293018 537449 293034
rect 537523 293102 537557 293118
rect 537523 293018 537557 293034
rect 538651 293102 538685 293118
rect 538651 293018 538685 293034
rect 538759 293102 538793 293118
rect 538759 293018 538793 293034
rect 539887 293102 539921 293118
rect 539887 293018 539921 293034
rect 539995 293102 540029 293118
rect 539995 293018 540029 293034
rect 541123 293102 541157 293118
rect 541123 293018 541157 293034
rect 541231 293102 541265 293118
rect 541231 293018 541265 293034
rect 542359 293102 542393 293118
rect 542359 293018 542393 293034
rect 542467 293102 542501 293118
rect 542467 293018 542501 293034
rect 543595 293102 543629 293118
rect 543595 293018 543629 293034
rect 543703 293102 543737 293118
rect 543703 293018 543737 293034
rect 544831 293102 544865 293118
rect 544831 293018 544865 293034
rect 536364 292972 536380 293006
rect 537356 292972 537372 293006
rect 537600 292972 537616 293006
rect 538592 292972 538608 293006
rect 538836 292972 538852 293006
rect 539828 292972 539844 293006
rect 540072 292972 540088 293006
rect 541064 292972 541080 293006
rect 541308 292972 541324 293006
rect 542300 292972 542316 293006
rect 542544 292972 542560 293006
rect 543536 292972 543552 293006
rect 543780 292972 543796 293006
rect 544772 292972 544788 293006
rect 536185 292892 536219 292954
rect 544933 292892 544967 292954
rect 536185 292858 536281 292892
rect 544871 292858 544967 292892
rect 536185 292664 536281 292698
rect 544871 292664 544967 292698
rect 536185 292602 536219 292664
rect 544933 292602 544967 292664
rect 536364 292550 536380 292584
rect 537356 292550 537372 292584
rect 537600 292550 537616 292584
rect 538592 292550 538608 292584
rect 538836 292550 538852 292584
rect 539828 292550 539844 292584
rect 540072 292550 540088 292584
rect 541064 292550 541080 292584
rect 541308 292550 541324 292584
rect 542300 292550 542316 292584
rect 542544 292550 542560 292584
rect 543536 292550 543552 292584
rect 543780 292550 543796 292584
rect 544772 292550 544788 292584
rect 536287 292522 536321 292538
rect 536287 292438 536321 292454
rect 537415 292522 537449 292538
rect 537415 292438 537449 292454
rect 537523 292522 537557 292538
rect 537523 292438 537557 292454
rect 538651 292522 538685 292538
rect 538651 292438 538685 292454
rect 538759 292522 538793 292538
rect 538759 292438 538793 292454
rect 539887 292522 539921 292538
rect 539887 292438 539921 292454
rect 539995 292522 540029 292538
rect 539995 292438 540029 292454
rect 541123 292522 541157 292538
rect 541123 292438 541157 292454
rect 541231 292522 541265 292538
rect 541231 292438 541265 292454
rect 542359 292522 542393 292538
rect 542359 292438 542393 292454
rect 542467 292522 542501 292538
rect 542467 292438 542501 292454
rect 543595 292522 543629 292538
rect 543595 292438 543629 292454
rect 543703 292522 543737 292538
rect 543703 292438 543737 292454
rect 544831 292522 544865 292538
rect 544831 292438 544865 292454
rect 536364 292392 536380 292426
rect 537356 292392 537372 292426
rect 537600 292392 537616 292426
rect 538592 292392 538608 292426
rect 538836 292392 538852 292426
rect 539828 292392 539844 292426
rect 540072 292392 540088 292426
rect 541064 292392 541080 292426
rect 541308 292392 541324 292426
rect 542300 292392 542316 292426
rect 542544 292392 542560 292426
rect 543536 292392 543552 292426
rect 543780 292392 543796 292426
rect 544772 292392 544788 292426
rect 536185 292312 536219 292374
rect 544933 292312 544967 292374
rect 536185 292278 536281 292312
rect 544871 292278 544967 292312
rect 537959 292222 538249 292278
rect 537959 292142 537979 292222
rect 538069 292142 538139 292222
rect 538229 292142 538249 292222
rect 537959 292118 538249 292142
rect 540439 292212 540729 292278
rect 540439 292142 540459 292212
rect 540539 292142 540629 292212
rect 540709 292142 540729 292212
rect 540439 292118 540729 292142
rect 542899 292212 543189 292278
rect 542899 292142 542919 292212
rect 542999 292142 543089 292212
rect 543169 292142 543189 292212
rect 542899 292118 543189 292142
rect 530592 292067 530688 292101
rect 533620 292067 533716 292101
rect 530592 292005 530626 292067
rect 533682 292005 533716 292067
rect 530592 290729 530626 290791
rect 536185 292084 536281 292118
rect 544871 292084 544967 292118
rect 536185 292022 536219 292084
rect 544933 292022 544967 292084
rect 536364 291970 536380 292004
rect 537356 291970 537372 292004
rect 537600 291970 537616 292004
rect 538592 291970 538608 292004
rect 538836 291970 538852 292004
rect 539828 291970 539844 292004
rect 540072 291970 540088 292004
rect 541064 291970 541080 292004
rect 541308 291970 541324 292004
rect 542300 291970 542316 292004
rect 542544 291970 542560 292004
rect 543536 291970 543552 292004
rect 543780 291970 543796 292004
rect 544772 291970 544788 292004
rect 536287 291942 536321 291958
rect 536287 291858 536321 291874
rect 537415 291942 537449 291958
rect 537415 291858 537449 291874
rect 537523 291942 537557 291958
rect 537523 291858 537557 291874
rect 538651 291942 538685 291958
rect 538651 291858 538685 291874
rect 538759 291942 538793 291958
rect 538759 291858 538793 291874
rect 539887 291942 539921 291958
rect 539887 291858 539921 291874
rect 539995 291942 540029 291958
rect 539995 291858 540029 291874
rect 541123 291942 541157 291958
rect 541123 291858 541157 291874
rect 541231 291942 541265 291958
rect 541231 291858 541265 291874
rect 542359 291942 542393 291958
rect 542359 291858 542393 291874
rect 542467 291942 542501 291958
rect 542467 291858 542501 291874
rect 543595 291942 543629 291958
rect 543595 291858 543629 291874
rect 543703 291942 543737 291958
rect 543703 291858 543737 291874
rect 544831 291942 544865 291958
rect 544831 291858 544865 291874
rect 536364 291812 536380 291846
rect 537356 291812 537372 291846
rect 537600 291812 537616 291846
rect 538592 291812 538608 291846
rect 538836 291812 538852 291846
rect 539828 291812 539844 291846
rect 540072 291812 540088 291846
rect 541064 291812 541080 291846
rect 541308 291812 541324 291846
rect 542300 291812 542316 291846
rect 542544 291812 542560 291846
rect 543536 291812 543552 291846
rect 543780 291812 543796 291846
rect 544772 291812 544788 291846
rect 536185 291732 536219 291794
rect 544933 291732 544967 291794
rect 536185 291698 536281 291732
rect 544871 291698 544967 291732
rect 547652 292067 547748 292101
rect 550680 292067 550776 292101
rect 547652 292005 547686 292067
rect 534345 291544 534441 291578
rect 546739 291544 546835 291578
rect 534345 291482 534379 291544
rect 546801 291482 546835 291544
rect 534524 291430 534540 291464
rect 535516 291430 535532 291464
rect 535760 291430 535776 291464
rect 536752 291430 536768 291464
rect 536996 291430 537012 291464
rect 537988 291430 538004 291464
rect 538232 291430 538248 291464
rect 539224 291430 539240 291464
rect 539468 291430 539484 291464
rect 540460 291430 540476 291464
rect 540704 291430 540720 291464
rect 541696 291430 541712 291464
rect 541940 291430 541956 291464
rect 542932 291430 542948 291464
rect 543176 291430 543192 291464
rect 544168 291430 544184 291464
rect 544412 291430 544428 291464
rect 545404 291430 545420 291464
rect 545648 291430 545664 291464
rect 546640 291430 546656 291464
rect 534447 291402 534481 291418
rect 534447 291318 534481 291334
rect 535575 291402 535609 291418
rect 535575 291318 535609 291334
rect 535683 291402 535717 291418
rect 535683 291318 535717 291334
rect 536811 291402 536845 291418
rect 536811 291318 536845 291334
rect 536919 291402 536953 291418
rect 536919 291318 536953 291334
rect 538047 291402 538081 291418
rect 538047 291318 538081 291334
rect 538155 291402 538189 291418
rect 538155 291318 538189 291334
rect 539283 291402 539317 291418
rect 539283 291318 539317 291334
rect 539391 291402 539425 291418
rect 539391 291318 539425 291334
rect 540519 291402 540553 291418
rect 540519 291318 540553 291334
rect 540627 291402 540661 291418
rect 540627 291318 540661 291334
rect 541755 291402 541789 291418
rect 541755 291318 541789 291334
rect 541863 291402 541897 291418
rect 541863 291318 541897 291334
rect 542991 291402 543025 291418
rect 542991 291318 543025 291334
rect 543099 291402 543133 291418
rect 543099 291318 543133 291334
rect 544227 291402 544261 291418
rect 544227 291318 544261 291334
rect 544335 291402 544369 291418
rect 544335 291318 544369 291334
rect 545463 291402 545497 291418
rect 545463 291318 545497 291334
rect 545571 291402 545605 291418
rect 545571 291318 545605 291334
rect 546699 291402 546733 291418
rect 546699 291318 546733 291334
rect 534524 291272 534540 291306
rect 535516 291272 535532 291306
rect 535760 291272 535776 291306
rect 536752 291272 536768 291306
rect 536996 291272 537012 291306
rect 537988 291272 538004 291306
rect 538232 291272 538248 291306
rect 539224 291272 539240 291306
rect 539468 291272 539484 291306
rect 540460 291272 540476 291306
rect 540704 291272 540720 291306
rect 541696 291272 541712 291306
rect 541940 291272 541956 291306
rect 542932 291272 542948 291306
rect 543176 291272 543192 291306
rect 544168 291272 544184 291306
rect 544412 291272 544428 291306
rect 545404 291272 545420 291306
rect 545648 291272 545664 291306
rect 546640 291272 546656 291306
rect 534345 291192 534379 291254
rect 546801 291192 546835 291254
rect 534345 291158 534441 291192
rect 546739 291158 546835 291192
rect 536099 291142 536409 291158
rect 536099 291062 536119 291142
rect 536209 291062 536299 291142
rect 536389 291062 536409 291142
rect 536099 291038 536409 291062
rect 538629 291142 538919 291158
rect 538629 291062 538649 291142
rect 538739 291062 538809 291142
rect 538899 291062 538919 291142
rect 538629 291038 538919 291062
rect 541099 291142 541389 291158
rect 541099 291062 541119 291142
rect 541209 291062 541279 291142
rect 541369 291062 541389 291142
rect 541099 291038 541389 291062
rect 543549 291142 543839 291158
rect 543549 291062 543569 291142
rect 543659 291062 543729 291142
rect 543819 291062 543839 291142
rect 543549 291038 543839 291062
rect 546049 291142 546339 291158
rect 546049 291062 546069 291142
rect 546159 291062 546229 291142
rect 546319 291062 546339 291142
rect 546049 291038 546339 291062
rect 531779 290729 531869 290742
rect 533682 290729 533716 290791
rect 530592 290695 530688 290729
rect 533620 290695 533716 290729
rect 534345 291004 534441 291038
rect 546739 291004 546835 291038
rect 534345 290942 534379 291004
rect 546801 290942 546835 291004
rect 534524 290890 534540 290924
rect 535516 290890 535532 290924
rect 535760 290890 535776 290924
rect 536752 290890 536768 290924
rect 536996 290890 537012 290924
rect 537988 290890 538004 290924
rect 538232 290890 538248 290924
rect 539224 290890 539240 290924
rect 539468 290890 539484 290924
rect 540460 290890 540476 290924
rect 540704 290890 540720 290924
rect 541696 290890 541712 290924
rect 541940 290890 541956 290924
rect 542932 290890 542948 290924
rect 543176 290890 543192 290924
rect 544168 290890 544184 290924
rect 544412 290890 544428 290924
rect 545404 290890 545420 290924
rect 545648 290890 545664 290924
rect 546640 290890 546656 290924
rect 534447 290862 534481 290878
rect 534447 290778 534481 290794
rect 535575 290862 535609 290878
rect 535575 290778 535609 290794
rect 535683 290862 535717 290878
rect 535683 290778 535717 290794
rect 536811 290862 536845 290878
rect 536811 290778 536845 290794
rect 536919 290862 536953 290878
rect 536919 290778 536953 290794
rect 538047 290862 538081 290878
rect 538047 290778 538081 290794
rect 538155 290862 538189 290878
rect 538155 290778 538189 290794
rect 539283 290862 539317 290878
rect 539283 290778 539317 290794
rect 539391 290862 539425 290878
rect 539391 290778 539425 290794
rect 540519 290862 540553 290878
rect 540519 290778 540553 290794
rect 540627 290862 540661 290878
rect 540627 290778 540661 290794
rect 541755 290862 541789 290878
rect 541755 290778 541789 290794
rect 541863 290862 541897 290878
rect 541863 290778 541897 290794
rect 542991 290862 543025 290878
rect 542991 290778 543025 290794
rect 543099 290862 543133 290878
rect 543099 290778 543133 290794
rect 544227 290862 544261 290878
rect 544227 290778 544261 290794
rect 544335 290862 544369 290878
rect 544335 290778 544369 290794
rect 545463 290862 545497 290878
rect 545463 290778 545497 290794
rect 545571 290862 545605 290878
rect 545571 290778 545605 290794
rect 546699 290862 546733 290878
rect 546699 290778 546733 290794
rect 534524 290732 534540 290766
rect 535516 290732 535532 290766
rect 535760 290732 535776 290766
rect 536752 290732 536768 290766
rect 536996 290732 537012 290766
rect 537988 290732 538004 290766
rect 538232 290732 538248 290766
rect 539224 290732 539240 290766
rect 539468 290732 539484 290766
rect 540460 290732 540476 290766
rect 540704 290732 540720 290766
rect 541696 290732 541712 290766
rect 541940 290732 541956 290766
rect 542932 290732 542948 290766
rect 543176 290732 543192 290766
rect 544168 290732 544184 290766
rect 544412 290732 544428 290766
rect 545404 290732 545420 290766
rect 545648 290732 545664 290766
rect 546640 290732 546656 290766
rect 531779 290631 531869 290695
rect 534345 290652 534379 290714
rect 546801 290652 546835 290714
rect 550742 292005 550776 292067
rect 547652 290729 547686 290791
rect 550742 290729 550776 290791
rect 547652 290695 547748 290729
rect 550680 290695 550776 290729
rect 530592 290597 530688 290631
rect 533620 290597 533716 290631
rect 534345 290618 534441 290652
rect 546739 290618 546835 290652
rect 549029 290631 549169 290695
rect 530592 290535 530626 290597
rect 533682 290535 533716 290597
rect 530592 289259 530626 289321
rect 547652 290597 547748 290631
rect 550680 290597 550776 290631
rect 547652 290535 547686 290597
rect 534345 290464 534441 290498
rect 546739 290464 546835 290498
rect 534345 290402 534379 290464
rect 546801 290402 546835 290464
rect 534524 290350 534540 290384
rect 535516 290350 535532 290384
rect 535760 290350 535776 290384
rect 536752 290350 536768 290384
rect 536996 290350 537012 290384
rect 537988 290350 538004 290384
rect 538232 290350 538248 290384
rect 539224 290350 539240 290384
rect 539468 290350 539484 290384
rect 540460 290350 540476 290384
rect 540704 290350 540720 290384
rect 541696 290350 541712 290384
rect 541940 290350 541956 290384
rect 542932 290350 542948 290384
rect 543176 290350 543192 290384
rect 544168 290350 544184 290384
rect 544412 290350 544428 290384
rect 545404 290350 545420 290384
rect 545648 290350 545664 290384
rect 546640 290350 546656 290384
rect 534447 290322 534481 290338
rect 534447 290238 534481 290254
rect 535575 290322 535609 290338
rect 535575 290238 535609 290254
rect 535683 290322 535717 290338
rect 535683 290238 535717 290254
rect 536811 290322 536845 290338
rect 536811 290238 536845 290254
rect 536919 290322 536953 290338
rect 536919 290238 536953 290254
rect 538047 290322 538081 290338
rect 538047 290238 538081 290254
rect 538155 290322 538189 290338
rect 538155 290238 538189 290254
rect 539283 290322 539317 290338
rect 539283 290238 539317 290254
rect 539391 290322 539425 290338
rect 539391 290238 539425 290254
rect 540519 290322 540553 290338
rect 540519 290238 540553 290254
rect 540627 290322 540661 290338
rect 540627 290238 540661 290254
rect 541755 290322 541789 290338
rect 541755 290238 541789 290254
rect 541863 290322 541897 290338
rect 541863 290238 541897 290254
rect 542991 290322 543025 290338
rect 542991 290238 543025 290254
rect 543099 290322 543133 290338
rect 543099 290238 543133 290254
rect 544227 290322 544261 290338
rect 544227 290238 544261 290254
rect 544335 290322 544369 290338
rect 544335 290238 544369 290254
rect 545463 290322 545497 290338
rect 545463 290238 545497 290254
rect 545571 290322 545605 290338
rect 545571 290238 545605 290254
rect 546699 290322 546733 290338
rect 546699 290238 546733 290254
rect 534524 290192 534540 290226
rect 535516 290192 535532 290226
rect 535760 290192 535776 290226
rect 536752 290192 536768 290226
rect 536996 290192 537012 290226
rect 537988 290192 538004 290226
rect 538232 290192 538248 290226
rect 539224 290192 539240 290226
rect 539468 290192 539484 290226
rect 540460 290192 540476 290226
rect 540704 290192 540720 290226
rect 541696 290192 541712 290226
rect 541940 290192 541956 290226
rect 542932 290192 542948 290226
rect 543176 290192 543192 290226
rect 544168 290192 544184 290226
rect 544412 290192 544428 290226
rect 545404 290192 545420 290226
rect 545648 290192 545664 290226
rect 546640 290192 546656 290226
rect 534345 290112 534379 290174
rect 546801 290112 546835 290174
rect 534345 290078 534441 290112
rect 546739 290078 546835 290112
rect 536099 290072 536409 290078
rect 536099 290062 536299 290072
rect 536099 289982 536119 290062
rect 536209 289992 536299 290062
rect 536389 289992 536409 290072
rect 536209 289982 536409 289992
rect 536099 289958 536409 289982
rect 538629 290062 538919 290078
rect 538629 289982 538649 290062
rect 538739 289982 538809 290062
rect 538899 289982 538919 290062
rect 538629 289958 538919 289982
rect 541099 290062 541389 290078
rect 541099 289982 541119 290062
rect 541209 289982 541279 290062
rect 541369 289982 541389 290062
rect 541099 289958 541389 289982
rect 543549 290062 543839 290078
rect 543549 289982 543569 290062
rect 543659 289982 543729 290062
rect 543819 289982 543839 290062
rect 543549 289958 543839 289982
rect 546049 290062 546339 290078
rect 546049 289982 546069 290062
rect 546159 289982 546229 290062
rect 546319 289982 546339 290062
rect 546049 289958 546339 289982
rect 534345 289924 534441 289958
rect 546739 289924 546835 289958
rect 534345 289862 534379 289924
rect 546801 289862 546835 289924
rect 534524 289810 534540 289844
rect 535516 289810 535532 289844
rect 535760 289810 535776 289844
rect 536752 289810 536768 289844
rect 536996 289810 537012 289844
rect 537988 289810 538004 289844
rect 538232 289810 538248 289844
rect 539224 289810 539240 289844
rect 539468 289810 539484 289844
rect 540460 289810 540476 289844
rect 540704 289810 540720 289844
rect 541696 289810 541712 289844
rect 541940 289810 541956 289844
rect 542932 289810 542948 289844
rect 543176 289810 543192 289844
rect 544168 289810 544184 289844
rect 544412 289810 544428 289844
rect 545404 289810 545420 289844
rect 545648 289810 545664 289844
rect 546640 289810 546656 289844
rect 534447 289782 534481 289798
rect 534447 289698 534481 289714
rect 535575 289782 535609 289798
rect 535575 289698 535609 289714
rect 535683 289782 535717 289798
rect 535683 289698 535717 289714
rect 536811 289782 536845 289798
rect 536811 289698 536845 289714
rect 536919 289782 536953 289798
rect 536919 289698 536953 289714
rect 538047 289782 538081 289798
rect 538047 289698 538081 289714
rect 538155 289782 538189 289798
rect 538155 289698 538189 289714
rect 539283 289782 539317 289798
rect 539283 289698 539317 289714
rect 539391 289782 539425 289798
rect 539391 289698 539425 289714
rect 540519 289782 540553 289798
rect 540519 289698 540553 289714
rect 540627 289782 540661 289798
rect 540627 289698 540661 289714
rect 541755 289782 541789 289798
rect 541755 289698 541789 289714
rect 541863 289782 541897 289798
rect 541863 289698 541897 289714
rect 542991 289782 543025 289798
rect 542991 289698 543025 289714
rect 543099 289782 543133 289798
rect 543099 289698 543133 289714
rect 544227 289782 544261 289798
rect 544227 289698 544261 289714
rect 544335 289782 544369 289798
rect 544335 289698 544369 289714
rect 545463 289782 545497 289798
rect 545463 289698 545497 289714
rect 545571 289782 545605 289798
rect 545571 289698 545605 289714
rect 546699 289782 546733 289798
rect 546699 289698 546733 289714
rect 534524 289652 534540 289686
rect 535516 289652 535532 289686
rect 535760 289652 535776 289686
rect 536752 289652 536768 289686
rect 536996 289652 537012 289686
rect 537988 289652 538004 289686
rect 538232 289652 538248 289686
rect 539224 289652 539240 289686
rect 539468 289652 539484 289686
rect 540460 289652 540476 289686
rect 540704 289652 540720 289686
rect 541696 289652 541712 289686
rect 541940 289652 541956 289686
rect 542932 289652 542948 289686
rect 543176 289652 543192 289686
rect 544168 289652 544184 289686
rect 544412 289652 544428 289686
rect 545404 289652 545420 289686
rect 545648 289652 545664 289686
rect 546640 289652 546656 289686
rect 534345 289572 534379 289634
rect 546801 289572 546835 289634
rect 534345 289538 534441 289572
rect 546739 289538 546835 289572
rect 533682 289259 533716 289321
rect 530592 289225 530688 289259
rect 533620 289225 533716 289259
rect 550742 290535 550776 290597
rect 547652 289259 547686 289321
rect 550742 289259 550776 289321
rect 547652 289225 547748 289259
rect 550680 289225 550776 289259
rect 536285 289144 536381 289178
rect 544845 289144 544941 289178
rect 536285 289082 536319 289144
rect 544907 289082 544941 289144
rect 536455 289030 536471 289064
rect 537447 289030 537463 289064
rect 537673 289030 537689 289064
rect 538665 289030 538681 289064
rect 538891 289030 538907 289064
rect 539883 289030 539899 289064
rect 540109 289030 540125 289064
rect 541101 289030 541117 289064
rect 541327 289030 541343 289064
rect 542319 289030 542335 289064
rect 542545 289030 542561 289064
rect 543537 289030 543553 289064
rect 543763 289030 543779 289064
rect 544755 289030 544771 289064
rect 536387 289002 536421 289018
rect 536387 288918 536421 288934
rect 537497 289002 537531 289018
rect 537497 288918 537531 288934
rect 537605 289002 537639 289018
rect 537605 288918 537639 288934
rect 538715 289002 538749 289018
rect 538715 288918 538749 288934
rect 538823 289002 538857 289018
rect 538823 288918 538857 288934
rect 539933 289002 539967 289018
rect 539933 288918 539967 288934
rect 540041 289002 540075 289018
rect 540041 288918 540075 288934
rect 541151 289002 541185 289018
rect 541151 288918 541185 288934
rect 541259 289002 541293 289018
rect 541259 288918 541293 288934
rect 542369 289002 542403 289018
rect 542369 288918 542403 288934
rect 542477 289002 542511 289018
rect 542477 288918 542511 288934
rect 543587 289002 543621 289018
rect 543587 288918 543621 288934
rect 543695 289002 543729 289018
rect 543695 288918 543729 288934
rect 544805 289002 544839 289018
rect 544805 288918 544839 288934
rect 536455 288872 536471 288906
rect 537447 288872 537463 288906
rect 537673 288872 537689 288906
rect 538665 288872 538681 288906
rect 538891 288872 538907 288906
rect 539883 288872 539899 288906
rect 540109 288872 540125 288906
rect 541101 288872 541117 288906
rect 541327 288872 541343 288906
rect 542319 288872 542335 288906
rect 542545 288872 542561 288906
rect 543537 288872 543553 288906
rect 543763 288872 543779 288906
rect 544755 288872 544771 288906
rect 536285 288792 536319 288854
rect 544907 288792 544941 288854
rect 536285 288758 536381 288792
rect 544845 288758 544941 288792
rect 568116 288824 568212 288858
rect 578368 288824 578464 288858
rect 568116 288762 568150 288824
rect 536285 288644 536381 288678
rect 544845 288644 544941 288678
rect 536285 288582 536319 288644
rect 544907 288582 544941 288644
rect 536455 288530 536471 288564
rect 537447 288530 537463 288564
rect 537673 288530 537689 288564
rect 538665 288530 538681 288564
rect 538891 288530 538907 288564
rect 539883 288530 539899 288564
rect 540109 288530 540125 288564
rect 541101 288530 541117 288564
rect 541327 288530 541343 288564
rect 542319 288530 542335 288564
rect 542545 288530 542561 288564
rect 543537 288530 543553 288564
rect 543763 288530 543779 288564
rect 544755 288530 544771 288564
rect 536387 288502 536421 288518
rect 536387 288418 536421 288434
rect 537497 288502 537531 288518
rect 537497 288418 537531 288434
rect 537605 288502 537639 288518
rect 537605 288418 537639 288434
rect 538715 288502 538749 288518
rect 538715 288418 538749 288434
rect 538823 288502 538857 288518
rect 538823 288418 538857 288434
rect 539933 288502 539967 288518
rect 539933 288418 539967 288434
rect 540041 288502 540075 288518
rect 540041 288418 540075 288434
rect 541151 288502 541185 288518
rect 541151 288418 541185 288434
rect 541259 288502 541293 288518
rect 541259 288418 541293 288434
rect 542369 288502 542403 288518
rect 542369 288418 542403 288434
rect 542477 288502 542511 288518
rect 542477 288418 542511 288434
rect 543587 288502 543621 288518
rect 543587 288418 543621 288434
rect 543695 288502 543729 288518
rect 543695 288418 543729 288434
rect 544805 288502 544839 288518
rect 544805 288418 544839 288434
rect 536455 288372 536471 288406
rect 537447 288372 537463 288406
rect 537673 288372 537689 288406
rect 538665 288372 538681 288406
rect 538891 288372 538907 288406
rect 539883 288372 539899 288406
rect 540109 288372 540125 288406
rect 541101 288372 541117 288406
rect 541327 288372 541343 288406
rect 542319 288372 542335 288406
rect 542545 288372 542561 288406
rect 543537 288372 543553 288406
rect 543763 288372 543779 288406
rect 544755 288372 544771 288406
rect 536285 288292 536319 288354
rect 544907 288292 544941 288354
rect 536285 288258 536381 288292
rect 544845 288258 544941 288292
rect 568218 288695 568252 288711
rect 568286 288710 568302 288744
rect 578278 288710 578294 288744
rect 568218 288645 568252 288661
rect 568286 288612 568302 288646
rect 578278 288612 578294 288646
rect 578328 288597 578362 288613
rect 536845 288144 536941 288178
rect 544187 288144 544283 288178
rect 536845 288082 536879 288144
rect 544249 288082 544283 288144
rect 537015 288030 537031 288064
rect 538007 288030 538023 288064
rect 538233 288030 538249 288064
rect 539225 288030 539241 288064
rect 539451 288030 539467 288064
rect 540443 288030 540459 288064
rect 540669 288030 540685 288064
rect 541661 288030 541677 288064
rect 541887 288030 541903 288064
rect 542879 288030 542895 288064
rect 543105 288030 543121 288064
rect 544097 288030 544113 288064
rect 536947 288002 536981 288018
rect 536947 287818 536981 287834
rect 538057 288002 538091 288018
rect 538057 287818 538091 287834
rect 538165 288002 538199 288018
rect 538165 287818 538199 287834
rect 539275 288002 539309 288018
rect 539275 287818 539309 287834
rect 539383 288002 539417 288018
rect 539383 287818 539417 287834
rect 540493 288002 540527 288018
rect 540493 287818 540527 287834
rect 540601 288002 540635 288018
rect 540601 287818 540635 287834
rect 541711 288002 541745 288018
rect 541711 287818 541745 287834
rect 541819 288002 541853 288018
rect 541819 287818 541853 287834
rect 542929 288002 542963 288018
rect 542929 287818 542963 287834
rect 543037 288002 543071 288018
rect 543037 287818 543071 287834
rect 544147 288002 544181 288018
rect 544147 287818 544181 287834
rect 537015 287772 537031 287806
rect 538007 287772 538023 287806
rect 538233 287772 538249 287806
rect 539225 287772 539241 287806
rect 539451 287772 539467 287806
rect 540443 287772 540459 287806
rect 540669 287772 540685 287806
rect 541661 287772 541677 287806
rect 541887 287772 541903 287806
rect 542879 287772 542895 287806
rect 543105 287772 543121 287806
rect 544097 287772 544113 287806
rect 536845 287692 536879 287754
rect 544249 287692 544283 287754
rect 536845 287658 536941 287692
rect 544187 287658 544283 287692
rect 568218 288499 568252 288515
rect 568286 288514 568302 288548
rect 578278 288514 578294 288548
rect 578328 288547 578362 288563
rect 568218 288449 568252 288465
rect 568286 288416 568302 288450
rect 578278 288416 578294 288450
rect 578328 288401 578362 288417
rect 568218 288303 568252 288319
rect 568286 288318 568302 288352
rect 578278 288318 578294 288352
rect 578328 288351 578362 288367
rect 568218 288253 568252 288269
rect 568286 288220 568302 288254
rect 578278 288220 578294 288254
rect 578328 288205 578362 288221
rect 568218 288107 568252 288123
rect 568286 288122 568302 288156
rect 578278 288122 578294 288156
rect 578328 288155 578362 288171
rect 568218 288057 568252 288073
rect 568286 288024 568302 288058
rect 578278 288024 578294 288058
rect 578328 288009 578362 288025
rect 568218 287911 568252 287927
rect 568286 287926 568302 287960
rect 578278 287926 578294 287960
rect 578328 287959 578362 287975
rect 568218 287861 568252 287877
rect 568286 287828 568302 287862
rect 578278 287828 578294 287862
rect 578328 287813 578362 287829
rect 568286 287730 568302 287764
rect 578278 287730 578294 287764
rect 578328 287763 578362 287779
rect 537539 287652 537709 287658
rect 537539 287562 537569 287652
rect 537679 287562 537709 287652
rect 537539 287558 537709 287562
rect 542449 287652 542619 287658
rect 542449 287562 542479 287652
rect 542589 287562 542619 287652
rect 568116 287650 568150 287712
rect 578430 287650 578464 288824
rect 568116 287616 568212 287650
rect 578368 287616 578464 287650
rect 542449 287558 542619 287562
rect 536845 287524 536941 287558
rect 544187 287524 544283 287558
rect 536845 287462 536879 287524
rect 544249 287462 544283 287524
rect 537015 287410 537031 287444
rect 538007 287410 538023 287444
rect 538233 287410 538249 287444
rect 539225 287410 539241 287444
rect 539451 287410 539467 287444
rect 540443 287410 540459 287444
rect 540669 287410 540685 287444
rect 541661 287410 541677 287444
rect 541887 287410 541903 287444
rect 542879 287410 542895 287444
rect 543105 287410 543121 287444
rect 544097 287410 544113 287444
rect 536947 287382 536981 287398
rect 536947 287198 536981 287214
rect 538057 287382 538091 287398
rect 538057 287198 538091 287214
rect 538165 287382 538199 287398
rect 538165 287198 538199 287214
rect 539275 287382 539309 287398
rect 539275 287198 539309 287214
rect 539383 287382 539417 287398
rect 539383 287198 539417 287214
rect 540493 287382 540527 287398
rect 540493 287198 540527 287214
rect 540601 287382 540635 287398
rect 540601 287198 540635 287214
rect 541711 287382 541745 287398
rect 541711 287198 541745 287214
rect 541819 287382 541853 287398
rect 541819 287198 541853 287214
rect 542929 287382 542963 287398
rect 542929 287198 542963 287214
rect 543037 287382 543071 287398
rect 543037 287198 543071 287214
rect 544147 287382 544181 287398
rect 544147 287198 544181 287214
rect 537015 287152 537031 287186
rect 538007 287152 538023 287186
rect 538233 287152 538249 287186
rect 539225 287152 539241 287186
rect 539451 287152 539467 287186
rect 540443 287152 540459 287186
rect 540669 287152 540685 287186
rect 541661 287152 541677 287186
rect 541887 287152 541903 287186
rect 542879 287152 542895 287186
rect 543105 287152 543121 287186
rect 544097 287152 544113 287186
rect 536845 287072 536879 287134
rect 544249 287072 544283 287134
rect 536845 287038 536941 287072
rect 544187 287038 544283 287072
rect 536285 286924 536381 286958
rect 544845 286924 544941 286958
rect 536285 286862 536319 286924
rect 544907 286862 544941 286924
rect 536455 286810 536471 286844
rect 537447 286810 537463 286844
rect 537673 286810 537689 286844
rect 538665 286810 538681 286844
rect 538891 286810 538907 286844
rect 539883 286810 539899 286844
rect 540109 286810 540125 286844
rect 541101 286810 541117 286844
rect 541327 286810 541343 286844
rect 542319 286810 542335 286844
rect 542545 286810 542561 286844
rect 543537 286810 543553 286844
rect 543763 286810 543779 286844
rect 544755 286810 544771 286844
rect 536387 286782 536421 286798
rect 536387 286598 536421 286614
rect 537497 286782 537531 286798
rect 537497 286598 537531 286614
rect 537605 286782 537639 286798
rect 537605 286598 537639 286614
rect 538715 286782 538749 286798
rect 538715 286598 538749 286614
rect 538823 286782 538857 286798
rect 538823 286598 538857 286614
rect 539933 286782 539967 286798
rect 539933 286598 539967 286614
rect 540041 286782 540075 286798
rect 540041 286598 540075 286614
rect 541151 286782 541185 286798
rect 541151 286598 541185 286614
rect 541259 286782 541293 286798
rect 541259 286598 541293 286614
rect 542369 286782 542403 286798
rect 542369 286598 542403 286614
rect 542477 286782 542511 286798
rect 542477 286598 542511 286614
rect 543587 286782 543621 286798
rect 543587 286598 543621 286614
rect 543695 286782 543729 286798
rect 543695 286598 543729 286614
rect 544805 286782 544839 286798
rect 544805 286598 544839 286614
rect 536455 286552 536471 286586
rect 537447 286552 537463 286586
rect 537673 286552 537689 286586
rect 538665 286552 538681 286586
rect 538891 286552 538907 286586
rect 539883 286552 539899 286586
rect 540109 286552 540125 286586
rect 541101 286552 541117 286586
rect 541327 286552 541343 286586
rect 542319 286552 542335 286586
rect 542545 286552 542561 286586
rect 543537 286552 543553 286586
rect 543763 286552 543779 286586
rect 544755 286552 544771 286586
rect 536285 286472 536319 286534
rect 544907 286472 544941 286534
rect 536285 286438 536381 286472
rect 544845 286438 544941 286472
rect 536285 286324 536381 286358
rect 544845 286324 544941 286358
rect 536285 286262 536319 286324
rect 544907 286262 544941 286324
rect 536455 286210 536471 286244
rect 537447 286210 537463 286244
rect 537673 286210 537689 286244
rect 538665 286210 538681 286244
rect 538891 286210 538907 286244
rect 539883 286210 539899 286244
rect 540109 286210 540125 286244
rect 541101 286210 541117 286244
rect 541327 286210 541343 286244
rect 542319 286210 542335 286244
rect 542545 286210 542561 286244
rect 543537 286210 543553 286244
rect 543763 286210 543779 286244
rect 544755 286210 544771 286244
rect 536387 286182 536421 286198
rect 536387 285998 536421 286014
rect 537497 286182 537531 286198
rect 537497 285998 537531 286014
rect 537605 286182 537639 286198
rect 537605 285998 537639 286014
rect 538715 286182 538749 286198
rect 538715 285998 538749 286014
rect 538823 286182 538857 286198
rect 538823 285998 538857 286014
rect 539933 286182 539967 286198
rect 539933 285998 539967 286014
rect 540041 286182 540075 286198
rect 540041 285998 540075 286014
rect 541151 286182 541185 286198
rect 541151 285998 541185 286014
rect 541259 286182 541293 286198
rect 541259 285998 541293 286014
rect 542369 286182 542403 286198
rect 542369 285998 542403 286014
rect 542477 286182 542511 286198
rect 542477 285998 542511 286014
rect 543587 286182 543621 286198
rect 543587 285998 543621 286014
rect 543695 286182 543729 286198
rect 543695 285998 543729 286014
rect 544805 286182 544839 286198
rect 544805 285998 544839 286014
rect 536455 285952 536471 285986
rect 537447 285952 537463 285986
rect 537673 285952 537689 285986
rect 538665 285952 538681 285986
rect 538891 285952 538907 285986
rect 539883 285952 539899 285986
rect 540109 285952 540125 285986
rect 541101 285952 541117 285986
rect 541327 285952 541343 285986
rect 542319 285952 542335 285986
rect 542545 285952 542561 285986
rect 543537 285952 543553 285986
rect 543763 285952 543779 285986
rect 544755 285952 544771 285986
rect 536285 285872 536319 285934
rect 544907 285872 544941 285934
rect 536285 285838 536381 285872
rect 544845 285838 544941 285872
rect 536830 285350 536926 285384
rect 544280 285350 544376 285384
rect 536830 285288 536864 285350
rect 544342 285288 544376 285350
rect 537009 285236 537025 285270
rect 538001 285236 538017 285270
rect 538245 285236 538261 285270
rect 539237 285236 539253 285270
rect 539481 285236 539497 285270
rect 540473 285236 540489 285270
rect 540717 285236 540733 285270
rect 541709 285236 541725 285270
rect 541953 285236 541969 285270
rect 542945 285236 542961 285270
rect 543189 285236 543205 285270
rect 544181 285236 544197 285270
rect 536932 285208 536966 285224
rect 536932 285024 536966 285040
rect 538060 285208 538094 285224
rect 538060 285024 538094 285040
rect 538168 285208 538202 285224
rect 538168 285024 538202 285040
rect 539296 285208 539330 285224
rect 539296 285024 539330 285040
rect 539404 285208 539438 285224
rect 539404 285024 539438 285040
rect 540532 285208 540566 285224
rect 540532 285024 540566 285040
rect 540640 285208 540674 285224
rect 540640 285024 540674 285040
rect 541768 285208 541802 285224
rect 541768 285024 541802 285040
rect 541876 285208 541910 285224
rect 541876 285024 541910 285040
rect 543004 285208 543038 285224
rect 543004 285024 543038 285040
rect 543112 285208 543146 285224
rect 543112 285024 543146 285040
rect 544240 285208 544274 285224
rect 544240 285024 544274 285040
rect 537009 284978 537025 285012
rect 538001 284978 538017 285012
rect 538245 284978 538261 285012
rect 539237 284978 539253 285012
rect 539481 284978 539497 285012
rect 540473 284978 540489 285012
rect 540717 284978 540733 285012
rect 541709 284978 541725 285012
rect 541953 284978 541969 285012
rect 542945 284978 542961 285012
rect 543189 284978 543205 285012
rect 544181 284978 544197 285012
rect 536830 284898 536864 284960
rect 544342 284898 544376 284960
rect 536830 284864 536926 284898
rect 544280 284864 544376 284898
rect 536830 284760 536926 284794
rect 544280 284760 544376 284794
rect 536830 284698 536864 284760
rect 544342 284698 544376 284760
rect 537009 284646 537025 284680
rect 538001 284646 538017 284680
rect 538245 284646 538261 284680
rect 539237 284646 539253 284680
rect 539481 284646 539497 284680
rect 540473 284646 540489 284680
rect 540717 284646 540733 284680
rect 541709 284646 541725 284680
rect 541953 284646 541969 284680
rect 542945 284646 542961 284680
rect 543189 284646 543205 284680
rect 544181 284646 544197 284680
rect 536932 284618 536966 284634
rect 536932 284434 536966 284450
rect 538060 284618 538094 284634
rect 538060 284434 538094 284450
rect 538168 284618 538202 284634
rect 538168 284434 538202 284450
rect 539296 284618 539330 284634
rect 539296 284434 539330 284450
rect 539404 284618 539438 284634
rect 539404 284434 539438 284450
rect 540532 284618 540566 284634
rect 540532 284434 540566 284450
rect 540640 284618 540674 284634
rect 540640 284434 540674 284450
rect 541768 284618 541802 284634
rect 541768 284434 541802 284450
rect 541876 284618 541910 284634
rect 541876 284434 541910 284450
rect 543004 284618 543038 284634
rect 543004 284434 543038 284450
rect 543112 284618 543146 284634
rect 543112 284434 543146 284450
rect 544240 284618 544274 284634
rect 544240 284434 544274 284450
rect 537009 284388 537025 284422
rect 538001 284388 538017 284422
rect 538245 284388 538261 284422
rect 539237 284388 539253 284422
rect 539481 284388 539497 284422
rect 540473 284388 540489 284422
rect 540717 284388 540733 284422
rect 541709 284388 541725 284422
rect 541953 284388 541969 284422
rect 542945 284388 542961 284422
rect 543189 284388 543205 284422
rect 544181 284388 544197 284422
rect 536830 284308 536864 284370
rect 544342 284308 544376 284370
rect 536830 284274 536926 284308
rect 544280 284274 544376 284308
rect 539600 283970 539696 284004
rect 541506 283970 541602 284004
rect 539600 283908 539634 283970
rect 541568 283908 541602 283970
rect 539770 283856 539786 283890
rect 540012 283856 540028 283890
rect 540238 283856 540254 283890
rect 540480 283856 540496 283890
rect 540706 283856 540722 283890
rect 540948 283856 540964 283890
rect 541174 283856 541190 283890
rect 541416 283856 541432 283890
rect 539702 283828 539736 283844
rect 539702 283644 539736 283660
rect 540062 283828 540096 283844
rect 540062 283644 540096 283660
rect 540170 283828 540204 283844
rect 540170 283644 540204 283660
rect 540530 283828 540564 283844
rect 540530 283644 540564 283660
rect 540638 283828 540672 283844
rect 540638 283644 540672 283660
rect 540998 283828 541032 283844
rect 540998 283644 541032 283660
rect 541106 283828 541140 283844
rect 541106 283644 541140 283660
rect 541466 283828 541500 283844
rect 541466 283644 541500 283660
rect 539770 283598 539786 283632
rect 540012 283598 540028 283632
rect 540238 283598 540254 283632
rect 540480 283598 540496 283632
rect 540706 283598 540722 283632
rect 540948 283598 540964 283632
rect 541174 283598 541190 283632
rect 541416 283598 541432 283632
rect 539600 283518 539634 283580
rect 541568 283518 541602 283580
rect 539600 283484 539696 283518
rect 541506 283484 541602 283518
rect 539820 283345 539916 283368
rect 541290 283345 541386 283368
rect 539820 283283 539854 283345
rect 541352 283283 541386 283345
rect 539990 283231 540006 283265
rect 540482 283231 540498 283265
rect 540708 283231 540724 283265
rect 541200 283231 541216 283265
rect 539922 283203 539956 283219
rect 539922 283119 539956 283135
rect 540532 283203 540566 283219
rect 540532 283119 540566 283135
rect 540640 283203 540674 283219
rect 540640 283119 540674 283135
rect 541250 283203 541284 283219
rect 541250 283119 541284 283135
rect 539990 283073 540006 283107
rect 540482 283073 540498 283107
rect 540708 283073 540724 283107
rect 541200 283073 541216 283107
rect 539820 282993 539854 283055
rect 541352 282993 541386 283055
rect 539820 282959 539916 282993
rect 541290 282959 541386 282993
rect 536885 282820 536981 282854
rect 544227 282820 544323 282854
rect 536885 282758 536919 282820
rect 544289 282758 544323 282820
rect 537055 282706 537071 282740
rect 538047 282706 538063 282740
rect 538273 282706 538289 282740
rect 539265 282706 539281 282740
rect 539491 282706 539507 282740
rect 540483 282706 540499 282740
rect 540709 282706 540725 282740
rect 541701 282706 541717 282740
rect 541927 282706 541943 282740
rect 542919 282706 542935 282740
rect 543145 282706 543161 282740
rect 544137 282706 544153 282740
rect 536987 282678 537021 282694
rect 536987 282494 537021 282510
rect 538097 282678 538131 282694
rect 538097 282494 538131 282510
rect 538205 282678 538239 282694
rect 538205 282494 538239 282510
rect 539315 282678 539349 282694
rect 539315 282494 539349 282510
rect 539423 282678 539457 282694
rect 539423 282494 539457 282510
rect 540533 282678 540567 282694
rect 540533 282494 540567 282510
rect 540641 282678 540675 282694
rect 540641 282494 540675 282510
rect 541751 282678 541785 282694
rect 541751 282494 541785 282510
rect 541859 282678 541893 282694
rect 541859 282494 541893 282510
rect 542969 282678 543003 282694
rect 542969 282494 543003 282510
rect 543077 282678 543111 282694
rect 543077 282494 543111 282510
rect 544187 282678 544221 282694
rect 544187 282494 544221 282510
rect 537055 282448 537071 282482
rect 538047 282448 538063 282482
rect 538273 282448 538289 282482
rect 539265 282448 539281 282482
rect 539491 282448 539507 282482
rect 540483 282448 540499 282482
rect 540709 282448 540725 282482
rect 541701 282448 541717 282482
rect 541927 282448 541943 282482
rect 542919 282448 542935 282482
rect 543145 282448 543161 282482
rect 544137 282448 544153 282482
rect 536885 282368 536919 282430
rect 544289 282368 544323 282430
rect 536885 282334 536981 282368
rect 544227 282334 544323 282368
rect 568136 281344 568232 281378
rect 578388 281344 578484 281378
rect 568136 281282 568170 281344
rect 537364 281058 537484 281074
rect 537364 280922 537484 280938
rect 543734 281058 543854 281074
rect 543734 280922 543854 280938
rect 568238 281215 568272 281231
rect 568306 281230 568322 281264
rect 578298 281230 578314 281264
rect 568238 281165 568272 281181
rect 568306 281132 568322 281166
rect 578298 281132 578314 281166
rect 578348 281117 578382 281133
rect 568238 281019 568272 281035
rect 568306 281034 568322 281068
rect 578298 281034 578314 281068
rect 578348 281067 578382 281083
rect 568238 280969 568272 280985
rect 568306 280936 568322 280970
rect 578298 280936 578314 280970
rect 578348 280921 578382 280937
rect 568238 280823 568272 280839
rect 568306 280838 568322 280872
rect 578298 280838 578314 280872
rect 578348 280871 578382 280887
rect 568238 280773 568272 280789
rect 568306 280740 568322 280774
rect 578298 280740 578314 280774
rect 578348 280725 578382 280741
rect 568238 280627 568272 280643
rect 568306 280642 568322 280676
rect 578298 280642 578314 280676
rect 578348 280675 578382 280691
rect 568238 280577 568272 280593
rect 568306 280544 568322 280578
rect 578298 280544 578314 280578
rect 578348 280529 578382 280545
rect 568238 280431 568272 280447
rect 568306 280446 568322 280480
rect 578298 280446 578314 280480
rect 578348 280479 578382 280495
rect 568238 280381 568272 280397
rect 568306 280348 568322 280382
rect 578298 280348 578314 280382
rect 578348 280333 578382 280349
rect 568306 280250 568322 280284
rect 578298 280250 578314 280284
rect 578348 280283 578382 280299
rect 568136 280170 568170 280232
rect 578450 280170 578484 281344
rect 568136 280136 568232 280170
rect 578388 280136 578484 280170
rect 11741 279723 11837 279757
rect 13051 279723 13147 279757
rect 11741 279661 11775 279723
rect 13113 279661 13147 279723
rect 13110 277920 13113 278580
rect 11741 276667 11775 276729
rect 13201 279723 13297 279757
rect 14511 279723 14607 279757
rect 13201 279661 13235 279723
rect 13147 277920 13201 278580
rect 13113 276667 13147 276729
rect 11741 276633 11837 276667
rect 13051 276633 13147 276667
rect 14573 279661 14607 279723
rect 537364 278058 537484 278074
rect 13201 276667 13235 276729
rect 537364 277922 537484 277938
rect 543734 278058 543854 278074
rect 543734 277922 543854 277938
rect 14573 276667 14607 276729
rect 13201 276633 13297 276667
rect 14511 276633 14607 276667
rect 12618 275914 12714 275948
rect 13888 275914 13984 275948
rect 12618 275852 12652 275914
rect 13950 275852 13984 275914
rect 31004 275900 31020 276140
rect 31260 275900 31276 276140
rect 32724 275900 32740 276140
rect 32980 275900 32996 276140
rect 34444 275900 34460 276140
rect 34700 275900 34716 276140
rect 35924 275900 35940 276140
rect 36180 275900 36196 276140
rect 37644 275900 37660 276140
rect 37900 275900 37916 276140
rect 39244 275900 39260 276140
rect 39500 275900 39516 276140
rect 40964 275900 40980 276140
rect 41220 275900 41236 276140
rect 42564 275900 42580 276140
rect 42820 275900 42836 276140
rect 44284 275900 44300 276140
rect 44540 275900 44556 276140
rect 12797 275800 12813 275834
rect 13789 275800 13805 275834
rect 12720 275772 12754 275788
rect 12720 275688 12754 275704
rect 13848 275772 13882 275788
rect 13848 275688 13882 275704
rect 12797 275642 12813 275676
rect 13789 275642 13805 275676
rect 12720 275614 12754 275630
rect 12720 275530 12754 275546
rect 13848 275614 13882 275630
rect 13848 275530 13882 275546
rect 12797 275484 12813 275518
rect 13789 275484 13805 275518
rect 12720 275456 12754 275472
rect 12720 275372 12754 275388
rect 13848 275456 13882 275472
rect 13848 275372 13882 275388
rect 12797 275326 12813 275360
rect 13789 275326 13805 275360
rect 12720 275298 12754 275314
rect 12720 275214 12754 275230
rect 13848 275298 13882 275314
rect 13848 275214 13882 275230
rect 12797 275168 12813 275202
rect 13789 275168 13805 275202
rect 12720 275140 12754 275156
rect 12720 275056 12754 275072
rect 13848 275140 13882 275156
rect 13848 275056 13882 275072
rect 12797 275010 12813 275044
rect 13789 275010 13805 275044
rect 12720 274982 12754 274998
rect 12720 274898 12754 274914
rect 13848 274982 13882 274998
rect 13848 274898 13882 274914
rect 12797 274852 12813 274886
rect 13789 274852 13805 274886
rect 12720 274824 12754 274840
rect 12720 274740 12754 274756
rect 13848 274824 13882 274840
rect 13848 274740 13882 274756
rect 12797 274694 12813 274728
rect 13789 274694 13805 274728
rect 12720 274666 12754 274682
rect 12720 274582 12754 274598
rect 13848 274666 13882 274682
rect 13848 274582 13882 274598
rect 12797 274536 12813 274570
rect 13789 274536 13805 274570
rect 12720 274508 12754 274524
rect 12720 274424 12754 274440
rect 13848 274508 13882 274524
rect 13848 274424 13882 274440
rect 12797 274378 12813 274412
rect 13789 274378 13805 274412
rect 12720 274350 12754 274366
rect 12720 274266 12754 274282
rect 13848 274350 13882 274366
rect 13848 274266 13882 274282
rect 537364 275058 537484 275074
rect 537364 274922 537484 274938
rect 543734 275058 543854 275074
rect 543734 274922 543854 274938
rect 21966 274556 22062 274590
rect 23218 274556 23314 274590
rect 21966 274494 22000 274556
rect 12797 274220 12813 274254
rect 13789 274220 13805 274254
rect 12720 274192 12754 274208
rect 12720 274108 12754 274124
rect 13848 274192 13882 274208
rect 13848 274108 13882 274124
rect 12797 274062 12813 274096
rect 13789 274062 13805 274096
rect 12720 274034 12754 274050
rect 12720 273950 12754 273966
rect 13848 274034 13882 274050
rect 13848 273950 13882 273966
rect 12797 273904 12813 273938
rect 13789 273904 13805 273938
rect 12720 273876 12754 273892
rect 12720 273792 12754 273808
rect 13848 273876 13882 273892
rect 13848 273792 13882 273808
rect 12797 273746 12813 273780
rect 13789 273746 13805 273780
rect 12720 273718 12754 273734
rect 12720 273634 12754 273650
rect 13848 273718 13882 273734
rect 13848 273634 13882 273650
rect 12797 273588 12813 273622
rect 13789 273588 13805 273622
rect 12720 273560 12754 273576
rect 12720 273476 12754 273492
rect 13848 273560 13882 273576
rect 13848 273476 13882 273492
rect 12797 273430 12813 273464
rect 13789 273430 13805 273464
rect 12720 273402 12754 273418
rect 12720 273318 12754 273334
rect 13848 273402 13882 273418
rect 13848 273318 13882 273334
rect 12797 273272 12813 273306
rect 13789 273272 13805 273306
rect 12720 273244 12754 273260
rect 12720 273160 12754 273176
rect 13848 273244 13882 273260
rect 13848 273160 13882 273176
rect 12797 273114 12813 273148
rect 13789 273114 13805 273148
rect 12720 273086 12754 273102
rect 12720 273002 12754 273018
rect 13848 273086 13882 273102
rect 13848 273002 13882 273018
rect 12797 272956 12813 272990
rect 13789 272956 13805 272990
rect 12720 272928 12754 272944
rect 12720 272844 12754 272860
rect 13848 272928 13882 272944
rect 13848 272844 13882 272860
rect 12797 272798 12813 272832
rect 13789 272798 13805 272832
rect 12720 272770 12754 272786
rect 12720 272686 12754 272702
rect 13848 272770 13882 272786
rect 13848 272686 13882 272702
rect 12797 272640 12813 272674
rect 13789 272640 13805 272674
rect 12720 272612 12754 272628
rect 12720 272528 12754 272544
rect 13848 272612 13882 272628
rect 13848 272528 13882 272544
rect 12797 272482 12813 272516
rect 13789 272482 13805 272516
rect 12720 272454 12754 272470
rect 12720 272370 12754 272386
rect 13848 272454 13882 272470
rect 13848 272370 13882 272386
rect 12797 272324 12813 272358
rect 13789 272324 13805 272358
rect 12720 272296 12754 272312
rect 12720 272212 12754 272228
rect 13848 272296 13882 272312
rect 13848 272212 13882 272228
rect 12797 272166 12813 272200
rect 13789 272166 13805 272200
rect 12720 272138 12754 272154
rect 12720 272054 12754 272070
rect 13848 272138 13882 272154
rect 13848 272054 13882 272070
rect 12797 272008 12813 272042
rect 13789 272008 13805 272042
rect 12720 271980 12754 271996
rect 12720 271896 12754 271912
rect 13848 271980 13882 271996
rect 13848 271896 13882 271912
rect 12797 271850 12813 271884
rect 13789 271850 13805 271884
rect 12720 271822 12754 271838
rect 12720 271738 12754 271754
rect 13848 271822 13882 271838
rect 13848 271738 13882 271754
rect 12797 271692 12813 271726
rect 13789 271692 13805 271726
rect 12720 271664 12754 271680
rect 12720 271580 12754 271596
rect 13848 271664 13882 271680
rect 13848 271580 13882 271596
rect 12797 271534 12813 271568
rect 13789 271534 13805 271568
rect 12720 271506 12754 271522
rect 12720 271422 12754 271438
rect 13848 271506 13882 271522
rect 13848 271422 13882 271438
rect 12797 271376 12813 271410
rect 13789 271376 13805 271410
rect 12720 271348 12754 271364
rect 12720 271264 12754 271280
rect 13848 271348 13882 271364
rect 13848 271264 13882 271280
rect 12797 271218 12813 271252
rect 13789 271218 13805 271252
rect 12720 271190 12754 271206
rect 12720 271106 12754 271122
rect 13848 271190 13882 271206
rect 13848 271106 13882 271122
rect 12797 271060 12813 271094
rect 13789 271060 13805 271094
rect 12720 271032 12754 271048
rect 12720 270948 12754 270964
rect 13848 271032 13882 271048
rect 13848 270948 13882 270964
rect 12797 270902 12813 270936
rect 13789 270902 13805 270936
rect 12720 270874 12754 270890
rect 12720 270790 12754 270806
rect 13848 270874 13882 270890
rect 13848 270790 13882 270806
rect 12797 270744 12813 270778
rect 13789 270744 13805 270778
rect 12720 270716 12754 270732
rect 12720 270632 12754 270648
rect 13848 270716 13882 270732
rect 13848 270632 13882 270648
rect 12797 270586 12813 270620
rect 13789 270586 13805 270620
rect 12720 270558 12754 270574
rect 12720 270474 12754 270490
rect 13848 270558 13882 270574
rect 13848 270474 13882 270490
rect 12797 270428 12813 270462
rect 13789 270428 13805 270462
rect 12720 270400 12754 270416
rect 12720 270316 12754 270332
rect 13848 270400 13882 270416
rect 13848 270316 13882 270332
rect 12797 270270 12813 270304
rect 13789 270270 13805 270304
rect 12720 270242 12754 270258
rect 12720 270158 12754 270174
rect 13848 270242 13882 270258
rect 13848 270158 13882 270174
rect 12797 270112 12813 270146
rect 13789 270112 13805 270146
rect 12720 270084 12754 270100
rect 12720 270000 12754 270016
rect 13848 270084 13882 270100
rect 13848 270000 13882 270016
rect 12797 269954 12813 269988
rect 13789 269954 13805 269988
rect 12720 269926 12754 269942
rect 12720 269842 12754 269858
rect 13848 269926 13882 269942
rect 13848 269842 13882 269858
rect 12797 269796 12813 269830
rect 13789 269796 13805 269830
rect 12720 269768 12754 269784
rect 12720 269684 12754 269700
rect 13848 269768 13882 269784
rect 13848 269684 13882 269700
rect 12797 269638 12813 269672
rect 13789 269638 13805 269672
rect 12720 269610 12754 269626
rect 12720 269526 12754 269542
rect 13848 269610 13882 269626
rect 13848 269526 13882 269542
rect 12797 269480 12813 269514
rect 13789 269480 13805 269514
rect 12618 269400 12652 269462
rect 14288 274412 14384 274446
rect 15558 274412 15654 274446
rect 14288 274350 14322 274412
rect 15620 274350 15654 274412
rect 14467 274298 14483 274332
rect 15459 274298 15475 274332
rect 14390 274270 14424 274286
rect 14390 274186 14424 274202
rect 15518 274270 15552 274286
rect 15518 274186 15552 274202
rect 14467 274140 14483 274174
rect 15459 274140 15475 274174
rect 14390 274112 14424 274128
rect 14390 274028 14424 274044
rect 15518 274112 15552 274128
rect 15518 274028 15552 274044
rect 14467 273982 14483 274016
rect 15459 273982 15475 274016
rect 14390 273954 14424 273970
rect 14390 273870 14424 273886
rect 15518 273954 15552 273970
rect 15518 273870 15552 273886
rect 14467 273824 14483 273858
rect 15459 273824 15475 273858
rect 14390 273796 14424 273812
rect 14390 273712 14424 273728
rect 15518 273796 15552 273812
rect 15518 273712 15552 273728
rect 14467 273666 14483 273700
rect 15459 273666 15475 273700
rect 15828 274412 15924 274446
rect 17098 274412 17194 274446
rect 15828 274350 15862 274412
rect 17160 274350 17194 274412
rect 16007 274298 16023 274332
rect 16999 274298 17015 274332
rect 15930 274270 15964 274286
rect 15930 274186 15964 274202
rect 17058 274270 17092 274286
rect 17058 274186 17092 274202
rect 16007 274140 16023 274174
rect 16999 274140 17015 274174
rect 15930 274112 15964 274128
rect 15930 274028 15964 274044
rect 17058 274112 17092 274128
rect 17058 274028 17092 274044
rect 16007 273982 16023 274016
rect 16999 273982 17015 274016
rect 15930 273954 15964 273970
rect 15930 273870 15964 273886
rect 17058 273954 17092 273970
rect 17058 273870 17092 273886
rect 16007 273824 16023 273858
rect 16999 273824 17015 273858
rect 15930 273796 15964 273812
rect 15930 273712 15964 273728
rect 17058 273796 17092 273812
rect 17058 273712 17092 273728
rect 14390 273638 14424 273654
rect 14390 273554 14424 273570
rect 15518 273638 15552 273654
rect 15518 273554 15552 273570
rect 14467 273508 14483 273542
rect 15459 273508 15475 273542
rect 14390 273480 14424 273496
rect 14390 273396 14424 273412
rect 15518 273480 15552 273496
rect 15518 273396 15552 273412
rect 14467 273350 14483 273384
rect 15459 273350 15475 273384
rect 14390 273322 14424 273338
rect 14390 273238 14424 273254
rect 15518 273322 15552 273338
rect 15518 273238 15552 273254
rect 14467 273192 14483 273226
rect 15459 273192 15475 273226
rect 14390 273164 14424 273180
rect 14390 273080 14424 273096
rect 15518 273164 15552 273180
rect 15518 273080 15552 273096
rect 16007 273666 16023 273700
rect 16999 273666 17015 273700
rect 15930 273638 15964 273654
rect 15930 273554 15964 273570
rect 17058 273638 17092 273654
rect 17058 273554 17092 273570
rect 16007 273508 16023 273542
rect 16999 273508 17015 273542
rect 15930 273480 15964 273496
rect 15930 273396 15964 273412
rect 17058 273480 17092 273496
rect 17058 273396 17092 273412
rect 16007 273350 16023 273384
rect 16999 273350 17015 273384
rect 15930 273322 15964 273338
rect 15930 273238 15964 273254
rect 17058 273322 17092 273338
rect 17058 273238 17092 273254
rect 16007 273192 16023 273226
rect 16999 273192 17015 273226
rect 14467 273034 14483 273068
rect 15459 273034 15475 273068
rect 14390 273006 14424 273022
rect 14390 272922 14424 272938
rect 15518 273006 15552 273022
rect 15518 272922 15552 272938
rect 14467 272876 14483 272910
rect 15459 272876 15475 272910
rect 14390 272848 14424 272864
rect 14390 272764 14424 272780
rect 15518 272848 15552 272864
rect 15518 272764 15552 272780
rect 14467 272718 14483 272752
rect 15459 272718 15475 272752
rect 14390 272690 14424 272706
rect 14390 272606 14424 272622
rect 15518 272690 15552 272706
rect 15518 272606 15552 272622
rect 14467 272560 14483 272594
rect 15459 272560 15475 272594
rect 14390 272532 14424 272548
rect 14390 272448 14424 272464
rect 15518 272532 15552 272548
rect 15518 272448 15552 272464
rect 14467 272402 14483 272436
rect 15459 272402 15475 272436
rect 14390 272374 14424 272390
rect 14390 272290 14424 272306
rect 15518 272374 15552 272390
rect 15518 272290 15552 272306
rect 14467 272244 14483 272278
rect 15459 272244 15475 272278
rect 14390 272216 14424 272232
rect 14390 272132 14424 272148
rect 15518 272216 15552 272232
rect 15518 272132 15552 272148
rect 15930 273164 15964 273180
rect 15930 273080 15964 273096
rect 17058 273164 17092 273180
rect 17058 273080 17092 273096
rect 16007 273034 16023 273068
rect 16999 273034 17015 273068
rect 15930 273006 15964 273022
rect 15930 272922 15964 272938
rect 17058 273006 17092 273022
rect 17058 272922 17092 272938
rect 16007 272876 16023 272910
rect 16999 272876 17015 272910
rect 15930 272848 15964 272864
rect 15930 272764 15964 272780
rect 17058 272848 17092 272864
rect 17058 272764 17092 272780
rect 16007 272718 16023 272752
rect 16999 272718 17015 272752
rect 15930 272690 15964 272706
rect 15930 272606 15964 272622
rect 17058 272690 17092 272706
rect 17058 272606 17092 272622
rect 16007 272560 16023 272594
rect 16999 272560 17015 272594
rect 15930 272532 15964 272548
rect 15930 272448 15964 272464
rect 17058 272532 17092 272548
rect 17058 272448 17092 272464
rect 16007 272402 16023 272436
rect 16999 272402 17015 272436
rect 15930 272374 15964 272390
rect 15930 272290 15964 272306
rect 17058 272374 17092 272390
rect 17058 272290 17092 272306
rect 16007 272244 16023 272278
rect 16999 272244 17015 272278
rect 14467 272086 14483 272120
rect 15459 272086 15475 272120
rect 14390 272058 14424 272074
rect 14390 271974 14424 271990
rect 15518 272058 15552 272074
rect 15518 271974 15552 271990
rect 14467 271928 14483 271962
rect 15459 271928 15475 271962
rect 14390 271900 14424 271916
rect 14390 271816 14424 271832
rect 15518 271900 15552 271916
rect 15518 271816 15552 271832
rect 14467 271770 14483 271804
rect 15459 271770 15475 271804
rect 14390 271742 14424 271758
rect 14390 271658 14424 271674
rect 15518 271742 15552 271758
rect 15518 271658 15552 271674
rect 14467 271612 14483 271646
rect 15459 271612 15475 271646
rect 15930 272216 15964 272232
rect 15930 272132 15964 272148
rect 17058 272216 17092 272232
rect 17058 272132 17092 272148
rect 16007 272086 16023 272120
rect 16999 272086 17015 272120
rect 15930 272058 15964 272074
rect 15930 271974 15964 271990
rect 17058 272058 17092 272074
rect 17058 271974 17092 271990
rect 16007 271928 16023 271962
rect 16999 271928 17015 271962
rect 15930 271900 15964 271916
rect 15930 271816 15964 271832
rect 17058 271900 17092 271916
rect 17058 271816 17092 271832
rect 16007 271770 16023 271804
rect 16999 271770 17015 271804
rect 15930 271742 15964 271758
rect 15930 271658 15964 271674
rect 17058 271742 17092 271758
rect 17058 271658 17092 271674
rect 14390 271584 14424 271600
rect 14390 271500 14424 271516
rect 15518 271584 15552 271600
rect 15518 271500 15552 271516
rect 14467 271454 14483 271488
rect 15459 271454 15475 271488
rect 14390 271426 14424 271442
rect 14390 271342 14424 271358
rect 15518 271426 15552 271442
rect 15518 271342 15552 271358
rect 14467 271296 14483 271330
rect 15459 271296 15475 271330
rect 14390 271268 14424 271284
rect 14390 271184 14424 271200
rect 15518 271268 15552 271284
rect 15518 271184 15552 271200
rect 14467 271138 14483 271172
rect 15459 271138 15475 271172
rect 14390 271110 14424 271126
rect 14390 271026 14424 271042
rect 15518 271110 15552 271126
rect 15518 271026 15552 271042
rect 14467 270980 14483 271014
rect 15459 270980 15475 271014
rect 14288 270900 14322 270962
rect 15620 270900 15654 270962
rect 14288 270866 14384 270900
rect 15558 270866 15654 270900
rect 16007 271612 16023 271646
rect 16999 271612 17015 271646
rect 15930 271584 15964 271600
rect 15930 271500 15964 271516
rect 17058 271584 17092 271600
rect 17058 271500 17092 271516
rect 16007 271454 16023 271488
rect 16999 271454 17015 271488
rect 15930 271426 15964 271442
rect 15930 271342 15964 271358
rect 17058 271426 17092 271442
rect 17058 271342 17092 271358
rect 16007 271296 16023 271330
rect 16999 271296 17015 271330
rect 15930 271268 15964 271284
rect 15930 271184 15964 271200
rect 17058 271268 17092 271284
rect 17058 271184 17092 271200
rect 16007 271138 16023 271172
rect 16999 271138 17015 271172
rect 15930 271110 15964 271126
rect 15930 271026 15964 271042
rect 17058 271110 17092 271126
rect 17058 271026 17092 271042
rect 16007 270980 16023 271014
rect 16999 270980 17015 271014
rect 15828 270900 15862 270962
rect 20446 274300 20542 274334
rect 21698 274300 21794 274334
rect 20446 274238 20480 274300
rect 21760 274238 21794 274300
rect 20616 274186 20632 274220
rect 21608 274186 21624 274220
rect 20548 274158 20582 274174
rect 20548 273974 20582 273990
rect 21658 274158 21692 274174
rect 21658 273974 21692 273990
rect 20616 273928 20632 273962
rect 21608 273928 21624 273962
rect 20548 273900 20582 273916
rect 20548 273716 20582 273732
rect 21658 273900 21692 273916
rect 21658 273716 21692 273732
rect 20616 273670 20632 273704
rect 21608 273670 21624 273704
rect 17405 273301 17501 273335
rect 18657 273301 18753 273335
rect 17405 273239 17439 273301
rect 18719 273239 18753 273301
rect 17575 273187 17591 273221
rect 18567 273187 18583 273221
rect 17507 273159 17541 273175
rect 17507 273075 17541 273091
rect 18617 273159 18651 273175
rect 18617 273075 18651 273091
rect 17575 273029 17591 273063
rect 18567 273029 18583 273063
rect 17507 273001 17541 273017
rect 17507 272917 17541 272933
rect 18617 273001 18651 273017
rect 18617 272917 18651 272933
rect 17575 272871 17591 272905
rect 18567 272871 18583 272905
rect 17507 272843 17541 272859
rect 17507 272759 17541 272775
rect 18617 272843 18651 272859
rect 18617 272759 18651 272775
rect 17575 272713 17591 272747
rect 18567 272713 18583 272747
rect 17507 272685 17541 272701
rect 17507 272601 17541 272617
rect 18617 272685 18651 272701
rect 18617 272601 18651 272617
rect 17575 272555 17591 272589
rect 18567 272555 18583 272589
rect 17507 272527 17541 272543
rect 17507 272443 17541 272459
rect 18617 272527 18651 272543
rect 18617 272443 18651 272459
rect 17575 272397 17591 272431
rect 18567 272397 18583 272431
rect 17507 272369 17541 272385
rect 17507 272285 17541 272301
rect 18617 272369 18651 272385
rect 18617 272285 18651 272301
rect 17575 272239 17591 272273
rect 18567 272239 18583 272273
rect 17507 272211 17541 272227
rect 17507 272127 17541 272143
rect 18617 272211 18651 272227
rect 18617 272127 18651 272143
rect 17575 272081 17591 272115
rect 18567 272081 18583 272115
rect 17405 272001 17439 272063
rect 18719 272001 18753 272063
rect 17405 271967 17501 272001
rect 18657 271967 18753 272001
rect 18925 273301 19021 273335
rect 20177 273301 20273 273335
rect 18925 273239 18959 273301
rect 20239 273239 20273 273301
rect 19095 273187 19111 273221
rect 20087 273187 20103 273221
rect 19027 273159 19061 273175
rect 19027 273075 19061 273091
rect 20137 273159 20171 273175
rect 20137 273075 20171 273091
rect 19095 273029 19111 273063
rect 20087 273029 20103 273063
rect 19027 273001 19061 273017
rect 19027 272917 19061 272933
rect 20137 273001 20171 273017
rect 20137 272917 20171 272933
rect 19095 272871 19111 272905
rect 20087 272871 20103 272905
rect 19027 272843 19061 272859
rect 19027 272759 19061 272775
rect 20137 272843 20171 272859
rect 20137 272759 20171 272775
rect 19095 272713 19111 272747
rect 20087 272713 20103 272747
rect 19027 272685 19061 272701
rect 19027 272601 19061 272617
rect 20137 272685 20171 272701
rect 20137 272601 20171 272617
rect 19095 272555 19111 272589
rect 20087 272555 20103 272589
rect 19027 272527 19061 272543
rect 19027 272443 19061 272459
rect 20137 272527 20171 272543
rect 20137 272443 20171 272459
rect 19095 272397 19111 272431
rect 20087 272397 20103 272431
rect 19027 272369 19061 272385
rect 19027 272285 19061 272301
rect 20137 272369 20171 272385
rect 20137 272285 20171 272301
rect 19095 272239 19111 272273
rect 20087 272239 20103 272273
rect 19027 272211 19061 272227
rect 19027 272127 19061 272143
rect 20137 272211 20171 272227
rect 20137 272127 20171 272143
rect 19095 272081 19111 272115
rect 20087 272081 20103 272115
rect 18925 272001 18959 272063
rect 20239 272001 20273 272063
rect 18925 271967 19021 272001
rect 20177 271967 20273 272001
rect 20548 273642 20582 273658
rect 20548 273458 20582 273474
rect 21658 273642 21692 273658
rect 21658 273458 21692 273474
rect 20616 273412 20632 273446
rect 21608 273412 21624 273446
rect 20548 273384 20582 273400
rect 20548 273200 20582 273216
rect 21658 273384 21692 273400
rect 21658 273200 21692 273216
rect 20616 273154 20632 273188
rect 21608 273154 21624 273188
rect 20548 273126 20582 273142
rect 20548 272942 20582 272958
rect 21658 273126 21692 273142
rect 21658 272942 21692 272958
rect 20616 272896 20632 272930
rect 21608 272896 21624 272930
rect 20548 272868 20582 272884
rect 20548 272684 20582 272700
rect 21658 272868 21692 272884
rect 21658 272684 21692 272700
rect 20616 272638 20632 272672
rect 21608 272638 21624 272672
rect 20548 272610 20582 272626
rect 20548 272426 20582 272442
rect 21658 272610 21692 272626
rect 21658 272426 21692 272442
rect 20616 272380 20632 272414
rect 21608 272380 21624 272414
rect 20548 272352 20582 272368
rect 20548 272168 20582 272184
rect 21658 272352 21692 272368
rect 21658 272168 21692 272184
rect 20616 272122 20632 272156
rect 21608 272122 21624 272156
rect 20548 272094 20582 272110
rect 20548 271910 20582 271926
rect 21658 272094 21692 272110
rect 21658 271910 21692 271926
rect 20616 271864 20632 271898
rect 21608 271864 21624 271898
rect 20548 271836 20582 271852
rect 20548 271652 20582 271668
rect 21658 271836 21692 271852
rect 21658 271652 21692 271668
rect 20616 271606 20632 271640
rect 21608 271606 21624 271640
rect 20548 271578 20582 271594
rect 20548 271394 20582 271410
rect 21658 271578 21692 271594
rect 21658 271394 21692 271410
rect 20616 271348 20632 271382
rect 21608 271348 21624 271382
rect 20548 271320 20582 271336
rect 20548 271136 20582 271152
rect 21658 271320 21692 271336
rect 21658 271136 21692 271152
rect 20616 271090 20632 271124
rect 21608 271090 21624 271124
rect 20446 271010 20480 271072
rect 21760 271010 21794 271072
rect 20446 270976 20542 271010
rect 21698 270976 21794 271010
rect 23280 274494 23314 274556
rect 22136 274442 22152 274476
rect 23128 274442 23144 274476
rect 22068 274414 22102 274430
rect 22068 274230 22102 274246
rect 23178 274414 23212 274430
rect 23178 274230 23212 274246
rect 22136 274184 22152 274218
rect 23128 274184 23144 274218
rect 22068 274156 22102 274172
rect 22068 273972 22102 273988
rect 23178 274156 23212 274172
rect 23178 273972 23212 273988
rect 22136 273926 22152 273960
rect 23128 273926 23144 273960
rect 22068 273898 22102 273914
rect 22068 273714 22102 273730
rect 23178 273898 23212 273914
rect 23178 273714 23212 273730
rect 22136 273668 22152 273702
rect 23128 273668 23144 273702
rect 22068 273640 22102 273656
rect 22068 273456 22102 273472
rect 23178 273640 23212 273656
rect 23178 273456 23212 273472
rect 22136 273410 22152 273444
rect 23128 273410 23144 273444
rect 22068 273382 22102 273398
rect 22068 273198 22102 273214
rect 23178 273382 23212 273398
rect 23178 273198 23212 273214
rect 22136 273152 22152 273186
rect 23128 273152 23144 273186
rect 22068 273124 22102 273140
rect 22068 272940 22102 272956
rect 23178 273124 23212 273140
rect 23178 272940 23212 272956
rect 22136 272894 22152 272928
rect 23128 272894 23144 272928
rect 22068 272866 22102 272882
rect 22068 272682 22102 272698
rect 23178 272866 23212 272882
rect 23178 272682 23212 272698
rect 22136 272636 22152 272670
rect 23128 272636 23144 272670
rect 22068 272608 22102 272624
rect 22068 272424 22102 272440
rect 23178 272608 23212 272624
rect 23178 272424 23212 272440
rect 22136 272378 22152 272412
rect 23128 272378 23144 272412
rect 22068 272350 22102 272366
rect 22068 272166 22102 272182
rect 23178 272350 23212 272366
rect 23178 272166 23212 272182
rect 22136 272120 22152 272154
rect 23128 272120 23144 272154
rect 22068 272092 22102 272108
rect 22068 271908 22102 271924
rect 23178 272092 23212 272108
rect 23178 271908 23212 271924
rect 22136 271862 22152 271896
rect 23128 271862 23144 271896
rect 17160 270900 17194 270962
rect 15828 270866 15924 270900
rect 17098 270866 17194 270900
rect 22068 271834 22102 271850
rect 22068 271650 22102 271666
rect 23178 271834 23212 271850
rect 23178 271650 23212 271666
rect 23998 273522 24094 273556
rect 25268 273522 25364 273556
rect 23998 273460 24032 273522
rect 25330 273460 25364 273522
rect 24177 273408 24193 273442
rect 25169 273408 25185 273442
rect 24100 273380 24134 273396
rect 24100 273196 24134 273212
rect 25228 273380 25262 273396
rect 25228 273196 25262 273212
rect 24177 273150 24193 273184
rect 25169 273150 25185 273184
rect 24100 273122 24134 273138
rect 24100 272938 24134 272954
rect 25228 273122 25262 273138
rect 25228 272938 25262 272954
rect 24177 272892 24193 272926
rect 25169 272892 25185 272926
rect 24100 272864 24134 272880
rect 24100 272680 24134 272696
rect 25228 272864 25262 272880
rect 25228 272680 25262 272696
rect 24177 272634 24193 272668
rect 25169 272634 25185 272668
rect 24100 272606 24134 272622
rect 24100 272422 24134 272438
rect 25228 272606 25262 272622
rect 25228 272422 25262 272438
rect 24177 272376 24193 272410
rect 25169 272376 25185 272410
rect 24100 272348 24134 272364
rect 24100 272164 24134 272180
rect 25228 272348 25262 272364
rect 25228 272164 25262 272180
rect 24177 272118 24193 272152
rect 25169 272118 25185 272152
rect 24100 272090 24134 272106
rect 24100 271906 24134 271922
rect 25228 272090 25262 272106
rect 25228 271906 25262 271922
rect 24177 271860 24193 271894
rect 25169 271860 25185 271894
rect 23998 271780 24032 271842
rect 25330 271780 25364 271842
rect 23998 271746 24094 271780
rect 25268 271746 25364 271780
rect 25498 273522 25594 273556
rect 26768 273522 26864 273556
rect 25498 273460 25532 273522
rect 26830 273460 26864 273522
rect 25677 273408 25693 273442
rect 26669 273408 26685 273442
rect 25600 273380 25634 273396
rect 25600 273196 25634 273212
rect 26728 273380 26762 273396
rect 26728 273196 26762 273212
rect 25677 273150 25693 273184
rect 26669 273150 26685 273184
rect 25600 273122 25634 273138
rect 25600 272938 25634 272954
rect 26728 273122 26762 273138
rect 26728 272938 26762 272954
rect 25677 272892 25693 272926
rect 26669 272892 26685 272926
rect 25600 272864 25634 272880
rect 25600 272680 25634 272696
rect 26728 272864 26762 272880
rect 26728 272680 26762 272696
rect 25677 272634 25693 272668
rect 26669 272634 26685 272668
rect 25600 272606 25634 272622
rect 25600 272422 25634 272438
rect 26728 272606 26762 272622
rect 26728 272422 26762 272438
rect 25677 272376 25693 272410
rect 26669 272376 26685 272410
rect 25600 272348 25634 272364
rect 25600 272164 25634 272180
rect 26728 272348 26762 272364
rect 26728 272164 26762 272180
rect 25677 272118 25693 272152
rect 26669 272118 26685 272152
rect 25600 272090 25634 272106
rect 25600 271906 25634 271922
rect 26728 272090 26762 272106
rect 26728 271906 26762 271922
rect 25677 271860 25693 271894
rect 26669 271860 26685 271894
rect 25498 271780 25532 271842
rect 28866 273507 28962 273541
rect 30118 273507 30214 273541
rect 28866 273445 28900 273507
rect 28116 273246 28212 273280
rect 28618 273246 28714 273280
rect 28116 273184 28150 273246
rect 27116 272890 27212 272924
rect 27868 272890 27964 272924
rect 27116 272828 27150 272890
rect 27930 272828 27964 272890
rect 27286 272776 27302 272810
rect 27778 272776 27794 272810
rect 27218 272748 27252 272764
rect 27218 272664 27252 272680
rect 27828 272748 27862 272764
rect 27828 272664 27862 272680
rect 27286 272618 27302 272652
rect 27778 272618 27794 272652
rect 27218 272590 27252 272606
rect 27218 272506 27252 272522
rect 27828 272590 27862 272606
rect 27828 272506 27862 272522
rect 27286 272460 27302 272494
rect 27778 272460 27794 272494
rect 27116 272380 27150 272442
rect 27930 272380 27964 272442
rect 27116 272346 27212 272380
rect 27868 272346 27964 272380
rect 28680 273184 28714 273246
rect 28286 273132 28302 273166
rect 28528 273132 28544 273166
rect 28218 273104 28252 273120
rect 28218 272920 28252 272936
rect 28578 273104 28612 273120
rect 28578 272920 28612 272936
rect 28286 272874 28302 272908
rect 28528 272874 28544 272908
rect 28218 272846 28252 272862
rect 28218 272662 28252 272678
rect 28578 272846 28612 272862
rect 28578 272662 28612 272678
rect 30180 273445 30214 273507
rect 29036 273393 29052 273427
rect 30028 273393 30044 273427
rect 28968 273365 29002 273381
rect 28968 273181 29002 273197
rect 30078 273365 30112 273381
rect 30078 273181 30112 273197
rect 29036 273135 29052 273169
rect 30028 273135 30044 273169
rect 28968 273107 29002 273123
rect 28968 272923 29002 272939
rect 30078 273107 30112 273123
rect 30078 272923 30112 272939
rect 29036 272877 29052 272911
rect 30028 272877 30044 272911
rect 28286 272616 28302 272650
rect 28528 272616 28544 272650
rect 28218 272588 28252 272604
rect 28218 272404 28252 272420
rect 28578 272588 28612 272604
rect 28578 272404 28612 272420
rect 28968 272849 29002 272865
rect 28968 272665 29002 272681
rect 30078 272849 30112 272865
rect 30078 272665 30112 272681
rect 30474 272829 30872 273941
rect 29036 272619 29052 272653
rect 30028 272619 30044 272653
rect 28286 272358 28302 272392
rect 28528 272358 28544 272392
rect 28218 272330 28252 272346
rect 28218 272146 28252 272162
rect 28578 272330 28612 272346
rect 28578 272146 28612 272162
rect 28286 272100 28302 272134
rect 28528 272100 28544 272134
rect 28116 272020 28150 272082
rect 28680 272020 28714 272082
rect 28116 271986 28212 272020
rect 28618 271986 28714 272020
rect 26830 271780 26864 271842
rect 25498 271746 25594 271780
rect 26768 271746 26864 271780
rect 28968 272591 29002 272607
rect 28968 272407 29002 272423
rect 30078 272591 30112 272607
rect 30078 272407 30112 272423
rect 29036 272361 29052 272395
rect 30028 272361 30044 272395
rect 28968 272333 29002 272349
rect 28968 272149 29002 272165
rect 30078 272333 30112 272349
rect 30078 272149 30112 272165
rect 29036 272103 29052 272137
rect 30028 272103 30044 272137
rect 28968 272075 29002 272091
rect 28968 271891 29002 271907
rect 30078 272075 30112 272091
rect 30078 271891 30112 271907
rect 29036 271845 29052 271879
rect 30028 271845 30044 271879
rect 28866 271765 28900 271827
rect 30180 271765 30214 271827
rect 28866 271731 28962 271765
rect 30118 271731 30214 271765
rect 22136 271604 22152 271638
rect 23128 271604 23144 271638
rect 22068 271576 22102 271592
rect 22068 271392 22102 271408
rect 23178 271576 23212 271592
rect 23178 271392 23212 271408
rect 22136 271346 22152 271380
rect 23128 271346 23144 271380
rect 22068 271318 22102 271334
rect 22068 271134 22102 271150
rect 23178 271318 23212 271334
rect 23178 271134 23212 271150
rect 22136 271088 22152 271122
rect 23128 271088 23144 271122
rect 22068 271060 22102 271076
rect 22068 270876 22102 270892
rect 23178 271060 23212 271076
rect 23178 270876 23212 270892
rect 22136 270830 22152 270864
rect 23128 270830 23144 270864
rect 21966 270750 22000 270812
rect 30474 271289 30872 272401
rect 537364 272058 537484 272074
rect 537364 271922 537484 271938
rect 543734 272058 543854 272074
rect 543734 271922 543854 271938
rect 23280 270750 23314 270812
rect 21966 270716 22062 270750
rect 23218 270716 23314 270750
rect 13950 269400 13984 269462
rect 12618 269366 12714 269400
rect 13888 269366 13984 269400
rect 31004 269200 31020 269440
rect 31260 269200 31276 269440
rect 32724 269200 32740 269440
rect 32980 269200 32996 269440
rect 34444 269200 34460 269440
rect 34700 269200 34716 269440
rect 35924 269200 35940 269440
rect 36180 269200 36196 269440
rect 37644 269200 37660 269440
rect 37900 269200 37916 269440
rect 39244 269200 39260 269440
rect 39500 269200 39516 269440
rect 40964 269200 40980 269440
rect 41220 269200 41236 269440
rect 42564 269200 42580 269440
rect 42820 269200 42836 269440
rect 44284 269200 44300 269440
rect 44540 269200 44556 269440
rect 537364 269058 537484 269074
rect 537364 268922 537484 268938
rect 543734 269058 543854 269074
rect 543734 268922 543854 268938
rect 11741 268653 11837 268687
rect 13051 268653 13147 268687
rect 11741 268591 11775 268653
rect 13113 268591 13147 268653
rect 13110 266670 13113 267330
rect 11741 265597 11775 265659
rect 13201 268653 13297 268687
rect 14511 268653 14607 268687
rect 13201 268591 13235 268653
rect 13147 266670 13201 267330
rect 13113 265597 13147 265659
rect 11741 265563 11837 265597
rect 13051 265563 13147 265597
rect 14573 268591 14607 268653
rect 13201 265597 13235 265659
rect 14573 265597 14607 265659
rect 13201 265563 13297 265597
rect 14511 265563 14607 265597
rect 5816 252444 5912 252478
rect 16068 252444 16164 252478
rect 5816 251270 5850 252444
rect 16130 252382 16164 252444
rect 5918 252315 5952 252331
rect 5986 252330 6002 252364
rect 15978 252330 15994 252364
rect 5918 252265 5952 252281
rect 5986 252232 6002 252266
rect 15978 252232 15994 252266
rect 16028 252217 16062 252233
rect 5918 252119 5952 252135
rect 5986 252134 6002 252168
rect 15978 252134 15994 252168
rect 16028 252167 16062 252183
rect 5918 252069 5952 252085
rect 5986 252036 6002 252070
rect 15978 252036 15994 252070
rect 16028 252021 16062 252037
rect 5918 251923 5952 251939
rect 5986 251938 6002 251972
rect 15978 251938 15994 251972
rect 16028 251971 16062 251987
rect 5918 251873 5952 251889
rect 5986 251840 6002 251874
rect 15978 251840 15994 251874
rect 16028 251825 16062 251841
rect 5918 251727 5952 251743
rect 5986 251742 6002 251776
rect 15978 251742 15994 251776
rect 16028 251775 16062 251791
rect 5918 251677 5952 251693
rect 5986 251644 6002 251678
rect 15978 251644 15994 251678
rect 16028 251629 16062 251645
rect 5918 251531 5952 251547
rect 5986 251546 6002 251580
rect 15978 251546 15994 251580
rect 16028 251579 16062 251595
rect 5918 251481 5952 251497
rect 5986 251448 6002 251482
rect 15978 251448 15994 251482
rect 16028 251433 16062 251449
rect 5986 251350 6002 251384
rect 15978 251350 15994 251384
rect 16028 251383 16062 251399
rect 16130 251270 16164 251332
rect 5816 251236 5912 251270
rect 16068 251236 16164 251270
rect 5816 242044 5912 242078
rect 16068 242044 16164 242078
rect 5816 240870 5850 242044
rect 16130 241982 16164 242044
rect 5918 241915 5952 241931
rect 5986 241930 6002 241964
rect 15978 241930 15994 241964
rect 5918 241865 5952 241881
rect 5986 241832 6002 241866
rect 15978 241832 15994 241866
rect 16028 241817 16062 241833
rect 5918 241719 5952 241735
rect 5986 241734 6002 241768
rect 15978 241734 15994 241768
rect 16028 241767 16062 241783
rect 5918 241669 5952 241685
rect 5986 241636 6002 241670
rect 15978 241636 15994 241670
rect 16028 241621 16062 241637
rect 5918 241523 5952 241539
rect 5986 241538 6002 241572
rect 15978 241538 15994 241572
rect 16028 241571 16062 241587
rect 5918 241473 5952 241489
rect 5986 241440 6002 241474
rect 15978 241440 15994 241474
rect 16028 241425 16062 241441
rect 5918 241327 5952 241343
rect 5986 241342 6002 241376
rect 15978 241342 15994 241376
rect 16028 241375 16062 241391
rect 5918 241277 5952 241293
rect 5986 241244 6002 241278
rect 15978 241244 15994 241278
rect 16028 241229 16062 241245
rect 5918 241131 5952 241147
rect 5986 241146 6002 241180
rect 15978 241146 15994 241180
rect 16028 241179 16062 241195
rect 5918 241081 5952 241097
rect 5986 241048 6002 241082
rect 15978 241048 15994 241082
rect 16028 241033 16062 241049
rect 5986 240950 6002 240984
rect 15978 240950 15994 240984
rect 16028 240983 16062 240999
rect 16130 240870 16164 240932
rect 5816 240836 5912 240870
rect 16068 240836 16164 240870
<< viali >>
rect 8420 304444 13560 304478
rect 6002 304330 15978 304364
rect 5918 304281 5952 304315
rect 6002 304232 15978 304266
rect 16028 304183 16062 304217
rect 6002 304134 15978 304168
rect 5918 304085 5952 304119
rect 6002 304036 15978 304070
rect 16028 303987 16062 304021
rect 6002 303938 15978 303972
rect 5918 303889 5952 303923
rect 6002 303840 15978 303874
rect 16028 303791 16062 303825
rect 6002 303742 15978 303776
rect 5918 303693 5952 303727
rect 6002 303644 15978 303678
rect 16028 303595 16062 303629
rect 6002 303546 15978 303580
rect 16130 303564 16164 304150
rect 5918 303497 5952 303531
rect 6002 303448 15978 303482
rect 16028 303399 16062 303433
rect 6002 303350 15978 303384
rect 8420 303236 13560 303270
rect 560097 305848 560131 305882
rect 560293 305848 560327 305882
rect 560489 305848 560523 305882
rect 560685 305848 560719 305882
rect 560881 305848 560915 305882
rect 559836 298240 559870 303380
rect 559950 295822 559984 305798
rect 560048 295822 560082 305798
rect 560146 295822 560180 305798
rect 560244 295822 560278 305798
rect 560342 295822 560376 305798
rect 560440 295822 560474 305798
rect 560538 295822 560572 305798
rect 560636 295822 560670 305798
rect 560734 295822 560768 305798
rect 560832 295822 560866 305798
rect 560930 295822 560964 305798
rect 561044 298240 561078 303380
rect 559999 295738 560033 295772
rect 560195 295738 560229 295772
rect 560391 295738 560425 295772
rect 560587 295738 560621 295772
rect 560783 295738 560817 295772
rect 560164 295636 560750 295670
rect 569297 305848 569331 305882
rect 569493 305848 569527 305882
rect 569689 305848 569723 305882
rect 569885 305848 569919 305882
rect 570081 305848 570115 305882
rect 569036 298240 569070 303380
rect 569150 295822 569184 305798
rect 569248 295822 569282 305798
rect 569346 295822 569380 305798
rect 569444 295822 569478 305798
rect 569542 295822 569576 305798
rect 569640 295822 569674 305798
rect 569738 295822 569772 305798
rect 569836 295822 569870 305798
rect 569934 295822 569968 305798
rect 570032 295822 570066 305798
rect 570130 295822 570164 305798
rect 570244 298240 570278 303380
rect 569199 295738 569233 295772
rect 569395 295738 569429 295772
rect 569591 295738 569625 295772
rect 569787 295738 569821 295772
rect 569983 295738 570017 295772
rect 569364 295636 569950 295670
rect 537969 294898 538059 294962
rect 538139 294898 538229 294962
rect 540459 294898 540549 294962
rect 540629 294898 540719 294962
rect 542919 294898 542999 294972
rect 543089 294898 543169 294972
rect 537969 294892 538059 294898
rect 538139 294892 538229 294898
rect 540459 294892 540549 294898
rect 540629 294892 540719 294898
rect 542919 294892 542999 294898
rect 543089 294892 543169 294898
rect 536380 294750 537356 294784
rect 537616 294750 538592 294784
rect 538852 294750 539828 294784
rect 540088 294750 541064 294784
rect 541324 294750 542300 294784
rect 542560 294750 543536 294784
rect 543796 294750 544772 294784
rect 536287 294654 536321 294722
rect 537415 294654 537449 294722
rect 537523 294654 537557 294722
rect 538651 294654 538685 294722
rect 538759 294654 538793 294722
rect 539887 294654 539921 294722
rect 539995 294654 540029 294722
rect 541123 294654 541157 294722
rect 541231 294654 541265 294722
rect 542359 294654 542393 294722
rect 542467 294654 542501 294722
rect 543595 294654 543629 294722
rect 543703 294654 543737 294722
rect 544831 294654 544865 294722
rect 536380 294592 537356 294626
rect 537616 294592 538592 294626
rect 538852 294592 539828 294626
rect 540088 294592 541064 294626
rect 541324 294592 542300 294626
rect 542560 294592 543536 294626
rect 543796 294592 544772 294626
rect 8420 294044 13560 294078
rect 6002 293930 15978 293964
rect 5918 293881 5952 293915
rect 6002 293832 15978 293866
rect 16028 293783 16062 293817
rect 6002 293734 15978 293768
rect 536380 294210 537356 294244
rect 537616 294210 538592 294244
rect 538852 294210 539828 294244
rect 540088 294210 541064 294244
rect 541324 294210 542300 294244
rect 542560 294210 543536 294244
rect 543796 294210 544772 294244
rect 536287 294114 536321 294182
rect 537415 294114 537449 294182
rect 537523 294114 537557 294182
rect 538651 294114 538685 294182
rect 538759 294114 538793 294182
rect 539887 294114 539921 294182
rect 539995 294114 540029 294182
rect 541123 294114 541157 294182
rect 541231 294114 541265 294182
rect 542359 294114 542393 294182
rect 542467 294114 542501 294182
rect 543595 294114 543629 294182
rect 543703 294114 543737 294182
rect 544831 294114 544865 294182
rect 536380 294052 537356 294086
rect 537616 294052 538592 294086
rect 538852 294052 539828 294086
rect 540088 294052 541064 294086
rect 541324 294052 542300 294086
rect 542560 294052 543536 294086
rect 543796 294052 544772 294086
rect 537979 293842 538069 293912
rect 538119 293842 538209 293912
rect 540459 293842 540549 293912
rect 540619 293852 540709 293922
rect 542919 293852 542999 293922
rect 543089 293852 543169 293922
rect 5918 293685 5952 293719
rect 6002 293636 15978 293670
rect 16028 293587 16062 293621
rect 6002 293538 15978 293572
rect 5918 293489 5952 293523
rect 6002 293440 15978 293474
rect 16028 293391 16062 293425
rect 6002 293342 15978 293376
rect 5918 293293 5952 293327
rect 6002 293244 15978 293278
rect 16028 293195 16062 293229
rect 6002 293146 15978 293180
rect 16130 293164 16164 293750
rect 536380 293670 537356 293704
rect 537616 293670 538592 293704
rect 538852 293670 539828 293704
rect 540088 293670 541064 293704
rect 541324 293670 542300 293704
rect 542560 293670 543536 293704
rect 543796 293670 544772 293704
rect 536287 293574 536321 293642
rect 537415 293574 537449 293642
rect 537523 293574 537557 293642
rect 538651 293574 538685 293642
rect 538759 293574 538793 293642
rect 539887 293574 539921 293642
rect 539995 293574 540029 293642
rect 541123 293574 541157 293642
rect 541231 293574 541265 293642
rect 542359 293574 542393 293642
rect 542467 293574 542501 293642
rect 543595 293574 543629 293642
rect 543703 293574 543737 293642
rect 544831 293574 544865 293642
rect 536380 293512 537356 293546
rect 537616 293512 538592 293546
rect 538852 293512 539828 293546
rect 540088 293512 541064 293546
rect 541324 293512 542300 293546
rect 542560 293512 543536 293546
rect 543796 293512 544772 293546
rect 537979 293302 538059 293382
rect 538149 293302 538229 293382
rect 540459 293302 540539 293382
rect 540629 293302 540709 293382
rect 542919 293302 542999 293382
rect 543089 293302 543169 293382
rect 5918 293097 5952 293131
rect 6002 293048 15978 293082
rect 16028 292999 16062 293033
rect 6002 292950 15978 292984
rect 8420 292836 13560 292870
rect 536380 293130 537356 293164
rect 537616 293130 538592 293164
rect 538852 293130 539828 293164
rect 540088 293130 541064 293164
rect 541324 293130 542300 293164
rect 542560 293130 543536 293164
rect 543796 293130 544772 293164
rect 536287 293034 536321 293102
rect 537415 293034 537449 293102
rect 537523 293034 537557 293102
rect 538651 293034 538685 293102
rect 538759 293034 538793 293102
rect 539887 293034 539921 293102
rect 539995 293034 540029 293102
rect 541123 293034 541157 293102
rect 541231 293034 541265 293102
rect 542359 293034 542393 293102
rect 542467 293034 542501 293102
rect 543595 293034 543629 293102
rect 543703 293034 543737 293102
rect 544831 293034 544865 293102
rect 536380 292972 537356 293006
rect 537616 292972 538592 293006
rect 538852 292972 539828 293006
rect 540088 292972 541064 293006
rect 541324 292972 542300 293006
rect 542560 292972 543536 293006
rect 543796 292972 544772 293006
rect 536380 292550 537356 292584
rect 537616 292550 538592 292584
rect 538852 292550 539828 292584
rect 540088 292550 541064 292584
rect 541324 292550 542300 292584
rect 542560 292550 543536 292584
rect 543796 292550 544772 292584
rect 536287 292454 536321 292522
rect 537415 292454 537449 292522
rect 537523 292454 537557 292522
rect 538651 292454 538685 292522
rect 538759 292454 538793 292522
rect 539887 292454 539921 292522
rect 539995 292454 540029 292522
rect 541123 292454 541157 292522
rect 541231 292454 541265 292522
rect 542359 292454 542393 292522
rect 542467 292454 542501 292522
rect 543595 292454 543629 292522
rect 543703 292454 543737 292522
rect 544831 292454 544865 292522
rect 536380 292392 537356 292426
rect 537616 292392 538592 292426
rect 538852 292392 539828 292426
rect 540088 292392 541064 292426
rect 541324 292392 542300 292426
rect 542560 292392 543536 292426
rect 543796 292392 544772 292426
rect 537979 292142 538069 292222
rect 538139 292142 538229 292222
rect 540459 292142 540539 292212
rect 540629 292142 540709 292212
rect 542919 292142 542999 292212
rect 543089 292142 543169 292212
rect 530740 290841 531137 291955
rect 533171 290841 533568 291955
rect 536380 291970 537356 292004
rect 537616 291970 538592 292004
rect 538852 291970 539828 292004
rect 540088 291970 541064 292004
rect 541324 291970 542300 292004
rect 542560 291970 543536 292004
rect 543796 291970 544772 292004
rect 536287 291874 536321 291942
rect 537415 291874 537449 291942
rect 537523 291874 537557 291942
rect 538651 291874 538685 291942
rect 538759 291874 538793 291942
rect 539887 291874 539921 291942
rect 539995 291874 540029 291942
rect 541123 291874 541157 291942
rect 541231 291874 541265 291942
rect 542359 291874 542393 291942
rect 542467 291874 542501 291942
rect 543595 291874 543629 291942
rect 543703 291874 543737 291942
rect 544831 291874 544865 291942
rect 536380 291812 537356 291846
rect 537616 291812 538592 291846
rect 538852 291812 539828 291846
rect 540088 291812 541064 291846
rect 541324 291812 542300 291846
rect 542560 291812 543536 291846
rect 543796 291812 544772 291846
rect 534540 291430 535516 291464
rect 535776 291430 536752 291464
rect 537012 291430 537988 291464
rect 538248 291430 539224 291464
rect 539484 291430 540460 291464
rect 540720 291430 541696 291464
rect 541956 291430 542932 291464
rect 543192 291430 544168 291464
rect 544428 291430 545404 291464
rect 545664 291430 546640 291464
rect 534447 291334 534481 291402
rect 535575 291334 535609 291402
rect 535683 291334 535717 291402
rect 536811 291334 536845 291402
rect 536919 291334 536953 291402
rect 538047 291334 538081 291402
rect 538155 291334 538189 291402
rect 539283 291334 539317 291402
rect 539391 291334 539425 291402
rect 540519 291334 540553 291402
rect 540627 291334 540661 291402
rect 541755 291334 541789 291402
rect 541863 291334 541897 291402
rect 542991 291334 543025 291402
rect 543099 291334 543133 291402
rect 544227 291334 544261 291402
rect 544335 291334 544369 291402
rect 545463 291334 545497 291402
rect 545571 291334 545605 291402
rect 546699 291334 546733 291402
rect 534540 291272 535516 291306
rect 535776 291272 536752 291306
rect 537012 291272 537988 291306
rect 538248 291272 539224 291306
rect 539484 291272 540460 291306
rect 540720 291272 541696 291306
rect 541956 291272 542932 291306
rect 543192 291272 544168 291306
rect 544428 291272 545404 291306
rect 545664 291272 546640 291306
rect 536119 291062 536209 291142
rect 536299 291062 536389 291142
rect 538649 291062 538739 291142
rect 538809 291062 538899 291142
rect 541119 291062 541209 291142
rect 541279 291062 541369 291142
rect 543569 291062 543659 291142
rect 543729 291062 543819 291142
rect 546069 291062 546159 291142
rect 546229 291062 546319 291142
rect 534540 290890 535516 290924
rect 535776 290890 536752 290924
rect 537012 290890 537988 290924
rect 538248 290890 539224 290924
rect 539484 290890 540460 290924
rect 540720 290890 541696 290924
rect 541956 290890 542932 290924
rect 543192 290890 544168 290924
rect 544428 290890 545404 290924
rect 545664 290890 546640 290924
rect 534447 290794 534481 290862
rect 535575 290794 535609 290862
rect 535683 290794 535717 290862
rect 536811 290794 536845 290862
rect 536919 290794 536953 290862
rect 538047 290794 538081 290862
rect 538155 290794 538189 290862
rect 539283 290794 539317 290862
rect 539391 290794 539425 290862
rect 540519 290794 540553 290862
rect 540627 290794 540661 290862
rect 541755 290794 541789 290862
rect 541863 290794 541897 290862
rect 542991 290794 543025 290862
rect 543099 290794 543133 290862
rect 544227 290794 544261 290862
rect 544335 290794 544369 290862
rect 545463 290794 545497 290862
rect 545571 290794 545605 290862
rect 546699 290794 546733 290862
rect 534540 290732 535516 290766
rect 535776 290732 536752 290766
rect 537012 290732 537988 290766
rect 538248 290732 539224 290766
rect 539484 290732 540460 290766
rect 540720 290732 541696 290766
rect 541956 290732 542932 290766
rect 543192 290732 544168 290766
rect 544428 290732 545404 290766
rect 545664 290732 546640 290766
rect 547800 290841 548197 291955
rect 550231 290841 550628 291955
rect 530740 289371 531137 290485
rect 533171 289371 533568 290485
rect 534540 290350 535516 290384
rect 535776 290350 536752 290384
rect 537012 290350 537988 290384
rect 538248 290350 539224 290384
rect 539484 290350 540460 290384
rect 540720 290350 541696 290384
rect 541956 290350 542932 290384
rect 543192 290350 544168 290384
rect 544428 290350 545404 290384
rect 545664 290350 546640 290384
rect 534447 290254 534481 290322
rect 535575 290254 535609 290322
rect 535683 290254 535717 290322
rect 536811 290254 536845 290322
rect 536919 290254 536953 290322
rect 538047 290254 538081 290322
rect 538155 290254 538189 290322
rect 539283 290254 539317 290322
rect 539391 290254 539425 290322
rect 540519 290254 540553 290322
rect 540627 290254 540661 290322
rect 541755 290254 541789 290322
rect 541863 290254 541897 290322
rect 542991 290254 543025 290322
rect 543099 290254 543133 290322
rect 544227 290254 544261 290322
rect 544335 290254 544369 290322
rect 545463 290254 545497 290322
rect 545571 290254 545605 290322
rect 546699 290254 546733 290322
rect 534540 290192 535516 290226
rect 535776 290192 536752 290226
rect 537012 290192 537988 290226
rect 538248 290192 539224 290226
rect 539484 290192 540460 290226
rect 540720 290192 541696 290226
rect 541956 290192 542932 290226
rect 543192 290192 544168 290226
rect 544428 290192 545404 290226
rect 545664 290192 546640 290226
rect 536119 289982 536209 290062
rect 536299 289992 536389 290072
rect 538649 289982 538739 290062
rect 538809 289982 538899 290062
rect 541119 289982 541209 290062
rect 541279 289982 541369 290062
rect 543569 289982 543659 290062
rect 543729 289982 543819 290062
rect 546069 289982 546159 290062
rect 546229 289982 546319 290062
rect 534540 289810 535516 289844
rect 535776 289810 536752 289844
rect 537012 289810 537988 289844
rect 538248 289810 539224 289844
rect 539484 289810 540460 289844
rect 540720 289810 541696 289844
rect 541956 289810 542932 289844
rect 543192 289810 544168 289844
rect 544428 289810 545404 289844
rect 545664 289810 546640 289844
rect 534447 289714 534481 289782
rect 535575 289714 535609 289782
rect 535683 289714 535717 289782
rect 536811 289714 536845 289782
rect 536919 289714 536953 289782
rect 538047 289714 538081 289782
rect 538155 289714 538189 289782
rect 539283 289714 539317 289782
rect 539391 289714 539425 289782
rect 540519 289714 540553 289782
rect 540627 289714 540661 289782
rect 541755 289714 541789 289782
rect 541863 289714 541897 289782
rect 542991 289714 543025 289782
rect 543099 289714 543133 289782
rect 544227 289714 544261 289782
rect 544335 289714 544369 289782
rect 545463 289714 545497 289782
rect 545571 289714 545605 289782
rect 546699 289714 546733 289782
rect 534540 289652 535516 289686
rect 535776 289652 536752 289686
rect 537012 289652 537988 289686
rect 538248 289652 539224 289686
rect 539484 289652 540460 289686
rect 540720 289652 541696 289686
rect 541956 289652 542932 289686
rect 543192 289652 544168 289686
rect 544428 289652 545404 289686
rect 545664 289652 546640 289686
rect 531759 289225 531849 289252
rect 531969 289225 532059 289252
rect 547800 289371 548197 290485
rect 550231 289371 550628 290485
rect 549069 289225 549139 289242
rect 549229 289225 549299 289242
rect 531759 289122 531849 289225
rect 531969 289122 532059 289225
rect 549069 289152 549139 289225
rect 549229 289152 549299 289225
rect 536471 289030 537447 289064
rect 537689 289030 538665 289064
rect 538907 289030 539883 289064
rect 540125 289030 541101 289064
rect 541343 289030 542319 289064
rect 542561 289030 543537 289064
rect 543779 289030 544755 289064
rect 536387 288934 536421 289002
rect 537497 288934 537531 289002
rect 537605 288934 537639 289002
rect 538715 288934 538749 289002
rect 538823 288934 538857 289002
rect 539933 288934 539967 289002
rect 540041 288934 540075 289002
rect 541151 288934 541185 289002
rect 541259 288934 541293 289002
rect 542369 288934 542403 289002
rect 542477 288934 542511 289002
rect 543587 288934 543621 289002
rect 543695 288934 543729 289002
rect 544805 288934 544839 289002
rect 536471 288872 537447 288906
rect 537689 288872 538665 288906
rect 538907 288872 539883 288906
rect 540125 288872 541101 288906
rect 541343 288872 542319 288906
rect 542561 288872 543537 288906
rect 543779 288872 544755 288906
rect 538279 288758 538389 288772
rect 539139 288758 539249 288772
rect 540349 288758 540459 288772
rect 541199 288758 541309 288772
rect 542769 288758 542879 288772
rect 543649 288758 543759 288772
rect 570720 288824 575860 288858
rect 538279 288678 538389 288758
rect 539139 288678 539249 288758
rect 540349 288678 540459 288758
rect 541199 288678 541309 288758
rect 542769 288678 542879 288758
rect 543649 288678 543759 288758
rect 538279 288662 538389 288678
rect 539139 288662 539249 288678
rect 540349 288662 540459 288678
rect 541199 288662 541309 288678
rect 542769 288662 542879 288678
rect 543649 288662 543759 288678
rect 536471 288530 537447 288564
rect 537689 288530 538665 288564
rect 538907 288530 539883 288564
rect 540125 288530 541101 288564
rect 541343 288530 542319 288564
rect 542561 288530 543537 288564
rect 543779 288530 544755 288564
rect 536387 288434 536421 288502
rect 537497 288434 537531 288502
rect 537605 288434 537639 288502
rect 538715 288434 538749 288502
rect 538823 288434 538857 288502
rect 539933 288434 539967 288502
rect 540041 288434 540075 288502
rect 541151 288434 541185 288502
rect 541259 288434 541293 288502
rect 542369 288434 542403 288502
rect 542477 288434 542511 288502
rect 543587 288434 543621 288502
rect 543695 288434 543729 288502
rect 544805 288434 544839 288502
rect 536471 288372 537447 288406
rect 537689 288372 538665 288406
rect 538907 288372 539883 288406
rect 540125 288372 541101 288406
rect 541343 288372 542319 288406
rect 542561 288372 543537 288406
rect 543779 288372 544755 288406
rect 568302 288710 578278 288744
rect 568218 288661 568252 288695
rect 568302 288612 578278 288646
rect 578328 288563 578362 288597
rect 537031 288030 538007 288064
rect 538249 288030 539225 288064
rect 539467 288030 540443 288064
rect 540685 288030 541661 288064
rect 541903 288030 542879 288064
rect 543121 288030 544097 288064
rect 536947 287834 536981 288002
rect 538057 287834 538091 288002
rect 538165 287834 538199 288002
rect 539275 287834 539309 288002
rect 539383 287834 539417 288002
rect 540493 287834 540527 288002
rect 540601 287834 540635 288002
rect 541711 287834 541745 288002
rect 541819 287834 541853 288002
rect 542929 287834 542963 288002
rect 543037 287834 543071 288002
rect 544147 287834 544181 288002
rect 537031 287772 538007 287806
rect 538249 287772 539225 287806
rect 539467 287772 540443 287806
rect 540685 287772 541661 287806
rect 541903 287772 542879 287806
rect 543121 287772 544097 287806
rect 568116 287944 568150 288530
rect 568302 288514 578278 288548
rect 568218 288465 568252 288499
rect 568302 288416 578278 288450
rect 578328 288367 578362 288401
rect 568302 288318 578278 288352
rect 568218 288269 568252 288303
rect 568302 288220 578278 288254
rect 578328 288171 578362 288205
rect 568302 288122 578278 288156
rect 568218 288073 568252 288107
rect 568302 288024 578278 288058
rect 578328 287975 578362 288009
rect 568302 287926 578278 287960
rect 568218 287877 568252 287911
rect 568302 287828 578278 287862
rect 578328 287779 578362 287813
rect 568302 287730 578278 287764
rect 537569 287562 537679 287652
rect 542479 287562 542589 287652
rect 570720 287616 575860 287650
rect 537031 287410 538007 287444
rect 538249 287410 539225 287444
rect 539467 287410 540443 287444
rect 540685 287410 541661 287444
rect 541903 287410 542879 287444
rect 543121 287410 544097 287444
rect 536947 287214 536981 287382
rect 538057 287214 538091 287382
rect 538165 287214 538199 287382
rect 539275 287214 539309 287382
rect 539383 287214 539417 287382
rect 540493 287214 540527 287382
rect 540601 287214 540635 287382
rect 541711 287214 541745 287382
rect 541819 287214 541853 287382
rect 542929 287214 542963 287382
rect 543037 287214 543071 287382
rect 544147 287214 544181 287382
rect 537031 287152 538007 287186
rect 538249 287152 539225 287186
rect 539467 287152 540443 287186
rect 540685 287152 541661 287186
rect 541903 287152 542879 287186
rect 543121 287152 544097 287186
rect 536471 286810 537447 286844
rect 537689 286810 538665 286844
rect 538907 286810 539883 286844
rect 540125 286810 541101 286844
rect 541343 286810 542319 286844
rect 542561 286810 543537 286844
rect 543779 286810 544755 286844
rect 536387 286614 536421 286782
rect 537497 286614 537531 286782
rect 537605 286614 537639 286782
rect 538715 286614 538749 286782
rect 538823 286614 538857 286782
rect 539933 286614 539967 286782
rect 540041 286614 540075 286782
rect 541151 286614 541185 286782
rect 541259 286614 541293 286782
rect 542369 286614 542403 286782
rect 542477 286614 542511 286782
rect 543587 286614 543621 286782
rect 543695 286614 543729 286782
rect 544805 286614 544839 286782
rect 536471 286552 537447 286586
rect 537689 286552 538665 286586
rect 538907 286552 539883 286586
rect 540125 286552 541101 286586
rect 541343 286552 542319 286586
rect 542561 286552 543537 286586
rect 543779 286552 544755 286586
rect 537509 286438 537629 286452
rect 538729 286438 538849 286452
rect 539939 286438 540059 286452
rect 541159 286438 541279 286452
rect 542389 286438 542509 286442
rect 543599 286438 543719 286452
rect 537509 286358 537629 286438
rect 538729 286358 538849 286438
rect 539939 286358 540059 286438
rect 541159 286358 541279 286438
rect 542389 286358 542509 286438
rect 543599 286358 543719 286438
rect 537509 286352 537629 286358
rect 538729 286352 538849 286358
rect 539939 286352 540059 286358
rect 541159 286352 541279 286358
rect 542389 286342 542509 286358
rect 543599 286352 543719 286358
rect 536471 286210 537447 286244
rect 537689 286210 538665 286244
rect 538907 286210 539883 286244
rect 540125 286210 541101 286244
rect 541343 286210 542319 286244
rect 542561 286210 543537 286244
rect 543779 286210 544755 286244
rect 536387 286014 536421 286182
rect 537497 286014 537531 286182
rect 537605 286014 537639 286182
rect 538715 286014 538749 286182
rect 538823 286014 538857 286182
rect 539933 286014 539967 286182
rect 540041 286014 540075 286182
rect 541151 286014 541185 286182
rect 541259 286014 541293 286182
rect 542369 286014 542403 286182
rect 542477 286014 542511 286182
rect 543587 286014 543621 286182
rect 543695 286014 543729 286182
rect 544805 286014 544839 286182
rect 536471 285952 537447 285986
rect 537689 285952 538665 285986
rect 538907 285952 539883 285986
rect 540125 285952 541101 285986
rect 541343 285952 542319 285986
rect 542561 285952 543537 285986
rect 543779 285952 544755 285986
rect 537384 285384 537544 285478
rect 538444 285384 538604 285478
rect 539904 285384 540064 285478
rect 541124 285384 541284 285478
rect 542604 285384 542764 285478
rect 543604 285384 543764 285478
rect 537384 285350 537544 285384
rect 538444 285350 538604 285384
rect 539904 285350 540064 285384
rect 541124 285350 541284 285384
rect 542604 285350 542764 285384
rect 543604 285350 543764 285384
rect 537384 285318 537544 285350
rect 538444 285318 538604 285350
rect 539904 285318 540064 285350
rect 541124 285318 541284 285350
rect 542604 285318 542764 285350
rect 543604 285318 543764 285350
rect 537025 285236 538001 285270
rect 538261 285236 539237 285270
rect 539497 285236 540473 285270
rect 540733 285236 541709 285270
rect 541969 285236 542945 285270
rect 543205 285236 544181 285270
rect 536932 285040 536966 285208
rect 538060 285040 538094 285208
rect 538168 285040 538202 285208
rect 539296 285040 539330 285208
rect 539404 285040 539438 285208
rect 540532 285040 540566 285208
rect 540640 285040 540674 285208
rect 541768 285040 541802 285208
rect 541876 285040 541910 285208
rect 543004 285040 543038 285208
rect 543112 285040 543146 285208
rect 544240 285040 544274 285208
rect 537025 284978 538001 285012
rect 538261 284978 539237 285012
rect 539497 284978 540473 285012
rect 540733 284978 541709 285012
rect 541969 284978 542945 285012
rect 543205 284978 544181 285012
rect 537384 284864 537544 284898
rect 538444 284864 538604 284898
rect 539904 284864 540064 284898
rect 541124 284864 541284 284898
rect 542604 284864 542764 284898
rect 543604 284864 543764 284898
rect 537384 284794 537544 284864
rect 538444 284794 538604 284864
rect 539904 284794 540064 284864
rect 541124 284794 541284 284864
rect 542604 284794 542764 284864
rect 543604 284794 543764 284864
rect 537384 284760 537544 284794
rect 538444 284760 538604 284794
rect 539904 284760 540064 284794
rect 541124 284760 541284 284794
rect 542604 284760 542764 284794
rect 543604 284760 543764 284794
rect 537384 284738 537544 284760
rect 538444 284738 538604 284760
rect 539904 284738 540064 284760
rect 541124 284738 541284 284760
rect 542604 284738 542764 284760
rect 543604 284738 543764 284760
rect 537025 284646 538001 284680
rect 538261 284646 539237 284680
rect 539497 284646 540473 284680
rect 540733 284646 541709 284680
rect 541969 284646 542945 284680
rect 543205 284646 544181 284680
rect 536932 284450 536966 284618
rect 538060 284450 538094 284618
rect 538168 284450 538202 284618
rect 539296 284450 539330 284618
rect 539404 284450 539438 284618
rect 540532 284450 540566 284618
rect 540640 284450 540674 284618
rect 541768 284450 541802 284618
rect 541876 284450 541910 284618
rect 543004 284450 543038 284618
rect 543112 284450 543146 284618
rect 544240 284450 544274 284618
rect 537025 284388 538001 284422
rect 538261 284388 539237 284422
rect 539497 284388 540473 284422
rect 540733 284388 541709 284422
rect 541969 284388 542945 284422
rect 543205 284388 544181 284422
rect 539786 283856 540012 283890
rect 540254 283856 540480 283890
rect 540722 283856 540948 283890
rect 541190 283856 541416 283890
rect 539702 283660 539736 283828
rect 540062 283660 540096 283828
rect 540170 283660 540204 283828
rect 540530 283660 540564 283828
rect 540638 283660 540672 283828
rect 540998 283660 541032 283828
rect 541106 283660 541140 283828
rect 541466 283660 541500 283828
rect 539786 283598 540012 283632
rect 540254 283598 540480 283632
rect 540722 283598 540948 283632
rect 541190 283598 541416 283632
rect 539764 283484 539984 283518
rect 540284 283484 540504 283518
rect 540704 283484 540924 283518
rect 541254 283484 541474 283518
rect 539764 283379 539984 283484
rect 540284 283379 540504 283484
rect 540704 283379 540924 283484
rect 541254 283379 541474 283484
rect 539764 283368 539916 283379
rect 539916 283368 539984 283379
rect 540284 283368 540504 283379
rect 540704 283368 540924 283379
rect 541254 283368 541290 283379
rect 541290 283368 541474 283379
rect 540006 283231 540482 283265
rect 540724 283231 541200 283265
rect 539922 283135 539956 283203
rect 540532 283135 540566 283203
rect 540640 283135 540674 283203
rect 541250 283135 541284 283203
rect 540006 283073 540482 283107
rect 540724 283073 541200 283107
rect 537404 282854 537584 282958
rect 538544 282854 538724 282958
rect 539524 282854 539704 282968
rect 540294 282959 540474 282968
rect 540734 282959 540914 282968
rect 540294 282854 540474 282959
rect 540734 282854 540914 282959
rect 541454 282854 541634 282958
rect 542524 282854 542704 282968
rect 543524 282854 543704 282968
rect 537404 282828 537584 282854
rect 538544 282828 538724 282854
rect 539524 282838 539704 282854
rect 540294 282838 540474 282854
rect 540734 282838 540914 282854
rect 541454 282828 541634 282854
rect 542524 282838 542704 282854
rect 543524 282838 543704 282854
rect 537071 282706 538047 282740
rect 538289 282706 539265 282740
rect 539507 282706 540483 282740
rect 540725 282706 541701 282740
rect 541943 282706 542919 282740
rect 543161 282706 544137 282740
rect 536987 282510 537021 282678
rect 538097 282510 538131 282678
rect 538205 282510 538239 282678
rect 539315 282510 539349 282678
rect 539423 282510 539457 282678
rect 540533 282510 540567 282678
rect 540641 282510 540675 282678
rect 541751 282510 541785 282678
rect 541859 282510 541893 282678
rect 542969 282510 543003 282678
rect 543077 282510 543111 282678
rect 544187 282510 544221 282678
rect 537071 282448 538047 282482
rect 538289 282448 539265 282482
rect 539507 282448 540483 282482
rect 540725 282448 541701 282482
rect 541943 282448 542919 282482
rect 543161 282448 544137 282482
rect 537777 281587 538891 281984
rect 539297 281587 540411 281984
rect 540807 281593 541921 281990
rect 542317 281593 543431 281990
rect 570740 281344 575880 281378
rect 537364 280938 537484 281058
rect 543734 280938 543854 281058
rect 568322 281230 578298 281264
rect 568238 281181 568272 281215
rect 568322 281132 578298 281166
rect 578348 281083 578382 281117
rect 568136 280464 568170 281050
rect 568322 281034 578298 281068
rect 568238 280985 568272 281019
rect 568322 280936 578298 280970
rect 578348 280887 578382 280921
rect 568322 280838 578298 280872
rect 568238 280789 568272 280823
rect 568322 280740 578298 280774
rect 578348 280691 578382 280725
rect 568322 280642 578298 280676
rect 568238 280593 568272 280627
rect 568322 280544 578298 280578
rect 578348 280495 578382 280529
rect 568322 280446 578298 280480
rect 568238 280397 568272 280431
rect 568322 280348 578298 280382
rect 578348 280299 578382 280333
rect 568322 280250 578298 280284
rect 570740 280136 575880 280170
rect 11887 279212 13001 279609
rect 11887 276781 13001 277178
rect 13347 279212 14461 279609
rect 14540 278370 14573 278550
rect 14573 278370 14607 278550
rect 14607 278370 14640 278550
rect 14540 277950 14573 278130
rect 14573 277950 14607 278130
rect 14607 277950 14640 278130
rect 13347 276781 14461 277178
rect 537364 277938 537484 278058
rect 543734 277938 543854 278058
rect 31020 275900 31260 276140
rect 32740 275900 32980 276140
rect 34460 275900 34700 276140
rect 35940 275900 36180 276140
rect 37660 275900 37900 276140
rect 39260 275900 39500 276140
rect 40980 275900 41220 276140
rect 42580 275900 42820 276140
rect 44300 275900 44540 276140
rect 12813 275800 13789 275834
rect 12720 275704 12754 275772
rect 13848 275704 13882 275772
rect 12813 275642 13789 275676
rect 12720 275546 12754 275614
rect 13848 275546 13882 275614
rect 12813 275484 13789 275518
rect 12720 275388 12754 275456
rect 13848 275388 13882 275456
rect 12813 275326 13789 275360
rect 12720 275230 12754 275298
rect 13848 275230 13882 275298
rect 12813 275168 13789 275202
rect 12720 275072 12754 275140
rect 13848 275072 13882 275140
rect 12813 275010 13789 275044
rect 12720 274914 12754 274982
rect 13848 274914 13882 274982
rect 12813 274852 13789 274886
rect 12720 274756 12754 274824
rect 13848 274756 13882 274824
rect 12813 274694 13789 274728
rect 12720 274598 12754 274666
rect 13848 274598 13882 274666
rect 12813 274536 13789 274570
rect 12720 274440 12754 274508
rect 13848 274440 13882 274508
rect 12813 274378 13789 274412
rect 12618 271029 12652 274285
rect 12720 274282 12754 274350
rect 13848 274282 13882 274350
rect 537364 274938 537484 275058
rect 543734 274938 543854 275058
rect 12813 274220 13789 274254
rect 12720 274124 12754 274192
rect 13848 274124 13882 274192
rect 12813 274062 13789 274096
rect 12720 273966 12754 274034
rect 13848 273966 13882 274034
rect 12813 273904 13789 273938
rect 12720 273808 12754 273876
rect 13848 273808 13882 273876
rect 12813 273746 13789 273780
rect 12720 273650 12754 273718
rect 13848 273650 13882 273718
rect 12813 273588 13789 273622
rect 12720 273492 12754 273560
rect 13848 273492 13882 273560
rect 12813 273430 13789 273464
rect 12720 273334 12754 273402
rect 13848 273334 13882 273402
rect 12813 273272 13789 273306
rect 12720 273176 12754 273244
rect 13848 273176 13882 273244
rect 12813 273114 13789 273148
rect 12720 273018 12754 273086
rect 13848 273018 13882 273086
rect 12813 272956 13789 272990
rect 12720 272860 12754 272928
rect 13848 272860 13882 272928
rect 12813 272798 13789 272832
rect 12720 272702 12754 272770
rect 13848 272702 13882 272770
rect 12813 272640 13789 272674
rect 12720 272544 12754 272612
rect 13848 272544 13882 272612
rect 12813 272482 13789 272516
rect 12720 272386 12754 272454
rect 13848 272386 13882 272454
rect 12813 272324 13789 272358
rect 12720 272228 12754 272296
rect 13848 272228 13882 272296
rect 12813 272166 13789 272200
rect 12720 272070 12754 272138
rect 13848 272070 13882 272138
rect 12813 272008 13789 272042
rect 12720 271912 12754 271980
rect 13848 271912 13882 271980
rect 12813 271850 13789 271884
rect 12720 271754 12754 271822
rect 13848 271754 13882 271822
rect 12813 271692 13789 271726
rect 12720 271596 12754 271664
rect 13848 271596 13882 271664
rect 12813 271534 13789 271568
rect 12720 271438 12754 271506
rect 13848 271438 13882 271506
rect 12813 271376 13789 271410
rect 12720 271280 12754 271348
rect 13848 271280 13882 271348
rect 12813 271218 13789 271252
rect 12720 271122 12754 271190
rect 13848 271122 13882 271190
rect 12813 271060 13789 271094
rect 12720 270964 12754 271032
rect 13848 270964 13882 271032
rect 13950 271029 13984 274285
rect 12813 270902 13789 270936
rect 12720 270806 12754 270874
rect 13848 270806 13882 270874
rect 12813 270744 13789 270778
rect 12720 270648 12754 270716
rect 13848 270648 13882 270716
rect 12813 270586 13789 270620
rect 12720 270490 12754 270558
rect 13848 270490 13882 270558
rect 12813 270428 13789 270462
rect 12720 270332 12754 270400
rect 13848 270332 13882 270400
rect 12813 270270 13789 270304
rect 12720 270174 12754 270242
rect 13848 270174 13882 270242
rect 12813 270112 13789 270146
rect 12720 270016 12754 270084
rect 13848 270016 13882 270084
rect 12813 269954 13789 269988
rect 12720 269858 12754 269926
rect 13848 269858 13882 269926
rect 12813 269796 13789 269830
rect 12720 269700 12754 269768
rect 13848 269700 13882 269768
rect 12813 269638 13789 269672
rect 12720 269542 12754 269610
rect 13848 269542 13882 269610
rect 12813 269480 13789 269514
rect 14483 274298 15459 274332
rect 14390 274202 14424 274270
rect 15518 274202 15552 274270
rect 14483 274140 15459 274174
rect 14390 274044 14424 274112
rect 15518 274044 15552 274112
rect 14483 273982 15459 274016
rect 14390 273886 14424 273954
rect 15518 273886 15552 273954
rect 14483 273824 15459 273858
rect 14390 273728 14424 273796
rect 15518 273728 15552 273796
rect 14483 273666 15459 273700
rect 16023 274298 16999 274332
rect 15930 274202 15964 274270
rect 17058 274202 17092 274270
rect 16023 274140 16999 274174
rect 15930 274044 15964 274112
rect 17058 274044 17092 274112
rect 16023 273982 16999 274016
rect 15930 273886 15964 273954
rect 17058 273886 17092 273954
rect 16023 273824 16999 273858
rect 15930 273728 15964 273796
rect 17058 273728 17092 273796
rect 14390 273570 14424 273638
rect 15518 273570 15552 273638
rect 14288 271778 14322 273534
rect 14483 273508 15459 273542
rect 14390 273412 14424 273480
rect 15518 273412 15552 273480
rect 14483 273350 15459 273384
rect 14390 273254 14424 273322
rect 15518 273254 15552 273322
rect 14483 273192 15459 273226
rect 14390 273096 14424 273164
rect 15518 273096 15552 273164
rect 15620 273110 15654 273680
rect 15654 273110 15828 273680
rect 15828 273110 15860 273680
rect 16023 273666 16999 273700
rect 15930 273570 15964 273638
rect 17058 273570 17092 273638
rect 16023 273508 16999 273542
rect 15930 273412 15964 273480
rect 17058 273412 17092 273480
rect 16023 273350 16999 273384
rect 15930 273254 15964 273322
rect 17058 273254 17092 273322
rect 16023 273192 16999 273226
rect 14483 273034 15459 273068
rect 14390 272938 14424 273006
rect 15518 272938 15552 273006
rect 14483 272876 15459 272910
rect 14390 272780 14424 272848
rect 15518 272780 15552 272848
rect 14483 272718 15459 272752
rect 14390 272622 14424 272690
rect 15518 272622 15552 272690
rect 14483 272560 15459 272594
rect 14390 272464 14424 272532
rect 15518 272464 15552 272532
rect 14483 272402 15459 272436
rect 14390 272306 14424 272374
rect 15518 272306 15552 272374
rect 14483 272244 15459 272278
rect 14390 272148 14424 272216
rect 15518 272148 15552 272216
rect 15930 273096 15964 273164
rect 17058 273096 17092 273164
rect 16023 273034 16999 273068
rect 15930 272938 15964 273006
rect 17058 272938 17092 273006
rect 16023 272876 16999 272910
rect 15930 272780 15964 272848
rect 17058 272780 17092 272848
rect 16023 272718 16999 272752
rect 15930 272622 15964 272690
rect 17058 272622 17092 272690
rect 16023 272560 16999 272594
rect 15930 272464 15964 272532
rect 17058 272464 17092 272532
rect 16023 272402 16999 272436
rect 15930 272306 15964 272374
rect 17058 272306 17092 272374
rect 16023 272244 16999 272278
rect 14483 272086 15459 272120
rect 14390 271990 14424 272058
rect 15518 271990 15552 272058
rect 14483 271928 15459 271962
rect 14390 271832 14424 271900
rect 15518 271832 15552 271900
rect 14483 271770 15459 271804
rect 14390 271674 14424 271742
rect 15518 271674 15552 271742
rect 14483 271612 15459 271646
rect 15620 271640 15654 272210
rect 15654 271640 15828 272210
rect 15828 271640 15860 272210
rect 15930 272148 15964 272216
rect 17058 272148 17092 272216
rect 16023 272086 16999 272120
rect 15930 271990 15964 272058
rect 17058 271990 17092 272058
rect 16023 271928 16999 271962
rect 15930 271832 15964 271900
rect 17058 271832 17092 271900
rect 16023 271770 16999 271804
rect 15930 271674 15964 271742
rect 17058 271674 17092 271742
rect 14390 271516 14424 271584
rect 15518 271516 15552 271584
rect 14483 271454 15459 271488
rect 14390 271358 14424 271426
rect 15518 271358 15552 271426
rect 14483 271296 15459 271330
rect 14390 271200 14424 271268
rect 15518 271200 15552 271268
rect 14483 271138 15459 271172
rect 14390 271042 14424 271110
rect 15518 271042 15552 271110
rect 14483 270980 15459 271014
rect 16023 271612 16999 271646
rect 15930 271516 15964 271584
rect 17058 271516 17092 271584
rect 16023 271454 16999 271488
rect 15930 271358 15964 271426
rect 17058 271358 17092 271426
rect 16023 271296 16999 271330
rect 15930 271200 15964 271268
rect 17058 271200 17092 271268
rect 16023 271138 16999 271172
rect 15930 271042 15964 271110
rect 17058 271042 17092 271110
rect 16023 270980 16999 271014
rect 20632 274186 21608 274220
rect 20548 273990 20582 274158
rect 21658 273990 21692 274158
rect 20632 273928 21608 273962
rect 20548 273732 20582 273900
rect 21658 273732 21692 273900
rect 20632 273670 21608 273704
rect 17591 273187 18567 273221
rect 17507 273091 17541 273159
rect 18617 273091 18651 273159
rect 17591 273029 18567 273063
rect 17405 272326 17439 272976
rect 17507 272933 17541 273001
rect 18617 272933 18651 273001
rect 17591 272871 18567 272905
rect 17507 272775 17541 272843
rect 18617 272775 18651 272843
rect 17591 272713 18567 272747
rect 17507 272617 17541 272685
rect 18617 272617 18651 272685
rect 17591 272555 18567 272589
rect 17507 272459 17541 272527
rect 18617 272459 18651 272527
rect 17591 272397 18567 272431
rect 17507 272301 17541 272369
rect 18617 272301 18651 272369
rect 18719 272326 18753 272976
rect 17591 272239 18567 272273
rect 17507 272143 17541 272211
rect 18617 272143 18651 272211
rect 17591 272081 18567 272115
rect 19111 273187 20087 273221
rect 19027 273091 19061 273159
rect 20137 273091 20171 273159
rect 19111 273029 20087 273063
rect 18925 272326 18959 272976
rect 19027 272933 19061 273001
rect 20137 272933 20171 273001
rect 19111 272871 20087 272905
rect 19027 272775 19061 272843
rect 20137 272775 20171 272843
rect 19111 272713 20087 272747
rect 19027 272617 19061 272685
rect 20137 272617 20171 272685
rect 19111 272555 20087 272589
rect 19027 272459 19061 272527
rect 20137 272459 20171 272527
rect 19111 272397 20087 272431
rect 19027 272301 19061 272369
rect 20137 272301 20171 272369
rect 20239 272326 20273 272976
rect 19111 272239 20087 272273
rect 19027 272143 19061 272211
rect 20137 272143 20171 272211
rect 19111 272081 20087 272115
rect 20446 271833 20480 273477
rect 20548 273474 20582 273642
rect 21658 273474 21692 273642
rect 20632 273412 21608 273446
rect 20548 273216 20582 273384
rect 21658 273216 21692 273384
rect 20632 273154 21608 273188
rect 20548 272958 20582 273126
rect 21658 272958 21692 273126
rect 20632 272896 21608 272930
rect 20548 272700 20582 272868
rect 21658 272700 21692 272868
rect 20632 272638 21608 272672
rect 20548 272442 20582 272610
rect 21658 272442 21692 272610
rect 20632 272380 21608 272414
rect 20548 272184 20582 272352
rect 21658 272184 21692 272352
rect 20632 272122 21608 272156
rect 20548 271926 20582 272094
rect 21658 271926 21692 272094
rect 20632 271864 21608 271898
rect 20548 271668 20582 271836
rect 21658 271668 21692 271836
rect 21760 271833 21794 273477
rect 20632 271606 21608 271640
rect 20548 271410 20582 271578
rect 21658 271410 21692 271578
rect 20632 271348 21608 271382
rect 20548 271152 20582 271320
rect 21658 271152 21692 271320
rect 20632 271090 21608 271124
rect 22152 274442 23128 274476
rect 22068 274246 22102 274414
rect 23178 274246 23212 274414
rect 22152 274184 23128 274218
rect 22068 273988 22102 274156
rect 23178 273988 23212 274156
rect 22152 273926 23128 273960
rect 22068 273730 22102 273898
rect 23178 273730 23212 273898
rect 22152 273668 23128 273702
rect 21966 271702 22000 273604
rect 22068 273472 22102 273640
rect 23178 273472 23212 273640
rect 22152 273410 23128 273444
rect 22068 273214 22102 273382
rect 23178 273214 23212 273382
rect 22152 273152 23128 273186
rect 22068 272956 22102 273124
rect 23178 272956 23212 273124
rect 22152 272894 23128 272928
rect 22068 272698 22102 272866
rect 23178 272698 23212 272866
rect 22152 272636 23128 272670
rect 22068 272440 22102 272608
rect 23178 272440 23212 272608
rect 22152 272378 23128 272412
rect 22068 272182 22102 272350
rect 23178 272182 23212 272350
rect 22152 272120 23128 272154
rect 22068 271924 22102 272092
rect 23178 271924 23212 272092
rect 22152 271862 23128 271896
rect 22068 271666 22102 271834
rect 23178 271666 23212 271834
rect 23280 271702 23314 273604
rect 24570 273556 24800 273560
rect 26080 273556 26310 273560
rect 24570 273522 24800 273556
rect 24570 273520 24800 273522
rect 24193 273408 25169 273442
rect 24100 273212 24134 273380
rect 25228 273212 25262 273380
rect 24193 273150 25169 273184
rect 24100 272954 24134 273122
rect 25228 272954 25262 273122
rect 24193 272892 25169 272926
rect 24100 272696 24134 272864
rect 25228 272696 25262 272864
rect 24193 272634 25169 272668
rect 24100 272438 24134 272606
rect 25228 272438 25262 272606
rect 24193 272376 25169 272410
rect 24100 272180 24134 272348
rect 25228 272180 25262 272348
rect 24193 272118 25169 272152
rect 24100 271922 24134 272090
rect 25228 271922 25262 272090
rect 24193 271860 25169 271894
rect 24570 271746 24800 271780
rect 26080 273522 26310 273556
rect 26080 273520 26310 273522
rect 25693 273408 26669 273442
rect 25600 273212 25634 273380
rect 26728 273212 26762 273380
rect 25693 273150 26669 273184
rect 25600 272954 25634 273122
rect 26728 272954 26762 273122
rect 25693 272892 26669 272926
rect 25600 272696 25634 272864
rect 26728 272696 26762 272864
rect 25693 272634 26669 272668
rect 25600 272438 25634 272606
rect 26728 272438 26762 272606
rect 25693 272376 26669 272410
rect 25600 272180 25634 272348
rect 26728 272180 26762 272348
rect 25693 272118 26669 272152
rect 25600 271922 25634 272090
rect 26728 271922 26762 272090
rect 25693 271860 26669 271894
rect 28370 273280 28450 273300
rect 28370 273246 28450 273280
rect 28370 273220 28450 273246
rect 27420 272924 27650 272930
rect 27420 272890 27650 272924
rect 27302 272776 27778 272810
rect 27218 272680 27252 272748
rect 27828 272680 27862 272748
rect 27302 272618 27778 272652
rect 27218 272522 27252 272590
rect 27828 272522 27862 272590
rect 27302 272460 27778 272494
rect 27420 272346 27650 272380
rect 27420 272340 27650 272346
rect 28302 273132 28528 273166
rect 28218 272936 28252 273104
rect 28578 272936 28612 273104
rect 28302 272874 28528 272908
rect 28218 272678 28252 272846
rect 28578 272678 28612 272846
rect 29052 273393 30028 273427
rect 28968 273197 29002 273365
rect 30078 273197 30112 273365
rect 29052 273135 30028 273169
rect 28968 272939 29002 273107
rect 30078 272939 30112 273107
rect 29052 272877 30028 272911
rect 28302 272616 28528 272650
rect 28218 272420 28252 272588
rect 28578 272420 28612 272588
rect 28680 272500 28714 272740
rect 28714 272500 28720 272740
rect 28860 272500 28866 272740
rect 28866 272500 28900 272740
rect 28968 272681 29002 272849
rect 30078 272681 30112 272849
rect 29052 272619 30028 272653
rect 28302 272358 28528 272392
rect 28218 272162 28252 272330
rect 28578 272162 28612 272330
rect 28302 272100 28528 272134
rect 28370 272020 28460 272050
rect 28370 271986 28460 272020
rect 28370 271960 28460 271986
rect 26080 271746 26310 271780
rect 28968 272423 29002 272591
rect 30078 272423 30112 272591
rect 30180 272500 30214 272740
rect 30214 272500 30220 272740
rect 29052 272361 30028 272395
rect 28968 272165 29002 272333
rect 30078 272165 30112 272333
rect 29052 272103 30028 272137
rect 28968 271907 29002 272075
rect 30078 271907 30112 272075
rect 29052 271845 30028 271879
rect 24570 271740 24800 271746
rect 26080 271740 26310 271746
rect 22152 271604 23128 271638
rect 22068 271408 22102 271576
rect 23178 271408 23212 271576
rect 22152 271346 23128 271380
rect 22068 271150 22102 271318
rect 23178 271150 23212 271318
rect 22152 271088 23128 271122
rect 22068 270892 22102 271060
rect 23178 270892 23212 271060
rect 22152 270830 23128 270864
rect 537364 271938 537484 272058
rect 543734 271938 543854 272058
rect 31020 269200 31260 269440
rect 32740 269200 32980 269440
rect 34460 269200 34700 269440
rect 35940 269200 36180 269440
rect 37660 269200 37900 269440
rect 39260 269200 39500 269440
rect 40980 269200 41220 269440
rect 42580 269200 42820 269440
rect 44300 269200 44540 269440
rect 537364 268938 537484 269058
rect 543734 268938 543854 269058
rect 11887 268142 13001 268539
rect 11887 265711 13001 266108
rect 13347 268142 14461 268539
rect 537777 267356 538891 267753
rect 539297 267356 540411 267753
rect 540807 267362 541921 267759
rect 542317 267362 543431 267759
rect 14540 267120 14573 267300
rect 14573 267120 14607 267300
rect 14607 267120 14640 267300
rect 14540 266700 14573 266880
rect 14573 266700 14607 266880
rect 14607 266700 14640 266880
rect 13347 265711 14461 266108
rect 8420 252444 13560 252478
rect 6002 252330 15978 252364
rect 5918 252281 5952 252315
rect 6002 252232 15978 252266
rect 16028 252183 16062 252217
rect 6002 252134 15978 252168
rect 5918 252085 5952 252119
rect 6002 252036 15978 252070
rect 16028 251987 16062 252021
rect 6002 251938 15978 251972
rect 5918 251889 5952 251923
rect 6002 251840 15978 251874
rect 16028 251791 16062 251825
rect 6002 251742 15978 251776
rect 5918 251693 5952 251727
rect 6002 251644 15978 251678
rect 16028 251595 16062 251629
rect 6002 251546 15978 251580
rect 16130 251564 16164 252150
rect 5918 251497 5952 251531
rect 6002 251448 15978 251482
rect 16028 251399 16062 251433
rect 6002 251350 15978 251384
rect 8420 251236 13560 251270
rect 8420 242044 13560 242078
rect 6002 241930 15978 241964
rect 5918 241881 5952 241915
rect 6002 241832 15978 241866
rect 16028 241783 16062 241817
rect 6002 241734 15978 241768
rect 5918 241685 5952 241719
rect 6002 241636 15978 241670
rect 16028 241587 16062 241621
rect 6002 241538 15978 241572
rect 5918 241489 5952 241523
rect 6002 241440 15978 241474
rect 16028 241391 16062 241425
rect 6002 241342 15978 241376
rect 5918 241293 5952 241327
rect 6002 241244 15978 241278
rect 16028 241195 16062 241229
rect 6002 241146 15978 241180
rect 16130 241164 16164 241750
rect 5918 241097 5952 241131
rect 6002 241048 15978 241082
rect 16028 240999 16062 241033
rect 6002 240950 15978 240984
rect 8420 240836 13560 240870
<< metal1 >>
rect 65040 702260 65940 702300
rect 23380 702180 24340 702200
rect 23380 702060 23400 702180
rect 23520 702060 23600 702180
rect 23720 702060 23800 702180
rect 23920 702060 24000 702180
rect 24120 702060 24200 702180
rect 24320 702060 24340 702180
rect 23380 702040 24340 702060
rect 65040 702080 65060 702260
rect 65240 702080 65400 702260
rect 65580 702080 65740 702260
rect 65920 702080 65940 702260
rect 573240 702240 574140 702280
rect 65040 702040 65940 702080
rect 563800 702120 565120 702160
rect 563800 702020 563840 702120
rect 563940 702020 563980 702120
rect 564080 702020 564120 702120
rect 564220 702020 564260 702120
rect 564360 702020 564400 702120
rect 564500 702020 564540 702120
rect 564640 702020 564680 702120
rect 564780 702020 564820 702120
rect 564920 702020 564960 702120
rect 565060 702020 565120 702120
rect 563800 701980 565120 702020
rect 563800 701880 563840 701980
rect 563940 701880 563980 701980
rect 564080 701880 564120 701980
rect 564220 701880 564260 701980
rect 564360 701880 564400 701980
rect 564500 701880 564540 701980
rect 564640 701880 564680 701980
rect 564780 701880 564820 701980
rect 564920 701880 564960 701980
rect 565060 701880 565120 701980
rect 563800 701840 565120 701880
rect 573240 702140 573280 702240
rect 573380 702140 573420 702240
rect 573520 702140 573560 702240
rect 573660 702140 573700 702240
rect 573800 702140 573840 702240
rect 573940 702140 573980 702240
rect 574080 702140 574140 702240
rect 573240 701980 574140 702140
rect 573240 701880 573280 701980
rect 573380 701880 573420 701980
rect 573520 701880 573560 701980
rect 573660 701880 573700 701980
rect 573800 701880 573840 701980
rect 573940 701880 573980 701980
rect 574080 701880 574140 701980
rect 573240 701840 574140 701880
rect 565040 699740 573080 700240
rect 24440 693020 24600 693060
rect 24440 692900 24460 693020
rect 24580 692900 24600 693020
rect 24440 692840 24600 692900
rect 24440 692720 24460 692840
rect 24580 692720 24600 692840
rect 24440 692660 24600 692720
rect 24440 692540 24460 692660
rect 24580 692540 24600 692660
rect 64680 693000 64880 693040
rect 64680 692860 64720 693000
rect 64860 692860 64880 693000
rect 64680 692800 64880 692860
rect 64680 692660 64720 692800
rect 64860 692660 64880 692800
rect 64680 692620 64880 692660
rect 66040 693000 66240 693040
rect 66040 692860 66060 693000
rect 66200 692860 66240 693000
rect 66040 692800 66240 692860
rect 66040 692660 66060 692800
rect 66200 692660 66240 692800
rect 66040 692620 66240 692660
rect 75080 693000 75280 693040
rect 75080 692860 75120 693000
rect 75260 692860 75280 693000
rect 75080 692800 75280 692860
rect 75080 692660 75120 692800
rect 75260 692660 75280 692800
rect 75080 692620 75280 692660
rect 24440 692480 24600 692540
rect 24440 692360 24460 692480
rect 24580 692360 24600 692480
rect 24440 692300 24600 692360
rect 24440 692180 24460 692300
rect 24580 692180 24600 692300
rect 12800 691900 14120 691980
rect 12800 691700 12900 691900
rect 13100 691700 13200 691900
rect 13400 691700 13500 691900
rect 13700 691700 13800 691900
rect 14000 691700 14120 691900
rect 75220 691820 76500 691980
rect 12800 691600 14120 691700
rect 566260 691100 571840 691320
rect 566260 690900 566300 691100
rect 566500 690900 566700 691100
rect 566900 690900 567100 691100
rect 567300 690900 567500 691100
rect 567700 690900 567900 691100
rect 568100 690900 568300 691100
rect 568500 690900 568700 691100
rect 568900 690900 569100 691100
rect 569300 690900 569500 691100
rect 569700 690900 569900 691100
rect 570100 690900 570300 691100
rect 570500 690900 570700 691100
rect 570900 690900 571100 691100
rect 571300 690900 571500 691100
rect 571700 690900 571840 691100
rect 566260 690700 571840 690900
rect 566260 690500 566300 690700
rect 566500 690500 566700 690700
rect 566900 690500 567100 690700
rect 567300 690500 567500 690700
rect 567700 690500 567900 690700
rect 568100 690500 568300 690700
rect 568500 690500 568700 690700
rect 568900 690500 569100 690700
rect 569300 690500 569500 690700
rect 569700 690500 569900 690700
rect 570100 690500 570300 690700
rect 570500 690500 570700 690700
rect 570900 690500 571100 690700
rect 571300 690500 571500 690700
rect 571700 690500 571840 690700
rect 47100 690300 47400 690400
rect 47100 690200 47200 690300
rect 47300 690200 47400 690300
rect 47100 690010 47400 690200
rect 43870 689830 43950 690010
rect 45350 690000 47400 690010
rect 45350 689830 47200 690000
rect 47100 689800 47200 689830
rect 47300 689800 47400 690000
rect 47100 689600 47400 689800
rect 47100 689500 47200 689600
rect 47300 689500 47400 689600
rect 47100 689400 47400 689500
rect 566260 690300 571840 690500
rect 566260 690100 566300 690300
rect 566500 690100 566700 690300
rect 566900 690100 567100 690300
rect 567300 690100 567500 690300
rect 567700 690100 567900 690300
rect 568100 690100 568300 690300
rect 568500 690100 568700 690300
rect 568900 690100 569100 690300
rect 569300 690100 569500 690300
rect 569700 690100 569900 690300
rect 570100 690100 570300 690300
rect 570500 690100 570700 690300
rect 570900 690100 571100 690300
rect 571300 690100 571500 690300
rect 571700 690100 571840 690300
rect 566260 689900 571840 690100
rect 566260 689700 566300 689900
rect 566500 689700 566700 689900
rect 566900 689700 567100 689900
rect 567300 689700 567500 689900
rect 567700 689700 567900 689900
rect 568100 689700 568300 689900
rect 568500 689700 568700 689900
rect 568900 689700 569100 689900
rect 569300 689700 569500 689900
rect 569700 689700 569900 689900
rect 570100 689700 570300 689900
rect 570500 689700 570700 689900
rect 570900 689700 571100 689900
rect 571300 689700 571500 689900
rect 571700 689700 571840 689900
rect 566260 689520 571840 689700
rect 566260 689500 571820 689520
rect 566260 689300 566300 689500
rect 566500 689300 566700 689500
rect 566900 689300 567100 689500
rect 567300 689300 567500 689500
rect 567700 689300 567900 689500
rect 568100 689300 568300 689500
rect 568500 689300 568700 689500
rect 568900 689300 569100 689500
rect 569300 689300 569500 689500
rect 569700 689300 569900 689500
rect 570100 689300 570300 689500
rect 570500 689300 570700 689500
rect 570900 689300 571100 689500
rect 571300 689300 571500 689500
rect 571700 689300 571820 689500
rect 41900 688700 42200 688800
rect 41900 688600 42000 688700
rect 42100 688600 42200 688700
rect 41900 688500 42200 688600
rect 41900 688300 42000 688500
rect 42100 688490 42200 688500
rect 42100 688310 43870 688490
rect 42100 688300 42200 688310
rect 41900 688200 42200 688300
rect 41900 688100 42000 688200
rect 42100 688100 42200 688200
rect 41900 688000 42200 688100
rect 566260 685080 571820 689300
rect 548820 684860 571820 685080
rect 582320 684600 582660 684660
rect 548820 684360 554960 684580
rect 554420 682300 554960 684360
rect 582320 684520 582360 684600
rect 582440 684520 582540 684600
rect 582620 684520 582660 684600
rect 582320 684440 582660 684520
rect 582320 684360 582360 684440
rect 582440 684360 582540 684440
rect 582620 684360 582660 684440
rect 582320 684280 582660 684360
rect 582320 684200 582360 684280
rect 582440 684200 582540 684280
rect 582620 684200 582660 684280
rect 582320 684100 582660 684200
rect 582320 684020 582360 684100
rect 582440 684020 582540 684100
rect 582620 684020 582660 684100
rect 582320 683940 582660 684020
rect 582320 683860 582360 683940
rect 582440 683860 582540 683940
rect 582620 683860 582660 683940
rect 582320 683740 582660 683860
rect 554420 682200 563740 682300
rect 554420 682000 561700 682200
rect 561900 682000 562100 682200
rect 562300 682000 562500 682200
rect 562700 682000 562900 682200
rect 563100 682000 563300 682200
rect 563500 682000 563740 682200
rect 554420 681800 563740 682000
rect 554420 681600 561700 681800
rect 561900 681600 562100 681800
rect 562300 681600 562500 681800
rect 562700 681600 562900 681800
rect 563100 681600 563300 681800
rect 563500 681600 563740 681800
rect 554420 681400 563740 681600
rect 554420 681200 561700 681400
rect 561900 681200 562100 681400
rect 562300 681200 562500 681400
rect 562700 681200 562900 681400
rect 563100 681200 563300 681400
rect 563500 681200 563740 681400
rect 554420 681000 563740 681200
rect 554420 680800 561700 681000
rect 561900 680800 562100 681000
rect 562300 680800 562500 681000
rect 562700 680800 562900 681000
rect 563100 680800 563300 681000
rect 563500 680800 563740 681000
rect 554420 680600 563740 680800
rect 554420 680400 561700 680600
rect 561900 680400 562100 680600
rect 562300 680400 562500 680600
rect 562700 680400 562900 680600
rect 563100 680400 563300 680600
rect 563500 680400 563740 680600
rect 554420 680200 563740 680400
rect 554420 680000 561700 680200
rect 561900 680000 562100 680200
rect 562300 680000 562500 680200
rect 562700 680000 562900 680200
rect 563100 680000 563300 680200
rect 563500 680000 563740 680200
rect 554420 679800 563740 680000
rect 554420 679600 561700 679800
rect 561900 679600 562100 679800
rect 562300 679600 562500 679800
rect 562700 679600 562900 679800
rect 563100 679600 563300 679800
rect 563500 679600 563740 679800
rect 554420 679400 563740 679600
rect 554420 679200 561700 679400
rect 561900 679200 562100 679400
rect 562300 679200 562500 679400
rect 562700 679200 562900 679400
rect 563100 679200 563300 679400
rect 563500 679200 563740 679400
rect 554420 679000 563740 679200
rect 554420 678800 561700 679000
rect 561900 678800 562100 679000
rect 562300 678800 562500 679000
rect 562700 678800 562900 679000
rect 563100 678800 563300 679000
rect 563500 678800 563740 679000
rect 554420 678600 563740 678800
rect 554420 678400 561700 678600
rect 561900 678400 562100 678600
rect 562300 678400 562500 678600
rect 562700 678400 562900 678600
rect 563100 678400 563300 678600
rect 563500 678400 563740 678600
rect 554420 678340 563740 678400
rect 571800 677350 572390 683650
rect 571800 677300 572280 677350
rect 571800 677100 571900 677300
rect 572100 677100 572280 677300
rect 571800 677000 572280 677100
rect 571800 676800 571900 677000
rect 572100 676800 572280 677000
rect 571800 676700 572280 676800
rect 571800 676500 571900 676700
rect 572100 676500 572280 676700
rect 571800 676400 572280 676500
rect 571800 676200 571900 676400
rect 572100 676200 572280 676400
rect 571800 676100 572280 676200
rect 32600 663300 48300 663400
rect 32600 663000 32800 663300
rect 33100 663000 33300 663300
rect 33600 663000 33800 663300
rect 34100 663000 34300 663300
rect 34600 663000 34800 663300
rect 35100 663000 35300 663300
rect 35600 663000 35800 663300
rect 36100 663000 36300 663300
rect 36600 663000 36800 663300
rect 37100 663000 37300 663300
rect 37600 663000 37800 663300
rect 38100 663000 38300 663300
rect 38600 663000 38800 663300
rect 39100 663000 39300 663300
rect 39600 663000 39800 663300
rect 40100 663000 40300 663300
rect 40600 663000 48300 663300
rect 32600 662800 48300 663000
rect 569240 306240 570140 306280
rect 559800 306120 561120 306160
rect 559800 306020 559840 306120
rect 559940 306020 559980 306120
rect 560080 306020 560120 306120
rect 560220 306020 560260 306120
rect 560360 306020 560400 306120
rect 560500 306020 560540 306120
rect 560640 306020 560680 306120
rect 560780 306020 560820 306120
rect 560920 306020 560960 306120
rect 561060 306020 561120 306120
rect 559800 305980 561120 306020
rect 559800 305880 559840 305980
rect 559940 305880 559980 305980
rect 560080 305882 560120 305980
rect 560080 305880 560097 305882
rect 560220 305880 560260 305980
rect 560360 305880 560400 305980
rect 560500 305882 560540 305980
rect 560523 305880 560540 305882
rect 560640 305880 560680 305980
rect 560780 305880 560820 305980
rect 560920 305880 560960 305980
rect 561060 305880 561120 305980
rect 569240 306140 569280 306240
rect 569380 306140 569420 306240
rect 569520 306140 569560 306240
rect 569660 306140 569700 306240
rect 569800 306140 569840 306240
rect 569940 306140 569980 306240
rect 570080 306140 570140 306240
rect 569240 305980 570140 306140
rect 559800 305848 560097 305880
rect 560131 305848 560293 305880
rect 560327 305848 560489 305880
rect 560523 305848 560685 305880
rect 560719 305848 560881 305880
rect 560915 305848 561120 305880
rect 559800 305840 561120 305848
rect 16020 304490 16180 304500
rect 5900 304478 16180 304490
rect 5900 304444 8420 304478
rect 13560 304444 16180 304478
rect 5900 304440 16180 304444
rect 8408 304438 13572 304440
rect 9680 304380 9740 304390
rect 5990 304364 9680 304370
rect 9845 304380 9905 304390
rect 9740 304364 9845 304370
rect 10045 304380 10105 304390
rect 9905 304364 10045 304370
rect 10235 304380 10295 304390
rect 10105 304364 10235 304370
rect 10415 304380 10475 304390
rect 10295 304364 10415 304370
rect 10615 304380 10675 304390
rect 10475 304364 10615 304370
rect 10805 304380 10865 304390
rect 10675 304364 10805 304370
rect 10965 304380 11025 304390
rect 10865 304364 10965 304370
rect 11155 304380 11215 304390
rect 11025 304364 11155 304370
rect 11330 304380 11390 304390
rect 11215 304364 11330 304370
rect 11470 304380 11530 304390
rect 11390 304364 11470 304370
rect 11530 304364 15990 304370
rect 5990 304330 6002 304364
rect 15978 304330 15990 304364
rect 5910 304327 5950 304330
rect 5910 304315 5958 304327
rect 5990 304324 9680 304330
rect 5910 304281 5918 304315
rect 5952 304281 5958 304315
rect 9740 304324 9845 304330
rect 9680 304310 9740 304320
rect 9905 304324 10045 304330
rect 9845 304310 9905 304320
rect 10105 304324 10235 304330
rect 10045 304310 10105 304320
rect 10295 304324 10415 304330
rect 10235 304310 10295 304320
rect 10475 304324 10615 304330
rect 10415 304310 10475 304320
rect 10675 304324 10805 304330
rect 10615 304310 10675 304320
rect 10865 304324 10965 304330
rect 10805 304310 10865 304320
rect 11025 304324 11155 304330
rect 10965 304310 11025 304320
rect 11215 304324 11330 304330
rect 11155 304310 11215 304320
rect 11390 304324 11470 304330
rect 11330 304310 11390 304320
rect 11530 304324 15990 304330
rect 11470 304310 11530 304320
rect 5910 304270 5958 304281
rect 16020 304280 16180 304440
rect 15970 304272 16180 304280
rect 5990 304270 16180 304272
rect 5910 304266 16180 304270
rect 5910 304232 6002 304266
rect 15978 304232 16180 304266
rect 5910 304226 16180 304232
rect 5910 304220 6000 304226
rect 15970 304220 16180 304226
rect 5910 304131 5950 304220
rect 16020 304217 16180 304220
rect 9680 304180 9740 304190
rect 5990 304168 9680 304174
rect 9845 304180 9905 304190
rect 9740 304168 9845 304174
rect 10045 304180 10105 304190
rect 9905 304168 10045 304174
rect 10235 304180 10295 304190
rect 10105 304168 10235 304174
rect 10415 304180 10475 304190
rect 10295 304168 10415 304174
rect 10615 304180 10675 304190
rect 10475 304168 10615 304174
rect 10805 304180 10865 304190
rect 10675 304168 10805 304174
rect 10965 304180 11025 304190
rect 10865 304168 10965 304174
rect 11155 304180 11215 304190
rect 11025 304168 11155 304174
rect 11330 304180 11390 304190
rect 11215 304168 11330 304174
rect 11470 304180 11530 304190
rect 11390 304168 11470 304174
rect 16020 304183 16028 304217
rect 16062 304183 16180 304217
rect 11530 304168 15990 304174
rect 5990 304134 6002 304168
rect 15978 304134 15990 304168
rect 5910 304119 5958 304131
rect 5990 304128 9680 304134
rect 5910 304085 5918 304119
rect 5952 304085 5958 304119
rect 9740 304128 9845 304134
rect 9680 304110 9740 304120
rect 9905 304128 10045 304134
rect 9845 304110 9905 304120
rect 10105 304128 10235 304134
rect 10045 304110 10105 304120
rect 10295 304128 10415 304134
rect 10235 304110 10295 304120
rect 10475 304128 10615 304134
rect 10415 304110 10475 304120
rect 10675 304128 10805 304134
rect 10615 304110 10675 304120
rect 10865 304128 10965 304134
rect 10805 304110 10865 304120
rect 11025 304128 11155 304134
rect 10965 304110 11025 304120
rect 11215 304128 11330 304134
rect 11155 304110 11215 304120
rect 11390 304128 11470 304134
rect 11330 304110 11390 304120
rect 11530 304128 15990 304134
rect 16020 304150 16180 304183
rect 11470 304110 11530 304120
rect 5910 304080 5958 304085
rect 16020 304080 16130 304150
rect 5910 304076 6000 304080
rect 15970 304076 16130 304080
rect 5910 304070 16130 304076
rect 5910 304036 6002 304070
rect 15978 304036 16130 304070
rect 5910 304030 16130 304036
rect 5910 303935 5950 304030
rect 15970 304021 16130 304030
rect 15970 304020 16028 304021
rect 9680 303980 9740 303990
rect 5990 303972 9680 303978
rect 9845 303980 9905 303990
rect 9740 303972 9845 303978
rect 10045 303980 10105 303990
rect 9905 303972 10045 303978
rect 10235 303980 10295 303990
rect 10105 303972 10235 303978
rect 10415 303980 10475 303990
rect 10295 303972 10415 303978
rect 10615 303980 10675 303990
rect 10475 303972 10615 303978
rect 10805 303980 10865 303990
rect 10675 303972 10805 303978
rect 10965 303980 11025 303990
rect 10865 303972 10965 303978
rect 11155 303980 11215 303990
rect 11025 303972 11155 303978
rect 11330 303980 11390 303990
rect 11215 303972 11330 303978
rect 11470 303980 11530 303990
rect 11390 303972 11470 303978
rect 16020 303987 16028 304020
rect 16062 303987 16130 304021
rect 11530 303972 15990 303978
rect 5990 303938 6002 303972
rect 15978 303938 15990 303972
rect 5910 303923 5958 303935
rect 5990 303932 9680 303938
rect 5910 303889 5918 303923
rect 5952 303889 5958 303923
rect 9740 303932 9845 303938
rect 9680 303910 9740 303920
rect 9905 303932 10045 303938
rect 9845 303910 9905 303920
rect 10105 303932 10235 303938
rect 10045 303910 10105 303920
rect 10295 303932 10415 303938
rect 10235 303910 10295 303920
rect 10475 303932 10615 303938
rect 10415 303910 10475 303920
rect 10675 303932 10805 303938
rect 10615 303910 10675 303920
rect 10865 303932 10965 303938
rect 10805 303910 10865 303920
rect 11025 303932 11155 303938
rect 10965 303910 11025 303920
rect 11215 303932 11330 303938
rect 11155 303910 11215 303920
rect 11390 303932 11470 303938
rect 11330 303910 11390 303920
rect 11530 303932 15990 303938
rect 11470 303910 11530 303920
rect 16020 303890 16130 303987
rect 5910 303880 5958 303889
rect 15970 303880 16130 303890
rect 5910 303874 16130 303880
rect 5910 303840 6002 303874
rect 15978 303840 16130 303874
rect 5910 303834 16130 303840
rect 5910 303830 6000 303834
rect 15970 303830 16130 303834
rect 5910 303739 5950 303830
rect 16020 303825 16130 303830
rect 9680 303790 9740 303800
rect 5990 303776 9680 303782
rect 9845 303790 9905 303800
rect 9740 303776 9845 303782
rect 10045 303790 10105 303800
rect 9905 303776 10045 303782
rect 10235 303790 10295 303800
rect 10105 303776 10235 303782
rect 10415 303790 10475 303800
rect 10295 303776 10415 303782
rect 10615 303790 10675 303800
rect 10475 303776 10615 303782
rect 10805 303790 10865 303800
rect 10675 303776 10805 303782
rect 10965 303790 11025 303800
rect 10865 303776 10965 303782
rect 11155 303790 11215 303800
rect 11025 303776 11155 303782
rect 11330 303790 11390 303800
rect 11215 303776 11330 303782
rect 11470 303790 11530 303800
rect 11390 303776 11470 303782
rect 16020 303791 16028 303825
rect 16062 303791 16130 303825
rect 11530 303776 15990 303782
rect 5990 303742 6002 303776
rect 15978 303742 15990 303776
rect 5910 303727 5958 303739
rect 5990 303736 9680 303742
rect 5910 303693 5918 303727
rect 5952 303693 5958 303727
rect 9740 303736 9845 303742
rect 9680 303720 9740 303730
rect 9905 303736 10045 303742
rect 9845 303720 9905 303730
rect 10105 303736 10235 303742
rect 10045 303720 10105 303730
rect 10295 303736 10415 303742
rect 10235 303720 10295 303730
rect 10475 303736 10615 303742
rect 10415 303720 10475 303730
rect 10675 303736 10805 303742
rect 10615 303720 10675 303730
rect 10865 303736 10965 303742
rect 10805 303720 10865 303730
rect 11025 303736 11155 303742
rect 10965 303720 11025 303730
rect 11215 303736 11330 303742
rect 11155 303720 11215 303730
rect 11390 303736 11470 303742
rect 11330 303720 11390 303730
rect 11530 303736 15990 303742
rect 11470 303720 11530 303730
rect 5910 303690 5958 303693
rect 16020 303690 16130 303791
rect 5910 303684 6000 303690
rect 15970 303684 16130 303690
rect 5910 303678 16130 303684
rect 5910 303644 6002 303678
rect 15978 303644 16130 303678
rect 5910 303640 16130 303644
rect 5910 303543 5950 303640
rect 5990 303638 16130 303640
rect 15970 303630 16130 303638
rect 16020 303629 16130 303630
rect 9680 303590 9740 303600
rect 5990 303580 9680 303586
rect 9845 303590 9905 303600
rect 9740 303580 9845 303586
rect 10045 303590 10105 303600
rect 9905 303580 10045 303586
rect 10235 303590 10295 303600
rect 10105 303580 10235 303586
rect 10415 303590 10475 303600
rect 10295 303580 10415 303586
rect 10615 303590 10675 303600
rect 10475 303580 10615 303586
rect 10805 303590 10865 303600
rect 10675 303580 10805 303586
rect 10965 303590 11025 303600
rect 10865 303580 10965 303586
rect 11155 303590 11215 303600
rect 11025 303580 11155 303586
rect 11330 303590 11390 303600
rect 11215 303580 11330 303586
rect 11470 303590 11530 303600
rect 11390 303580 11470 303586
rect 16020 303595 16028 303629
rect 16062 303595 16130 303629
rect 11530 303580 15990 303586
rect 5990 303546 6002 303580
rect 15978 303546 15990 303580
rect 5910 303531 5958 303543
rect 5990 303540 9680 303546
rect 5910 303497 5918 303531
rect 5952 303497 5958 303531
rect 9740 303540 9845 303546
rect 9680 303520 9740 303530
rect 9905 303540 10045 303546
rect 9845 303520 9905 303530
rect 10105 303540 10235 303546
rect 10045 303520 10105 303530
rect 10295 303540 10415 303546
rect 10235 303520 10295 303530
rect 10475 303540 10615 303546
rect 10415 303520 10475 303530
rect 10675 303540 10805 303546
rect 10615 303520 10675 303530
rect 10865 303540 10965 303546
rect 10805 303520 10865 303530
rect 11025 303540 11155 303546
rect 10965 303520 11025 303530
rect 11215 303540 11330 303546
rect 11155 303520 11215 303530
rect 11390 303540 11470 303546
rect 11330 303520 11390 303530
rect 11530 303540 15990 303546
rect 16020 303564 16130 303595
rect 16164 303564 16180 304150
rect 11470 303520 11530 303530
rect 5910 303490 5958 303497
rect 16020 303490 16180 303564
rect 5910 303488 6000 303490
rect 15970 303488 16180 303490
rect 5910 303482 16180 303488
rect 5910 303448 6002 303482
rect 15978 303448 16180 303482
rect 5910 303442 16180 303448
rect 5910 303440 6000 303442
rect 15970 303440 16180 303442
rect 16020 303433 16180 303440
rect 9680 303400 9740 303410
rect 5990 303384 9680 303390
rect 9845 303390 9905 303400
rect 10045 303390 10105 303400
rect 10235 303390 10295 303400
rect 10415 303390 10475 303400
rect 10615 303390 10675 303400
rect 10805 303390 10865 303400
rect 10965 303390 11025 303400
rect 11155 303390 11215 303400
rect 11330 303390 11390 303400
rect 11470 303390 11530 303400
rect 16020 303399 16028 303433
rect 16062 303399 16180 303433
rect 9740 303384 9845 303390
rect 9905 303384 10045 303390
rect 10105 303384 10235 303390
rect 10295 303384 10415 303390
rect 10475 303384 10615 303390
rect 10675 303384 10805 303390
rect 10865 303384 10965 303390
rect 11025 303384 11155 303390
rect 11215 303384 11330 303390
rect 11390 303384 11470 303390
rect 11530 303384 15990 303390
rect 5990 303350 6002 303384
rect 15978 303350 15990 303384
rect 5990 303344 9680 303350
rect 9740 303344 9845 303350
rect 9680 303330 9740 303340
rect 9905 303344 10045 303350
rect 9845 303320 9905 303330
rect 10105 303344 10235 303350
rect 10045 303320 10105 303330
rect 10295 303344 10415 303350
rect 10235 303320 10295 303330
rect 10475 303344 10615 303350
rect 10415 303320 10475 303330
rect 10675 303344 10805 303350
rect 10615 303320 10675 303330
rect 10865 303344 10965 303350
rect 10805 303320 10865 303330
rect 11025 303344 11155 303350
rect 10965 303320 11025 303330
rect 11215 303344 11330 303350
rect 11155 303320 11215 303330
rect 11390 303344 11470 303350
rect 11330 303320 11390 303330
rect 11530 303344 15990 303350
rect 11470 303320 11530 303330
rect 16020 303280 16180 303399
rect 5900 303270 16180 303280
rect 5900 303236 8420 303270
rect 13560 303260 16180 303270
rect 13560 303236 15000 303260
rect 5900 303230 15000 303236
rect 14960 303120 15000 303230
rect 15140 303120 15200 303260
rect 15340 303230 16180 303260
rect 15340 303120 15380 303230
rect 16020 303220 16180 303230
rect 559830 303380 559880 305840
rect 14960 303080 15380 303120
rect 559830 298240 559836 303380
rect 559870 298240 559880 303380
rect 559944 305798 559990 305810
rect 560040 305800 560090 305840
rect 560240 305810 560290 305840
rect 559944 302120 559950 305798
rect 559984 302120 559990 305798
rect 560042 305798 560088 305800
rect 559930 302060 559940 302120
rect 560000 302060 560010 302120
rect 559944 301955 559950 302060
rect 559984 301955 559990 302060
rect 559920 301895 559930 301955
rect 559990 301895 560000 301955
rect 559944 301755 559950 301895
rect 559984 301755 559990 301895
rect 559920 301695 559930 301755
rect 559990 301695 560000 301755
rect 559944 301565 559950 301695
rect 559984 301565 559990 301695
rect 559920 301505 559930 301565
rect 559990 301505 560000 301565
rect 559944 301385 559950 301505
rect 559984 301385 559990 301505
rect 559920 301325 559930 301385
rect 559990 301325 560000 301385
rect 559944 301185 559950 301325
rect 559984 301185 559990 301325
rect 559920 301125 559930 301185
rect 559990 301125 560000 301185
rect 559944 300995 559950 301125
rect 559984 300995 559990 301125
rect 559920 300935 559930 300995
rect 559990 300935 560000 300995
rect 559944 300835 559950 300935
rect 559984 300835 559990 300935
rect 559920 300775 559930 300835
rect 559990 300775 560000 300835
rect 559944 300645 559950 300775
rect 559984 300645 559990 300775
rect 559920 300585 559930 300645
rect 559990 300585 560000 300645
rect 559944 300470 559950 300585
rect 559984 300470 559990 300585
rect 559920 300410 559930 300470
rect 559990 300410 560000 300470
rect 559944 300330 559950 300410
rect 559984 300330 559990 300410
rect 559920 300270 559930 300330
rect 559990 300270 560000 300330
rect 559830 295680 559880 298240
rect 559944 295822 559950 300270
rect 559984 295822 559990 300270
rect 560042 295830 560048 305798
rect 559944 295810 559990 295822
rect 560040 295822 560048 295830
rect 560082 295830 560088 305798
rect 560140 305798 560186 305810
rect 560140 302120 560146 305798
rect 560180 302120 560186 305798
rect 560238 305800 560290 305810
rect 560238 305798 560284 305800
rect 560120 302060 560130 302120
rect 560190 302060 560200 302120
rect 560140 301955 560146 302060
rect 560180 301955 560186 302060
rect 560120 301895 560130 301955
rect 560190 301895 560200 301955
rect 560140 301755 560146 301895
rect 560180 301755 560186 301895
rect 560120 301695 560130 301755
rect 560190 301695 560200 301755
rect 560140 301565 560146 301695
rect 560180 301565 560186 301695
rect 560120 301505 560130 301565
rect 560190 301505 560200 301565
rect 560140 301385 560146 301505
rect 560180 301385 560186 301505
rect 560120 301325 560130 301385
rect 560190 301325 560200 301385
rect 560140 301185 560146 301325
rect 560180 301185 560186 301325
rect 560120 301125 560130 301185
rect 560190 301125 560200 301185
rect 560140 300995 560146 301125
rect 560180 300995 560186 301125
rect 560120 300935 560130 300995
rect 560190 300935 560200 300995
rect 560140 300835 560146 300935
rect 560180 300835 560186 300935
rect 560120 300775 560130 300835
rect 560190 300775 560200 300835
rect 560140 300645 560146 300775
rect 560180 300645 560186 300775
rect 560120 300585 560130 300645
rect 560190 300585 560200 300645
rect 560140 300470 560146 300585
rect 560180 300470 560186 300585
rect 560120 300410 560130 300470
rect 560190 300410 560200 300470
rect 560140 300330 560146 300410
rect 560180 300330 560186 300410
rect 560120 300270 560130 300330
rect 560190 300270 560200 300330
rect 560082 295822 560090 295830
rect 560040 295780 560090 295822
rect 560140 295822 560146 300270
rect 560180 295822 560186 300270
rect 560238 295830 560244 305798
rect 560140 295810 560186 295822
rect 560230 295822 560244 295830
rect 560278 295830 560284 305798
rect 560336 305798 560382 305810
rect 560430 305800 560480 305840
rect 560336 302120 560342 305798
rect 560376 302120 560382 305798
rect 560434 305798 560480 305800
rect 560320 302060 560330 302120
rect 560390 302060 560400 302120
rect 560336 301955 560342 302060
rect 560376 301955 560382 302060
rect 560320 301895 560330 301955
rect 560390 301895 560400 301955
rect 560336 301755 560342 301895
rect 560376 301755 560382 301895
rect 560320 301695 560330 301755
rect 560390 301695 560400 301755
rect 560336 301565 560342 301695
rect 560376 301565 560382 301695
rect 560320 301505 560330 301565
rect 560390 301505 560400 301565
rect 560336 301385 560342 301505
rect 560376 301385 560382 301505
rect 560320 301325 560330 301385
rect 560390 301325 560400 301385
rect 560336 301185 560342 301325
rect 560376 301185 560382 301325
rect 560320 301125 560330 301185
rect 560390 301125 560400 301185
rect 560336 300995 560342 301125
rect 560376 300995 560382 301125
rect 560320 300935 560330 300995
rect 560390 300935 560400 300995
rect 560336 300835 560342 300935
rect 560376 300835 560382 300935
rect 560320 300775 560330 300835
rect 560390 300775 560400 300835
rect 560336 300645 560342 300775
rect 560376 300645 560382 300775
rect 560320 300585 560330 300645
rect 560390 300585 560400 300645
rect 560336 300470 560342 300585
rect 560376 300470 560382 300585
rect 560320 300410 560330 300470
rect 560390 300410 560400 300470
rect 560336 300330 560342 300410
rect 560376 300330 560382 300410
rect 560320 300270 560330 300330
rect 560390 300270 560400 300330
rect 560278 295822 560290 295830
rect 560230 295780 560290 295822
rect 560336 295822 560342 300270
rect 560376 295822 560382 300270
rect 560434 295830 560440 305798
rect 560336 295810 560382 295822
rect 560430 295822 560440 295830
rect 560474 295830 560480 305798
rect 560532 305798 560578 305810
rect 560532 302120 560538 305798
rect 560572 302120 560578 305798
rect 560630 305800 560680 305840
rect 560820 305810 560870 305840
rect 560630 305798 560676 305800
rect 560510 302060 560520 302120
rect 560580 302060 560590 302120
rect 560532 301955 560538 302060
rect 560572 301955 560578 302060
rect 560510 301895 560520 301955
rect 560580 301895 560590 301955
rect 560532 301755 560538 301895
rect 560572 301755 560578 301895
rect 560510 301695 560520 301755
rect 560580 301695 560590 301755
rect 560532 301565 560538 301695
rect 560572 301565 560578 301695
rect 560510 301505 560520 301565
rect 560580 301505 560590 301565
rect 560532 301385 560538 301505
rect 560572 301385 560578 301505
rect 560510 301325 560520 301385
rect 560580 301325 560590 301385
rect 560532 301185 560538 301325
rect 560572 301185 560578 301325
rect 560510 301125 560520 301185
rect 560580 301125 560590 301185
rect 560532 300995 560538 301125
rect 560572 300995 560578 301125
rect 560510 300935 560520 300995
rect 560580 300935 560590 300995
rect 560532 300835 560538 300935
rect 560572 300835 560578 300935
rect 560510 300775 560520 300835
rect 560580 300775 560590 300835
rect 560532 300645 560538 300775
rect 560572 300645 560578 300775
rect 560510 300585 560520 300645
rect 560580 300585 560590 300645
rect 560532 300470 560538 300585
rect 560572 300470 560578 300585
rect 560510 300410 560520 300470
rect 560580 300410 560590 300470
rect 560532 300330 560538 300410
rect 560572 300330 560578 300410
rect 560510 300270 560520 300330
rect 560580 300270 560590 300330
rect 560474 295822 560490 295830
rect 560430 295780 560490 295822
rect 560532 295822 560538 300270
rect 560572 295822 560578 300270
rect 560630 295830 560636 305798
rect 560532 295810 560578 295822
rect 560620 295822 560636 295830
rect 560670 295830 560676 305798
rect 560728 305798 560774 305810
rect 560820 305800 560872 305810
rect 560728 302120 560734 305798
rect 560768 302120 560774 305798
rect 560826 305798 560872 305800
rect 560710 302060 560720 302120
rect 560780 302060 560790 302120
rect 560728 301955 560734 302060
rect 560768 301955 560774 302060
rect 560710 301895 560720 301955
rect 560780 301895 560790 301955
rect 560728 301755 560734 301895
rect 560768 301755 560774 301895
rect 560710 301695 560720 301755
rect 560780 301695 560790 301755
rect 560728 301565 560734 301695
rect 560768 301565 560774 301695
rect 560710 301505 560720 301565
rect 560780 301505 560790 301565
rect 560728 301385 560734 301505
rect 560768 301385 560774 301505
rect 560710 301325 560720 301385
rect 560780 301325 560790 301385
rect 560728 301185 560734 301325
rect 560768 301185 560774 301325
rect 560710 301125 560720 301185
rect 560780 301125 560790 301185
rect 560728 300995 560734 301125
rect 560768 300995 560774 301125
rect 560710 300935 560720 300995
rect 560780 300935 560790 300995
rect 560728 300835 560734 300935
rect 560768 300835 560774 300935
rect 560710 300775 560720 300835
rect 560780 300775 560790 300835
rect 560728 300645 560734 300775
rect 560768 300645 560774 300775
rect 560710 300585 560720 300645
rect 560780 300585 560790 300645
rect 560728 300470 560734 300585
rect 560768 300470 560774 300585
rect 560710 300410 560720 300470
rect 560780 300410 560790 300470
rect 560728 300330 560734 300410
rect 560768 300330 560774 300410
rect 560710 300270 560720 300330
rect 560780 300270 560790 300330
rect 560670 295822 560680 295830
rect 560620 295780 560680 295822
rect 560728 295822 560734 300270
rect 560768 295822 560774 300270
rect 560826 295830 560832 305798
rect 560728 295810 560774 295822
rect 560820 295822 560832 295830
rect 560866 295830 560872 305798
rect 560924 305798 560970 305810
rect 560924 302120 560930 305798
rect 560964 302120 560970 305798
rect 561040 304240 561090 305840
rect 569030 304240 569080 305900
rect 569240 305880 569280 305980
rect 569380 305880 569420 305980
rect 569520 305882 569560 305980
rect 569527 305880 569560 305882
rect 569660 305882 569700 305980
rect 569660 305880 569689 305882
rect 569800 305880 569840 305980
rect 569940 305880 569980 305980
rect 570080 305882 570140 305980
rect 570080 305880 570081 305882
rect 569240 305848 569297 305880
rect 569331 305848 569493 305880
rect 569527 305848 569689 305880
rect 569723 305848 569885 305880
rect 569919 305848 570081 305880
rect 570115 305848 570140 305882
rect 569240 305840 570140 305848
rect 561040 303740 569080 304240
rect 561040 303392 561090 303740
rect 561038 303380 561090 303392
rect 560910 302060 560920 302120
rect 560980 302060 560990 302120
rect 560924 301955 560930 302060
rect 560964 301955 560970 302060
rect 560910 301895 560920 301955
rect 560980 301895 560990 301955
rect 560924 301755 560930 301895
rect 560964 301755 560970 301895
rect 560910 301695 560920 301755
rect 560980 301695 560990 301755
rect 560924 301565 560930 301695
rect 560964 301565 560970 301695
rect 560910 301505 560920 301565
rect 560980 301505 560990 301565
rect 560924 301385 560930 301505
rect 560964 301385 560970 301505
rect 560910 301325 560920 301385
rect 560980 301325 560990 301385
rect 560924 301185 560930 301325
rect 560964 301185 560970 301325
rect 560910 301125 560920 301185
rect 560980 301125 560990 301185
rect 560924 300995 560930 301125
rect 560964 300995 560970 301125
rect 560910 300935 560920 300995
rect 560980 300935 560990 300995
rect 560924 300835 560930 300935
rect 560964 300835 560970 300935
rect 560910 300775 560920 300835
rect 560980 300775 560990 300835
rect 560924 300645 560930 300775
rect 560964 300645 560970 300775
rect 560910 300585 560920 300645
rect 560980 300585 560990 300645
rect 560924 300470 560930 300585
rect 560964 300470 560970 300585
rect 560910 300410 560920 300470
rect 560980 300410 560990 300470
rect 560924 300330 560930 300410
rect 560964 300330 560970 300410
rect 560910 300270 560920 300330
rect 560980 300270 560990 300330
rect 560866 295822 560880 295830
rect 560820 295780 560880 295822
rect 560924 295822 560930 300270
rect 560964 295822 560970 300270
rect 561038 298240 561044 303380
rect 561078 298240 561090 303380
rect 561038 298228 561090 298240
rect 560924 295810 560970 295822
rect 559980 295772 560880 295780
rect 559980 295740 559999 295772
rect 559987 295738 559999 295740
rect 560033 295740 560195 295772
rect 560033 295738 560045 295740
rect 559987 295732 560045 295738
rect 560183 295738 560195 295740
rect 560229 295740 560391 295772
rect 560229 295738 560241 295740
rect 560183 295732 560241 295738
rect 560379 295738 560391 295740
rect 560425 295740 560587 295772
rect 560425 295738 560437 295740
rect 560379 295732 560437 295738
rect 560575 295738 560587 295740
rect 560621 295740 560783 295772
rect 560621 295738 560633 295740
rect 560575 295732 560633 295738
rect 560771 295738 560783 295740
rect 560817 295740 560880 295772
rect 560817 295738 560829 295740
rect 560771 295732 560829 295738
rect 561040 295680 561090 298228
rect 559830 295670 561090 295680
rect 559830 295636 560164 295670
rect 560750 295636 561090 295670
rect 559830 295630 561090 295636
rect 569030 303380 569080 303740
rect 569030 298240 569036 303380
rect 569070 298240 569080 303380
rect 569144 305798 569190 305810
rect 569240 305800 569290 305840
rect 569440 305810 569490 305840
rect 569144 302120 569150 305798
rect 569184 302120 569190 305798
rect 569242 305798 569288 305800
rect 569130 302060 569140 302120
rect 569200 302060 569210 302120
rect 569144 301955 569150 302060
rect 569184 301955 569190 302060
rect 569120 301895 569130 301955
rect 569190 301895 569200 301955
rect 569144 301755 569150 301895
rect 569184 301755 569190 301895
rect 569120 301695 569130 301755
rect 569190 301695 569200 301755
rect 569144 301565 569150 301695
rect 569184 301565 569190 301695
rect 569120 301505 569130 301565
rect 569190 301505 569200 301565
rect 569144 301385 569150 301505
rect 569184 301385 569190 301505
rect 569120 301325 569130 301385
rect 569190 301325 569200 301385
rect 569144 301185 569150 301325
rect 569184 301185 569190 301325
rect 569120 301125 569130 301185
rect 569190 301125 569200 301185
rect 569144 300995 569150 301125
rect 569184 300995 569190 301125
rect 569120 300935 569130 300995
rect 569190 300935 569200 300995
rect 569144 300835 569150 300935
rect 569184 300835 569190 300935
rect 569120 300775 569130 300835
rect 569190 300775 569200 300835
rect 569144 300645 569150 300775
rect 569184 300645 569190 300775
rect 569120 300585 569130 300645
rect 569190 300585 569200 300645
rect 569144 300470 569150 300585
rect 569184 300470 569190 300585
rect 569120 300410 569130 300470
rect 569190 300410 569200 300470
rect 569144 300330 569150 300410
rect 569184 300330 569190 300410
rect 569120 300270 569130 300330
rect 569190 300270 569200 300330
rect 569030 295680 569080 298240
rect 569144 295822 569150 300270
rect 569184 295822 569190 300270
rect 569242 295830 569248 305798
rect 569144 295810 569190 295822
rect 569240 295822 569248 295830
rect 569282 295830 569288 305798
rect 569340 305798 569386 305810
rect 569340 302120 569346 305798
rect 569380 302120 569386 305798
rect 569438 305800 569490 305810
rect 569438 305798 569484 305800
rect 569320 302060 569330 302120
rect 569390 302060 569400 302120
rect 569340 301955 569346 302060
rect 569380 301955 569386 302060
rect 569320 301895 569330 301955
rect 569390 301895 569400 301955
rect 569340 301755 569346 301895
rect 569380 301755 569386 301895
rect 569320 301695 569330 301755
rect 569390 301695 569400 301755
rect 569340 301565 569346 301695
rect 569380 301565 569386 301695
rect 569320 301505 569330 301565
rect 569390 301505 569400 301565
rect 569340 301385 569346 301505
rect 569380 301385 569386 301505
rect 569320 301325 569330 301385
rect 569390 301325 569400 301385
rect 569340 301185 569346 301325
rect 569380 301185 569386 301325
rect 569320 301125 569330 301185
rect 569390 301125 569400 301185
rect 569340 300995 569346 301125
rect 569380 300995 569386 301125
rect 569320 300935 569330 300995
rect 569390 300935 569400 300995
rect 569340 300835 569346 300935
rect 569380 300835 569386 300935
rect 569320 300775 569330 300835
rect 569390 300775 569400 300835
rect 569340 300645 569346 300775
rect 569380 300645 569386 300775
rect 569320 300585 569330 300645
rect 569390 300585 569400 300645
rect 569340 300470 569346 300585
rect 569380 300470 569386 300585
rect 569320 300410 569330 300470
rect 569390 300410 569400 300470
rect 569340 300330 569346 300410
rect 569380 300330 569386 300410
rect 569320 300270 569330 300330
rect 569390 300270 569400 300330
rect 569282 295822 569290 295830
rect 569240 295780 569290 295822
rect 569340 295822 569346 300270
rect 569380 295822 569386 300270
rect 569438 295830 569444 305798
rect 569340 295810 569386 295822
rect 569430 295822 569444 295830
rect 569478 295830 569484 305798
rect 569536 305798 569582 305810
rect 569630 305800 569680 305840
rect 569536 302120 569542 305798
rect 569576 302120 569582 305798
rect 569634 305798 569680 305800
rect 569520 302060 569530 302120
rect 569590 302060 569600 302120
rect 569536 301955 569542 302060
rect 569576 301955 569582 302060
rect 569520 301895 569530 301955
rect 569590 301895 569600 301955
rect 569536 301755 569542 301895
rect 569576 301755 569582 301895
rect 569520 301695 569530 301755
rect 569590 301695 569600 301755
rect 569536 301565 569542 301695
rect 569576 301565 569582 301695
rect 569520 301505 569530 301565
rect 569590 301505 569600 301565
rect 569536 301385 569542 301505
rect 569576 301385 569582 301505
rect 569520 301325 569530 301385
rect 569590 301325 569600 301385
rect 569536 301185 569542 301325
rect 569576 301185 569582 301325
rect 569520 301125 569530 301185
rect 569590 301125 569600 301185
rect 569536 300995 569542 301125
rect 569576 300995 569582 301125
rect 569520 300935 569530 300995
rect 569590 300935 569600 300995
rect 569536 300835 569542 300935
rect 569576 300835 569582 300935
rect 569520 300775 569530 300835
rect 569590 300775 569600 300835
rect 569536 300645 569542 300775
rect 569576 300645 569582 300775
rect 569520 300585 569530 300645
rect 569590 300585 569600 300645
rect 569536 300470 569542 300585
rect 569576 300470 569582 300585
rect 569520 300410 569530 300470
rect 569590 300410 569600 300470
rect 569536 300330 569542 300410
rect 569576 300330 569582 300410
rect 569520 300270 569530 300330
rect 569590 300270 569600 300330
rect 569478 295822 569490 295830
rect 569430 295780 569490 295822
rect 569536 295822 569542 300270
rect 569576 295822 569582 300270
rect 569634 295830 569640 305798
rect 569536 295810 569582 295822
rect 569630 295822 569640 295830
rect 569674 295830 569680 305798
rect 569732 305798 569778 305810
rect 569732 302120 569738 305798
rect 569772 302120 569778 305798
rect 569830 305800 569880 305840
rect 570020 305810 570070 305840
rect 569830 305798 569876 305800
rect 569710 302060 569720 302120
rect 569780 302060 569790 302120
rect 569732 301955 569738 302060
rect 569772 301955 569778 302060
rect 569710 301895 569720 301955
rect 569780 301895 569790 301955
rect 569732 301755 569738 301895
rect 569772 301755 569778 301895
rect 569710 301695 569720 301755
rect 569780 301695 569790 301755
rect 569732 301565 569738 301695
rect 569772 301565 569778 301695
rect 569710 301505 569720 301565
rect 569780 301505 569790 301565
rect 569732 301385 569738 301505
rect 569772 301385 569778 301505
rect 569710 301325 569720 301385
rect 569780 301325 569790 301385
rect 569732 301185 569738 301325
rect 569772 301185 569778 301325
rect 569710 301125 569720 301185
rect 569780 301125 569790 301185
rect 569732 300995 569738 301125
rect 569772 300995 569778 301125
rect 569710 300935 569720 300995
rect 569780 300935 569790 300995
rect 569732 300835 569738 300935
rect 569772 300835 569778 300935
rect 569710 300775 569720 300835
rect 569780 300775 569790 300835
rect 569732 300645 569738 300775
rect 569772 300645 569778 300775
rect 569710 300585 569720 300645
rect 569780 300585 569790 300645
rect 569732 300470 569738 300585
rect 569772 300470 569778 300585
rect 569710 300410 569720 300470
rect 569780 300410 569790 300470
rect 569732 300330 569738 300410
rect 569772 300330 569778 300410
rect 569710 300270 569720 300330
rect 569780 300270 569790 300330
rect 569674 295822 569690 295830
rect 569630 295780 569690 295822
rect 569732 295822 569738 300270
rect 569772 295822 569778 300270
rect 569830 295830 569836 305798
rect 569732 295810 569778 295822
rect 569820 295822 569836 295830
rect 569870 295830 569876 305798
rect 569928 305798 569974 305810
rect 570020 305800 570072 305810
rect 569928 302120 569934 305798
rect 569968 302120 569974 305798
rect 570026 305798 570072 305800
rect 569910 302060 569920 302120
rect 569980 302060 569990 302120
rect 569928 301955 569934 302060
rect 569968 301955 569974 302060
rect 569910 301895 569920 301955
rect 569980 301895 569990 301955
rect 569928 301755 569934 301895
rect 569968 301755 569974 301895
rect 569910 301695 569920 301755
rect 569980 301695 569990 301755
rect 569928 301565 569934 301695
rect 569968 301565 569974 301695
rect 569910 301505 569920 301565
rect 569980 301505 569990 301565
rect 569928 301385 569934 301505
rect 569968 301385 569974 301505
rect 569910 301325 569920 301385
rect 569980 301325 569990 301385
rect 569928 301185 569934 301325
rect 569968 301185 569974 301325
rect 569910 301125 569920 301185
rect 569980 301125 569990 301185
rect 569928 300995 569934 301125
rect 569968 300995 569974 301125
rect 569910 300935 569920 300995
rect 569980 300935 569990 300995
rect 569928 300835 569934 300935
rect 569968 300835 569974 300935
rect 569910 300775 569920 300835
rect 569980 300775 569990 300835
rect 569928 300645 569934 300775
rect 569968 300645 569974 300775
rect 569910 300585 569920 300645
rect 569980 300585 569990 300645
rect 569928 300470 569934 300585
rect 569968 300470 569974 300585
rect 569910 300410 569920 300470
rect 569980 300410 569990 300470
rect 569928 300330 569934 300410
rect 569968 300330 569974 300410
rect 569910 300270 569920 300330
rect 569980 300270 569990 300330
rect 569870 295822 569880 295830
rect 569820 295780 569880 295822
rect 569928 295822 569934 300270
rect 569968 295822 569974 300270
rect 570026 295830 570032 305798
rect 569928 295810 569974 295822
rect 570020 295822 570032 295830
rect 570066 295830 570072 305798
rect 570124 305798 570170 305810
rect 570124 302120 570130 305798
rect 570164 302120 570170 305798
rect 570240 303392 570290 305900
rect 570238 303380 570290 303392
rect 570110 302060 570120 302120
rect 570180 302060 570190 302120
rect 570124 301955 570130 302060
rect 570164 301955 570170 302060
rect 570110 301895 570120 301955
rect 570180 301895 570190 301955
rect 570124 301755 570130 301895
rect 570164 301755 570170 301895
rect 570110 301695 570120 301755
rect 570180 301695 570190 301755
rect 570124 301565 570130 301695
rect 570164 301565 570170 301695
rect 570110 301505 570120 301565
rect 570180 301505 570190 301565
rect 570124 301385 570130 301505
rect 570164 301385 570170 301505
rect 570110 301325 570120 301385
rect 570180 301325 570190 301385
rect 570124 301185 570130 301325
rect 570164 301185 570170 301325
rect 570110 301125 570120 301185
rect 570180 301125 570190 301185
rect 570124 300995 570130 301125
rect 570164 300995 570170 301125
rect 570110 300935 570120 300995
rect 570180 300935 570190 300995
rect 570124 300835 570130 300935
rect 570164 300835 570170 300935
rect 570110 300775 570120 300835
rect 570180 300775 570190 300835
rect 570124 300645 570130 300775
rect 570164 300645 570170 300775
rect 570110 300585 570120 300645
rect 570180 300585 570190 300645
rect 570124 300470 570130 300585
rect 570164 300470 570170 300585
rect 570110 300410 570120 300470
rect 570180 300410 570190 300470
rect 570124 300330 570130 300410
rect 570164 300330 570170 300410
rect 570110 300270 570120 300330
rect 570180 300270 570190 300330
rect 570066 295822 570080 295830
rect 570020 295780 570080 295822
rect 570124 295822 570130 300270
rect 570164 295822 570170 300270
rect 570238 298240 570244 303380
rect 570278 298240 570290 303380
rect 570238 298228 570290 298240
rect 570124 295810 570170 295822
rect 569180 295772 570080 295780
rect 569180 295740 569199 295772
rect 569187 295738 569199 295740
rect 569233 295740 569395 295772
rect 569233 295738 569245 295740
rect 569187 295732 569245 295738
rect 569383 295738 569395 295740
rect 569429 295740 569591 295772
rect 569429 295738 569441 295740
rect 569383 295732 569441 295738
rect 569579 295738 569591 295740
rect 569625 295740 569787 295772
rect 569625 295738 569637 295740
rect 569579 295732 569637 295738
rect 569775 295738 569787 295740
rect 569821 295740 569983 295772
rect 569821 295738 569833 295740
rect 569775 295732 569833 295738
rect 569971 295738 569983 295740
rect 570017 295740 570080 295772
rect 570017 295738 570029 295740
rect 569971 295732 570029 295738
rect 570240 295680 570290 298228
rect 569030 295670 570290 295680
rect 569030 295636 569364 295670
rect 569950 295636 570290 295670
rect 569030 295630 570290 295636
rect 562260 295100 567840 295320
rect 542907 294972 543011 294978
rect 537957 294962 538071 294968
rect 537957 294892 537969 294962
rect 538059 294892 538071 294962
rect 537957 294886 538071 294892
rect 538127 294962 538241 294968
rect 538127 294892 538139 294962
rect 538229 294892 538241 294962
rect 538127 294886 538241 294892
rect 540447 294962 540561 294968
rect 540447 294892 540459 294962
rect 540549 294892 540561 294962
rect 540447 294886 540561 294892
rect 540617 294962 540731 294968
rect 540617 294892 540629 294962
rect 540719 294892 540731 294962
rect 540617 294886 540731 294892
rect 542907 294892 542919 294972
rect 542999 294892 543011 294972
rect 542907 294886 543011 294892
rect 543077 294972 543181 294978
rect 543077 294892 543089 294972
rect 543169 294892 543181 294972
rect 543077 294886 543181 294892
rect 562260 294900 562300 295100
rect 562500 294900 562700 295100
rect 562900 294900 563100 295100
rect 563300 294900 563500 295100
rect 563700 294900 563900 295100
rect 564100 294900 564300 295100
rect 564500 294900 564700 295100
rect 564900 294900 565100 295100
rect 565300 294900 565500 295100
rect 565700 294900 565900 295100
rect 566100 294900 566300 295100
rect 566500 294900 566700 295100
rect 566900 294900 567100 295100
rect 567300 294900 567500 295100
rect 567700 294900 567840 295100
rect 537959 294802 537969 294852
rect 536359 294784 537969 294802
rect 538049 294802 538059 294852
rect 538129 294802 538139 294852
rect 538049 294784 538139 294802
rect 538219 294802 538229 294852
rect 540449 294802 540459 294852
rect 538219 294784 540459 294802
rect 540539 294802 540549 294852
rect 540619 294802 540629 294852
rect 540539 294784 540629 294802
rect 540709 294802 540719 294852
rect 542909 294802 542919 294842
rect 540709 294784 542919 294802
rect 542999 294802 543009 294842
rect 543079 294802 543089 294842
rect 542999 294784 543089 294802
rect 543169 294802 543179 294842
rect 543169 294784 544799 294802
rect 536359 294762 536380 294784
rect 536368 294750 536380 294762
rect 537356 294762 537616 294784
rect 537356 294750 537368 294762
rect 536368 294744 537368 294750
rect 537604 294750 537616 294762
rect 538592 294762 538852 294784
rect 538592 294750 538604 294762
rect 537604 294744 538604 294750
rect 538840 294750 538852 294762
rect 539828 294762 540088 294784
rect 539828 294750 539840 294762
rect 538840 294744 539840 294750
rect 540076 294750 540088 294762
rect 541064 294762 541324 294784
rect 541064 294750 541076 294762
rect 540076 294744 541076 294750
rect 541312 294750 541324 294762
rect 542300 294762 542560 294784
rect 543536 294762 543796 294784
rect 542300 294750 542312 294762
rect 541312 294744 542312 294750
rect 542548 294750 542560 294762
rect 543536 294750 543548 294762
rect 542548 294744 543548 294750
rect 543784 294750 543796 294762
rect 544772 294762 544799 294784
rect 544772 294750 544784 294762
rect 543784 294744 544784 294750
rect 536281 294722 536327 294734
rect 536281 294672 536287 294722
rect 536269 294654 536287 294672
rect 536321 294712 536327 294722
rect 537409 294722 537455 294734
rect 537517 294722 537563 294734
rect 537409 294712 537415 294722
rect 536321 294682 537415 294712
rect 536321 294654 537089 294682
rect 536269 294626 537089 294654
rect 537169 294626 537239 294682
rect 537319 294654 537415 294682
rect 537557 294712 537563 294722
rect 538645 294722 538691 294734
rect 538753 294722 538799 294734
rect 539881 294722 539927 294734
rect 539989 294722 540035 294734
rect 538645 294712 538651 294722
rect 537557 294654 538651 294712
rect 538793 294712 538799 294722
rect 539879 294712 539887 294722
rect 538793 294682 539887 294712
rect 538793 294654 539579 294682
rect 537319 294652 537419 294654
rect 537549 294652 538659 294654
rect 538789 294652 539579 294654
rect 537319 294626 539579 294652
rect 539659 294626 539729 294682
rect 539809 294654 539887 294682
rect 540029 294712 540035 294722
rect 541117 294722 541163 294734
rect 541225 294722 541271 294734
rect 541117 294712 541123 294722
rect 540029 294654 541123 294712
rect 541265 294712 541271 294722
rect 542353 294722 542399 294734
rect 542461 294722 542507 294734
rect 543589 294722 543635 294734
rect 543697 294722 543743 294734
rect 542353 294712 542359 294722
rect 541265 294682 542359 294712
rect 541265 294654 542059 294682
rect 539809 294652 539889 294654
rect 540019 294652 541129 294654
rect 541259 294652 542059 294654
rect 539809 294626 542059 294652
rect 542139 294626 542209 294682
rect 542289 294654 542359 294682
rect 542501 294712 542509 294722
rect 543589 294712 543595 294722
rect 542501 294654 543595 294712
rect 543737 294712 543743 294722
rect 544825 294722 544871 294734
rect 544825 294712 544831 294722
rect 543737 294654 544831 294712
rect 544865 294672 544871 294722
rect 562260 294700 567840 294900
rect 544865 294654 544879 294672
rect 542289 294652 542369 294654
rect 542499 294652 543599 294654
rect 543729 294652 544879 294654
rect 542289 294626 544879 294652
rect 536269 294592 536380 294626
rect 537356 294592 537616 294626
rect 538592 294592 538852 294626
rect 539828 294592 540088 294626
rect 541064 294592 541324 294626
rect 542300 294592 542560 294626
rect 543536 294592 543796 294626
rect 544772 294592 544879 294626
rect 536269 294572 536699 294592
rect 536689 294532 536699 294572
rect 536779 294572 536869 294592
rect 536779 294532 536789 294572
rect 536859 294532 536869 294572
rect 536949 294572 539219 294592
rect 536949 294532 536959 294572
rect 539209 294532 539219 294572
rect 539299 294572 539389 294592
rect 539299 294532 539309 294572
rect 539379 294532 539389 294572
rect 539469 294572 541709 294592
rect 539469 294532 539479 294572
rect 541699 294532 541709 294572
rect 541789 294572 541879 294592
rect 541789 294532 541799 294572
rect 541869 294532 541879 294572
rect 541959 294572 544159 294592
rect 541959 294532 541969 294572
rect 544149 294532 544159 294572
rect 544239 294572 544329 294592
rect 544239 294532 544249 294572
rect 544319 294532 544329 294572
rect 544409 294572 544879 294592
rect 544409 294532 544419 294572
rect 562260 294500 562300 294700
rect 562500 294500 562700 294700
rect 562900 294500 563100 294700
rect 563300 294500 563500 294700
rect 563700 294500 563900 294700
rect 564100 294500 564300 294700
rect 564500 294500 564700 294700
rect 564900 294500 565100 294700
rect 565300 294500 565500 294700
rect 565700 294500 565900 294700
rect 566100 294500 566300 294700
rect 566500 294500 566700 294700
rect 566900 294500 567100 294700
rect 567300 294500 567500 294700
rect 567700 294500 567840 294700
rect 537959 294262 537969 294312
rect 536359 294244 537969 294262
rect 538049 294262 538059 294312
rect 538129 294262 538139 294312
rect 538049 294244 538139 294262
rect 538219 294262 538229 294312
rect 540449 294262 540459 294312
rect 538219 294244 540459 294262
rect 540539 294262 540549 294312
rect 540619 294262 540629 294312
rect 540539 294244 540629 294262
rect 540709 294262 540719 294312
rect 542909 294262 542919 294302
rect 540709 294244 542919 294262
rect 542999 294262 543009 294302
rect 543079 294262 543089 294302
rect 542999 294244 543089 294262
rect 543169 294262 543179 294302
rect 562260 294300 567840 294500
rect 543169 294244 544799 294262
rect 14960 294200 15380 294240
rect 536359 294222 536380 294244
rect 536368 294210 536380 294222
rect 537356 294222 537616 294244
rect 537356 294210 537368 294222
rect 536368 294204 537368 294210
rect 537604 294210 537616 294222
rect 538592 294222 538852 294244
rect 538592 294210 538604 294222
rect 537604 294204 538604 294210
rect 538840 294210 538852 294222
rect 539828 294222 540088 294244
rect 539828 294210 539840 294222
rect 538840 294204 539840 294210
rect 540076 294210 540088 294222
rect 541064 294222 541324 294244
rect 541064 294210 541076 294222
rect 540076 294204 541076 294210
rect 541312 294210 541324 294222
rect 542300 294222 542560 294244
rect 543536 294222 543796 294244
rect 542300 294210 542312 294222
rect 541312 294204 542312 294210
rect 542548 294210 542560 294222
rect 543536 294210 543548 294222
rect 542548 294204 543548 294210
rect 543784 294210 543796 294222
rect 544772 294222 544799 294244
rect 544772 294210 544784 294222
rect 543784 294204 544784 294210
rect 14960 294090 15000 294200
rect 5900 294078 15000 294090
rect 5900 294044 8420 294078
rect 13560 294060 15000 294078
rect 15140 294060 15200 294200
rect 15340 294090 15380 294200
rect 536281 294182 536327 294194
rect 536281 294132 536287 294182
rect 536279 294114 536287 294132
rect 536321 294172 536327 294182
rect 537409 294182 537455 294194
rect 537517 294182 537563 294194
rect 537409 294172 537415 294182
rect 536321 294142 537415 294172
rect 536321 294114 537089 294142
rect 15340 294060 16170 294090
rect 13560 294044 16170 294060
rect 5900 294040 16170 294044
rect 8408 294038 13572 294040
rect 9680 293980 9740 293990
rect 5990 293964 9680 293970
rect 9845 293980 9905 293990
rect 9740 293964 9845 293970
rect 10045 293980 10105 293990
rect 9905 293964 10045 293970
rect 10235 293980 10295 293990
rect 10105 293964 10235 293970
rect 10415 293980 10475 293990
rect 10295 293964 10415 293970
rect 10615 293980 10675 293990
rect 10475 293964 10615 293970
rect 10805 293980 10865 293990
rect 10675 293964 10805 293970
rect 10965 293980 11025 293990
rect 10865 293964 10965 293970
rect 11155 293980 11215 293990
rect 11025 293964 11155 293970
rect 11330 293980 11390 293990
rect 11215 293964 11330 293970
rect 11470 293980 11530 293990
rect 11390 293964 11470 293970
rect 11530 293964 15990 293970
rect 5700 293920 5960 293940
rect 5990 293930 6002 293964
rect 15978 293930 15990 293964
rect 5990 293924 9680 293930
rect 5700 293740 5740 293920
rect 5920 293915 5960 293920
rect 5952 293881 5960 293915
rect 9740 293924 9845 293930
rect 9680 293910 9740 293920
rect 9905 293924 10045 293930
rect 9845 293910 9905 293920
rect 10105 293924 10235 293930
rect 10045 293910 10105 293920
rect 10295 293924 10415 293930
rect 10235 293910 10295 293920
rect 10475 293924 10615 293930
rect 10415 293910 10475 293920
rect 10675 293924 10805 293930
rect 10615 293910 10675 293920
rect 10865 293924 10965 293930
rect 10805 293910 10865 293920
rect 11025 293924 11155 293930
rect 10965 293910 11025 293920
rect 11215 293924 11330 293930
rect 11155 293910 11215 293920
rect 11390 293924 11470 293930
rect 11330 293910 11390 293920
rect 11530 293924 15990 293930
rect 11470 293910 11530 293920
rect 5920 293870 5960 293881
rect 15970 293872 16060 293880
rect 5990 293870 16060 293872
rect 5920 293866 16060 293870
rect 5920 293832 6002 293866
rect 15978 293832 16060 293866
rect 5920 293829 16060 293832
rect 5920 293826 16068 293829
rect 5920 293820 6000 293826
rect 15970 293820 16068 293826
rect 5920 293740 5960 293820
rect 16020 293817 16068 293820
rect 9680 293780 9740 293790
rect 5700 293719 5960 293740
rect 5990 293768 9680 293774
rect 9845 293780 9905 293790
rect 9740 293768 9845 293774
rect 10045 293780 10105 293790
rect 9905 293768 10045 293774
rect 10235 293780 10295 293790
rect 10105 293768 10235 293774
rect 10415 293780 10475 293790
rect 10295 293768 10415 293774
rect 10615 293780 10675 293790
rect 10475 293768 10615 293774
rect 10805 293780 10865 293790
rect 10675 293768 10805 293774
rect 10965 293780 11025 293790
rect 10865 293768 10965 293774
rect 11155 293780 11215 293790
rect 11025 293768 11155 293774
rect 11330 293780 11390 293790
rect 11215 293768 11330 293774
rect 11470 293780 11530 293790
rect 11390 293768 11470 293774
rect 16020 293783 16028 293817
rect 16062 293783 16068 293817
rect 11530 293768 15990 293774
rect 5990 293734 6002 293768
rect 15978 293734 15990 293768
rect 5990 293728 9680 293734
rect 5700 293685 5918 293719
rect 5952 293685 5960 293719
rect 9740 293728 9845 293734
rect 9680 293710 9740 293720
rect 9905 293728 10045 293734
rect 9845 293710 9905 293720
rect 10105 293728 10235 293734
rect 10045 293710 10105 293720
rect 10295 293728 10415 293734
rect 10235 293710 10295 293720
rect 10475 293728 10615 293734
rect 10415 293710 10475 293720
rect 10675 293728 10805 293734
rect 10615 293710 10675 293720
rect 10865 293728 10965 293734
rect 10805 293710 10865 293720
rect 11025 293728 11155 293734
rect 10965 293710 11025 293720
rect 11215 293728 11330 293734
rect 11155 293710 11215 293720
rect 11390 293728 11470 293734
rect 11330 293710 11390 293720
rect 11530 293728 15990 293734
rect 16020 293771 16068 293783
rect 11470 293710 11530 293720
rect 5700 293680 5960 293685
rect 16020 293680 16060 293771
rect 5700 293676 6000 293680
rect 15970 293676 16060 293680
rect 5700 293670 16060 293676
rect 5700 293636 6002 293670
rect 15978 293636 16060 293670
rect 5700 293633 16060 293636
rect 16120 293750 16170 294040
rect 536279 294086 537089 294114
rect 537169 294086 537239 294142
rect 537319 294114 537415 294142
rect 537557 294172 537563 294182
rect 538645 294182 538691 294194
rect 538753 294182 538799 294194
rect 539881 294182 539927 294194
rect 539989 294182 540035 294194
rect 538645 294172 538651 294182
rect 537557 294114 538651 294172
rect 538793 294172 538799 294182
rect 539879 294172 539887 294182
rect 538793 294142 539887 294172
rect 538793 294114 539579 294142
rect 537319 294112 537419 294114
rect 537549 294112 538659 294114
rect 538789 294112 539579 294114
rect 537319 294086 539579 294112
rect 539659 294086 539729 294142
rect 539809 294114 539887 294142
rect 540029 294172 540035 294182
rect 541117 294182 541163 294194
rect 541225 294182 541271 294194
rect 541117 294172 541123 294182
rect 540029 294114 541123 294172
rect 541265 294172 541271 294182
rect 542353 294182 542399 294194
rect 542461 294182 542507 294194
rect 543589 294182 543635 294194
rect 543697 294182 543743 294194
rect 542353 294172 542359 294182
rect 541265 294142 542359 294172
rect 541265 294114 542059 294142
rect 539809 294112 539889 294114
rect 540019 294112 541129 294114
rect 541259 294112 542059 294114
rect 539809 294086 542059 294112
rect 542139 294086 542209 294142
rect 542289 294114 542359 294142
rect 542501 294172 542509 294182
rect 543589 294172 543595 294182
rect 542501 294114 543595 294172
rect 543737 294172 543743 294182
rect 544825 294182 544871 294194
rect 544825 294172 544831 294182
rect 543737 294114 544831 294172
rect 544865 294114 544871 294182
rect 542289 294112 542369 294114
rect 542499 294112 543599 294114
rect 543729 294112 544871 294114
rect 542289 294102 544871 294112
rect 542289 294086 544859 294102
rect 536279 294052 536380 294086
rect 537356 294052 537616 294086
rect 538592 294052 538852 294086
rect 539828 294052 540088 294086
rect 541064 294052 541324 294086
rect 542300 294052 542560 294086
rect 543536 294052 543796 294086
rect 544772 294052 544859 294086
rect 536279 294032 536699 294052
rect 536689 293992 536699 294032
rect 536779 294032 536869 294052
rect 536779 293992 536789 294032
rect 536859 293992 536869 294032
rect 536949 294032 539219 294052
rect 536949 293992 536959 294032
rect 539209 293992 539219 294032
rect 539299 294032 539389 294052
rect 539299 293992 539309 294032
rect 539379 293992 539389 294032
rect 539469 294032 541709 294052
rect 539469 293992 539479 294032
rect 541699 293992 541709 294032
rect 541789 294032 541879 294052
rect 541789 293992 541799 294032
rect 541869 293992 541879 294032
rect 541959 294032 544159 294052
rect 541959 293992 541969 294032
rect 544149 293982 544159 294032
rect 544239 294032 544329 294052
rect 544239 293982 544249 294032
rect 544319 293982 544329 294032
rect 544409 294032 544859 294052
rect 562260 294100 562300 294300
rect 562500 294100 562700 294300
rect 562900 294100 563100 294300
rect 563300 294100 563500 294300
rect 563700 294100 563900 294300
rect 564100 294100 564300 294300
rect 564500 294100 564700 294300
rect 564900 294100 565100 294300
rect 565300 294100 565500 294300
rect 565700 294100 565900 294300
rect 566100 294100 566300 294300
rect 566500 294100 566700 294300
rect 566900 294100 567100 294300
rect 567300 294100 567500 294300
rect 567700 294100 567840 294300
rect 544409 293982 544419 294032
rect 537969 293918 538229 293952
rect 540607 293922 540721 293928
rect 537967 293912 538229 293918
rect 537967 293842 537979 293912
rect 538069 293842 538119 293912
rect 538209 293842 538229 293912
rect 537967 293836 538229 293842
rect 540447 293912 540561 293918
rect 540447 293842 540459 293912
rect 540549 293842 540561 293912
rect 540607 293852 540619 293922
rect 540709 293852 540721 293922
rect 540607 293846 540721 293852
rect 542907 293922 543011 293928
rect 542907 293852 542919 293922
rect 542999 293852 543011 293922
rect 542907 293846 543011 293852
rect 543077 293922 543181 293928
rect 543077 293852 543089 293922
rect 543169 293852 543181 293922
rect 543077 293846 543181 293852
rect 562260 293900 567840 294100
rect 540447 293836 540561 293842
rect 537969 293802 538229 293836
rect 5700 293630 16068 293633
rect 5700 293580 5960 293630
rect 15970 293621 16068 293630
rect 15970 293620 16028 293621
rect 5700 293400 5740 293580
rect 5920 293523 5960 293580
rect 9680 293580 9740 293590
rect 5990 293572 9680 293578
rect 9845 293580 9905 293590
rect 9740 293572 9845 293578
rect 10045 293580 10105 293590
rect 9905 293572 10045 293578
rect 10235 293580 10295 293590
rect 10105 293572 10235 293578
rect 10415 293580 10475 293590
rect 10295 293572 10415 293578
rect 10615 293580 10675 293590
rect 10475 293572 10615 293578
rect 10805 293580 10865 293590
rect 10675 293572 10805 293578
rect 10965 293580 11025 293590
rect 10865 293572 10965 293578
rect 11155 293580 11215 293590
rect 11025 293572 11155 293578
rect 11330 293580 11390 293590
rect 11215 293572 11330 293578
rect 11470 293580 11530 293590
rect 11390 293572 11470 293578
rect 16020 293587 16028 293620
rect 16062 293587 16068 293621
rect 11530 293572 15990 293578
rect 5990 293538 6002 293572
rect 15978 293538 15990 293572
rect 5990 293532 9680 293538
rect 5952 293489 5960 293523
rect 9740 293532 9845 293538
rect 9680 293510 9740 293520
rect 9905 293532 10045 293538
rect 9845 293510 9905 293520
rect 10105 293532 10235 293538
rect 10045 293510 10105 293520
rect 10295 293532 10415 293538
rect 10235 293510 10295 293520
rect 10475 293532 10615 293538
rect 10415 293510 10475 293520
rect 10675 293532 10805 293538
rect 10615 293510 10675 293520
rect 10865 293532 10965 293538
rect 10805 293510 10865 293520
rect 11025 293532 11155 293538
rect 10965 293510 11025 293520
rect 11215 293532 11330 293538
rect 11155 293510 11215 293520
rect 11390 293532 11470 293538
rect 11330 293510 11390 293520
rect 11530 293532 15990 293538
rect 16020 293575 16068 293587
rect 11470 293510 11530 293520
rect 16020 293490 16060 293575
rect 5920 293480 5960 293489
rect 15970 293480 16060 293490
rect 5920 293474 16060 293480
rect 5920 293440 6002 293474
rect 15978 293440 16060 293474
rect 5920 293437 16060 293440
rect 5920 293434 16068 293437
rect 5920 293430 6000 293434
rect 15970 293430 16068 293434
rect 5920 293400 5960 293430
rect 16020 293425 16068 293430
rect 5700 293327 5960 293400
rect 9680 293390 9740 293400
rect 5990 293376 9680 293382
rect 9845 293390 9905 293400
rect 9740 293376 9845 293382
rect 10045 293390 10105 293400
rect 9905 293376 10045 293382
rect 10235 293390 10295 293400
rect 10105 293376 10235 293382
rect 10415 293390 10475 293400
rect 10295 293376 10415 293382
rect 10615 293390 10675 293400
rect 10475 293376 10615 293382
rect 10805 293390 10865 293400
rect 10675 293376 10805 293382
rect 10965 293390 11025 293400
rect 10865 293376 10965 293382
rect 11155 293390 11215 293400
rect 11025 293376 11155 293382
rect 11330 293390 11390 293400
rect 11215 293376 11330 293382
rect 11470 293390 11530 293400
rect 11390 293376 11470 293382
rect 16020 293391 16028 293425
rect 16062 293391 16068 293425
rect 11530 293376 15990 293382
rect 5990 293342 6002 293376
rect 15978 293342 15990 293376
rect 5990 293336 9680 293342
rect 5700 293293 5918 293327
rect 5952 293293 5960 293327
rect 9740 293336 9845 293342
rect 9680 293320 9740 293330
rect 9905 293336 10045 293342
rect 9845 293320 9905 293330
rect 10105 293336 10235 293342
rect 10045 293320 10105 293330
rect 10295 293336 10415 293342
rect 10235 293320 10295 293330
rect 10475 293336 10615 293342
rect 10415 293320 10475 293330
rect 10675 293336 10805 293342
rect 10615 293320 10675 293330
rect 10865 293336 10965 293342
rect 10805 293320 10865 293330
rect 11025 293336 11155 293342
rect 10965 293320 11025 293330
rect 11215 293336 11330 293342
rect 11155 293320 11215 293330
rect 11390 293336 11470 293342
rect 11330 293320 11390 293330
rect 11530 293336 15990 293342
rect 16020 293379 16068 293391
rect 11470 293320 11530 293330
rect 5700 293290 5960 293293
rect 16020 293290 16060 293379
rect 5700 293284 6000 293290
rect 15970 293284 16060 293290
rect 5700 293278 16060 293284
rect 5700 293244 6002 293278
rect 15978 293244 16060 293278
rect 5700 293241 16060 293244
rect 5700 293240 16068 293241
rect 5700 293060 5740 293240
rect 5920 293131 5960 293240
rect 5990 293238 16068 293240
rect 15970 293230 16068 293238
rect 16020 293229 16068 293230
rect 9680 293190 9740 293200
rect 5990 293180 9680 293186
rect 9845 293190 9905 293200
rect 9740 293180 9845 293186
rect 10045 293190 10105 293200
rect 9905 293180 10045 293186
rect 10235 293190 10295 293200
rect 10105 293180 10235 293186
rect 10415 293190 10475 293200
rect 10295 293180 10415 293186
rect 10615 293190 10675 293200
rect 10475 293180 10615 293186
rect 10805 293190 10865 293200
rect 10675 293180 10805 293186
rect 10965 293190 11025 293200
rect 10865 293180 10965 293186
rect 11155 293190 11215 293200
rect 11025 293180 11155 293186
rect 11330 293190 11390 293200
rect 11215 293180 11330 293186
rect 11470 293190 11530 293200
rect 11390 293180 11470 293186
rect 16020 293195 16028 293229
rect 16062 293195 16068 293229
rect 11530 293180 15990 293186
rect 5990 293146 6002 293180
rect 15978 293146 15990 293180
rect 5990 293140 9680 293146
rect 5952 293097 5960 293131
rect 9740 293140 9845 293146
rect 9680 293120 9740 293130
rect 9905 293140 10045 293146
rect 9845 293120 9905 293130
rect 10105 293140 10235 293146
rect 10045 293120 10105 293130
rect 10295 293140 10415 293146
rect 10235 293120 10295 293130
rect 10475 293140 10615 293146
rect 10415 293120 10475 293130
rect 10675 293140 10805 293146
rect 10615 293120 10675 293130
rect 10865 293140 10965 293146
rect 10805 293120 10865 293130
rect 11025 293140 11155 293146
rect 10965 293120 11025 293130
rect 11215 293140 11330 293146
rect 11155 293120 11215 293130
rect 11390 293140 11470 293146
rect 11330 293120 11390 293130
rect 11530 293140 15990 293146
rect 16020 293183 16068 293195
rect 11470 293120 11530 293130
rect 5920 293090 5960 293097
rect 16020 293090 16060 293183
rect 5920 293088 6000 293090
rect 15970 293088 16060 293090
rect 5920 293082 16060 293088
rect 5920 293060 6002 293082
rect 5700 293048 6002 293060
rect 15978 293048 16060 293082
rect 5700 293045 16060 293048
rect 16120 293164 16130 293750
rect 16164 293164 16170 293750
rect 537959 293722 537969 293772
rect 536359 293704 537969 293722
rect 538049 293722 538059 293772
rect 538129 293722 538139 293772
rect 538049 293704 538139 293722
rect 538219 293722 538229 293772
rect 540449 293722 540459 293782
rect 538219 293704 540459 293722
rect 540539 293722 540549 293782
rect 540619 293722 540629 293782
rect 540539 293704 540629 293722
rect 540709 293722 540719 293782
rect 542909 293722 542919 293762
rect 540709 293704 542919 293722
rect 542999 293722 543009 293762
rect 543079 293722 543089 293762
rect 542999 293704 543089 293722
rect 543169 293722 543179 293762
rect 543169 293704 544799 293722
rect 536359 293682 536380 293704
rect 536368 293670 536380 293682
rect 537356 293682 537616 293704
rect 537356 293670 537368 293682
rect 536368 293664 537368 293670
rect 537604 293670 537616 293682
rect 538592 293682 538852 293704
rect 538592 293670 538604 293682
rect 537604 293664 538604 293670
rect 538840 293670 538852 293682
rect 539828 293682 540088 293704
rect 539828 293670 539840 293682
rect 538840 293664 539840 293670
rect 540076 293670 540088 293682
rect 541064 293682 541324 293704
rect 541064 293670 541076 293682
rect 540076 293664 541076 293670
rect 541312 293670 541324 293682
rect 542300 293682 542560 293704
rect 543536 293682 543796 293704
rect 542300 293670 542312 293682
rect 541312 293664 542312 293670
rect 542548 293670 542560 293682
rect 543536 293670 543548 293682
rect 542548 293664 543548 293670
rect 543784 293670 543796 293682
rect 544772 293682 544799 293704
rect 562260 293700 562300 293900
rect 562500 293700 562700 293900
rect 562900 293700 563100 293900
rect 563300 293700 563500 293900
rect 563700 293700 563900 293900
rect 564100 293700 564300 293900
rect 564500 293700 564700 293900
rect 564900 293700 565100 293900
rect 565300 293700 565500 293900
rect 565700 293700 565900 293900
rect 566100 293700 566300 293900
rect 566500 293700 566700 293900
rect 566900 293700 567100 293900
rect 567300 293700 567500 293900
rect 567700 293700 567840 293900
rect 544772 293670 544784 293682
rect 543784 293664 544784 293670
rect 536281 293642 536327 293654
rect 536281 293574 536287 293642
rect 536321 293632 536327 293642
rect 537409 293642 537455 293654
rect 537517 293642 537563 293654
rect 537409 293632 537415 293642
rect 536321 293602 537415 293632
rect 536321 293574 537089 293602
rect 536281 293562 537089 293574
rect 536289 293546 537089 293562
rect 537169 293546 537239 293602
rect 537319 293574 537415 293602
rect 537557 293632 537563 293642
rect 538645 293642 538691 293654
rect 538753 293642 538799 293654
rect 539881 293642 539927 293654
rect 539989 293642 540035 293654
rect 538645 293632 538651 293642
rect 537557 293574 538651 293632
rect 538793 293632 538799 293642
rect 539879 293632 539887 293642
rect 538793 293602 539887 293632
rect 538793 293574 539579 293602
rect 537319 293572 537419 293574
rect 537549 293572 538659 293574
rect 538789 293572 539579 293574
rect 537319 293546 539579 293572
rect 539659 293546 539729 293602
rect 539809 293574 539887 293602
rect 540029 293632 540035 293642
rect 541117 293642 541163 293654
rect 541225 293642 541271 293654
rect 541117 293632 541123 293642
rect 540029 293574 541123 293632
rect 541265 293632 541271 293642
rect 542353 293642 542399 293654
rect 542461 293642 542507 293654
rect 543589 293642 543635 293654
rect 543697 293642 543743 293654
rect 542353 293632 542359 293642
rect 541265 293602 542359 293632
rect 541265 293574 542069 293602
rect 539809 293572 539889 293574
rect 540019 293572 541129 293574
rect 541259 293572 542069 293574
rect 539809 293546 542069 293572
rect 542149 293546 542209 293602
rect 542289 293574 542359 293602
rect 542501 293632 542509 293642
rect 543589 293632 543595 293642
rect 542501 293574 543595 293632
rect 543737 293632 543743 293642
rect 544825 293642 544871 293654
rect 544825 293632 544831 293642
rect 543737 293574 544831 293632
rect 544865 293574 544871 293642
rect 542289 293572 542369 293574
rect 542499 293572 543599 293574
rect 543729 293572 544871 293574
rect 542289 293562 544871 293572
rect 542289 293546 544869 293562
rect 536289 293512 536380 293546
rect 537356 293512 537616 293546
rect 538592 293512 538852 293546
rect 539828 293512 540088 293546
rect 541064 293512 541324 293546
rect 542300 293512 542560 293546
rect 543536 293512 543796 293546
rect 544772 293512 544869 293546
rect 536289 293492 536699 293512
rect 536689 293452 536699 293492
rect 536779 293492 536869 293512
rect 536779 293452 536789 293492
rect 536859 293452 536869 293492
rect 536949 293492 539219 293512
rect 536949 293452 536959 293492
rect 539209 293452 539219 293492
rect 539299 293492 539389 293512
rect 539299 293452 539309 293492
rect 539379 293452 539389 293492
rect 539469 293492 541709 293512
rect 539469 293452 539479 293492
rect 541699 293442 541709 293492
rect 541789 293492 541879 293512
rect 541789 293442 541799 293492
rect 541869 293442 541879 293492
rect 541959 293492 544159 293512
rect 541959 293442 541969 293492
rect 544149 293452 544159 293492
rect 544239 293492 544329 293512
rect 544239 293452 544249 293492
rect 544319 293452 544329 293492
rect 544409 293492 544869 293512
rect 562260 293520 567840 293700
rect 562260 293500 567820 293520
rect 544409 293452 544419 293492
rect 537967 293382 538071 293388
rect 537967 293302 537979 293382
rect 538059 293302 538071 293382
rect 537967 293296 538071 293302
rect 538137 293382 538241 293388
rect 538137 293302 538149 293382
rect 538229 293302 538241 293382
rect 538137 293296 538241 293302
rect 540447 293382 540551 293388
rect 540447 293302 540459 293382
rect 540539 293302 540551 293382
rect 540447 293296 540551 293302
rect 540617 293382 540721 293388
rect 540617 293302 540629 293382
rect 540709 293302 540721 293382
rect 540617 293296 540721 293302
rect 542907 293382 543011 293388
rect 542907 293302 542919 293382
rect 542999 293302 543011 293382
rect 542907 293296 543011 293302
rect 543077 293382 543181 293388
rect 543077 293302 543089 293382
rect 543169 293302 543181 293382
rect 543077 293296 543181 293302
rect 562260 293300 562300 293500
rect 562500 293300 562700 293500
rect 562900 293300 563100 293500
rect 563300 293300 563500 293500
rect 563700 293300 563900 293500
rect 564100 293300 564300 293500
rect 564500 293300 564700 293500
rect 564900 293300 565100 293500
rect 565300 293300 565500 293500
rect 565700 293300 565900 293500
rect 566100 293300 566300 293500
rect 566500 293300 566700 293500
rect 566900 293300 567100 293500
rect 567300 293300 567500 293500
rect 567700 293300 567820 293500
rect 537969 293192 537979 293252
rect 536369 293172 537979 293192
rect 538059 293192 538069 293252
rect 538139 293192 538149 293252
rect 538059 293172 538149 293192
rect 538229 293192 538239 293252
rect 540449 293192 540459 293262
rect 538229 293182 540459 293192
rect 540539 293192 540549 293262
rect 540619 293192 540629 293262
rect 540539 293182 540629 293192
rect 540709 293192 540719 293262
rect 542909 293192 542919 293252
rect 540709 293182 542919 293192
rect 538229 293172 542919 293182
rect 542999 293192 543009 293252
rect 543079 293192 543089 293252
rect 542999 293172 543089 293192
rect 543169 293192 543179 293252
rect 543169 293172 544809 293192
rect 536369 293170 544809 293172
rect 5700 293042 16068 293045
rect 5700 293040 6000 293042
rect 15970 293040 16068 293042
rect 16020 293033 16068 293040
rect 9680 293000 9740 293010
rect 5990 292984 9680 292990
rect 9845 292990 9905 293000
rect 10045 292990 10105 293000
rect 10235 292990 10295 293000
rect 10415 292990 10475 293000
rect 10615 292990 10675 293000
rect 10805 292990 10865 293000
rect 10965 292990 11025 293000
rect 11155 292990 11215 293000
rect 11330 292990 11390 293000
rect 11470 292990 11530 293000
rect 16020 292999 16028 293033
rect 16062 292999 16068 293033
rect 9740 292984 9845 292990
rect 9905 292984 10045 292990
rect 10105 292984 10235 292990
rect 10295 292984 10415 292990
rect 10475 292984 10615 292990
rect 10675 292984 10805 292990
rect 10865 292984 10965 292990
rect 11025 292984 11155 292990
rect 11215 292984 11330 292990
rect 11390 292984 11470 292990
rect 11530 292984 15990 292990
rect 5990 292950 6002 292984
rect 15978 292950 15990 292984
rect 16020 292987 16068 292999
rect 16020 292980 16060 292987
rect 5990 292944 9680 292950
rect 9740 292944 9845 292950
rect 9680 292930 9740 292940
rect 9905 292944 10045 292950
rect 9845 292920 9905 292930
rect 10105 292944 10235 292950
rect 10045 292920 10105 292930
rect 10295 292944 10415 292950
rect 10235 292920 10295 292930
rect 10475 292944 10615 292950
rect 10415 292920 10475 292930
rect 10675 292944 10805 292950
rect 10615 292920 10675 292930
rect 10865 292944 10965 292950
rect 10805 292920 10865 292930
rect 11025 292944 11155 292950
rect 10965 292920 11025 292930
rect 11215 292944 11330 292950
rect 11155 292920 11215 292930
rect 11390 292944 11470 292950
rect 11330 292920 11390 292930
rect 11530 292944 15990 292950
rect 11470 292920 11530 292930
rect 16120 292880 16170 293164
rect 536368 293164 544809 293170
rect 536368 293130 536380 293164
rect 537356 293152 537616 293164
rect 537356 293130 537368 293152
rect 536368 293124 537368 293130
rect 537604 293130 537616 293152
rect 538592 293152 538852 293164
rect 538592 293130 538604 293152
rect 537604 293124 538604 293130
rect 538840 293130 538852 293152
rect 539828 293152 540088 293164
rect 539828 293130 539840 293152
rect 538840 293124 539840 293130
rect 540076 293130 540088 293152
rect 541064 293152 541324 293164
rect 541064 293130 541076 293152
rect 540076 293124 541076 293130
rect 541312 293130 541324 293152
rect 542300 293152 542560 293164
rect 542300 293130 542312 293152
rect 541312 293124 542312 293130
rect 542548 293130 542560 293152
rect 543536 293152 543796 293164
rect 543536 293130 543548 293152
rect 542548 293124 543548 293130
rect 543784 293130 543796 293152
rect 544772 293152 544809 293164
rect 544772 293130 544784 293152
rect 543784 293124 544784 293130
rect 536281 293102 536327 293114
rect 536281 293034 536287 293102
rect 536321 293092 536327 293102
rect 537409 293102 537455 293114
rect 537517 293102 537563 293114
rect 537409 293092 537415 293102
rect 536321 293042 537415 293092
rect 536321 293034 536327 293042
rect 536281 293022 536327 293034
rect 537409 293034 537415 293042
rect 537557 293092 537563 293102
rect 538645 293102 538691 293114
rect 538753 293102 538799 293114
rect 539881 293102 539927 293114
rect 539989 293102 540035 293114
rect 538645 293092 538651 293102
rect 537557 293042 538651 293092
rect 537557 293034 537563 293042
rect 537409 293032 537419 293034
rect 537549 293032 537563 293034
rect 537409 293022 537455 293032
rect 537517 293022 537563 293032
rect 538645 293034 538651 293042
rect 538793 293092 538799 293102
rect 539879 293092 539887 293102
rect 538793 293042 539887 293092
rect 538793 293034 538799 293042
rect 538645 293032 538659 293034
rect 538789 293032 538799 293034
rect 539879 293034 539887 293042
rect 540029 293092 540035 293102
rect 541117 293102 541163 293114
rect 541225 293102 541271 293114
rect 542353 293102 542399 293114
rect 542461 293102 542507 293114
rect 541117 293092 541123 293102
rect 540029 293042 541123 293092
rect 540029 293034 540035 293042
rect 539879 293032 539889 293034
rect 540019 293032 540035 293034
rect 538645 293022 538691 293032
rect 538753 293022 538799 293032
rect 539881 293022 539927 293032
rect 539989 293022 540035 293032
rect 541117 293034 541123 293042
rect 541265 293092 541271 293102
rect 542349 293092 542359 293102
rect 541265 293042 542359 293092
rect 541265 293034 541271 293042
rect 541117 293032 541129 293034
rect 541259 293032 541271 293034
rect 542349 293032 542359 293042
rect 542501 293092 542507 293102
rect 543589 293102 543635 293114
rect 543697 293102 543743 293114
rect 543589 293092 543595 293102
rect 542501 293042 543595 293092
rect 542501 293034 542507 293042
rect 542489 293032 542507 293034
rect 541117 293022 541163 293032
rect 541225 293022 541271 293032
rect 542353 293022 542399 293032
rect 542461 293022 542507 293032
rect 543589 293034 543595 293042
rect 543737 293092 543743 293102
rect 544825 293102 544871 293114
rect 544825 293092 544831 293102
rect 543737 293042 544831 293092
rect 543737 293034 543743 293042
rect 543589 293032 543599 293034
rect 543729 293032 543743 293034
rect 543589 293022 543635 293032
rect 543697 293022 543743 293032
rect 544825 293034 544831 293042
rect 544865 293034 544871 293102
rect 544825 293022 544871 293034
rect 536368 293006 537368 293012
rect 536368 292992 536380 293006
rect 537356 292992 537368 293006
rect 537604 293006 538604 293012
rect 537604 292992 537616 293006
rect 536359 292972 536380 292992
rect 537356 292972 537616 292992
rect 538592 292992 538604 293006
rect 538840 293006 539840 293012
rect 538840 292992 538852 293006
rect 539828 292992 539840 293006
rect 540076 293006 541076 293012
rect 540076 292992 540088 293006
rect 538592 292972 538852 292992
rect 539828 292972 540088 292992
rect 541064 292992 541076 293006
rect 541312 293006 542312 293012
rect 541312 292992 541324 293006
rect 542300 292992 542312 293006
rect 542548 293006 543548 293012
rect 542548 292992 542560 293006
rect 543536 292992 543548 293006
rect 543784 293006 544784 293012
rect 543784 292992 543796 293006
rect 544772 292992 544784 293006
rect 541064 292972 541324 292992
rect 542300 292972 542560 292992
rect 543536 292972 543796 292992
rect 544772 292972 544799 292992
rect 536359 292952 536699 292972
rect 536689 292912 536699 292952
rect 536779 292952 536869 292972
rect 536779 292912 536789 292952
rect 536859 292912 536869 292952
rect 536949 292952 538379 292972
rect 536949 292912 536959 292952
rect 538359 292922 538379 292952
rect 538459 292922 538489 292972
rect 538569 292952 539209 292972
rect 538569 292922 538589 292952
rect 538359 292892 538589 292922
rect 539199 292912 539209 292952
rect 539289 292952 539379 292972
rect 539289 292912 539299 292952
rect 539369 292912 539379 292952
rect 539459 292952 540789 292972
rect 539459 292912 539469 292952
rect 540769 292922 540789 292952
rect 540869 292922 540899 292972
rect 540979 292952 541699 292972
rect 540979 292922 540999 292952
rect 540769 292912 540999 292922
rect 541689 292912 541699 292952
rect 541779 292952 541869 292972
rect 541779 292912 541789 292952
rect 541859 292912 541869 292952
rect 541949 292952 543249 292972
rect 541949 292912 541959 292952
rect 543229 292912 543249 292952
rect 543329 292912 543359 292972
rect 543439 292952 544189 292972
rect 543439 292912 543459 292952
rect 544179 292912 544189 292952
rect 544269 292952 544359 292972
rect 544269 292912 544279 292952
rect 544349 292912 544359 292952
rect 544439 292952 544799 292972
rect 544439 292912 544449 292952
rect 543229 292892 543459 292912
rect 5900 292870 16170 292880
rect 5900 292836 8420 292870
rect 13560 292860 16170 292870
rect 13560 292836 15000 292860
rect 5900 292830 15000 292836
rect 14960 292720 15000 292830
rect 15140 292720 15200 292860
rect 15340 292830 16170 292860
rect 15340 292720 15380 292830
rect 14960 292680 15380 292720
rect 537969 292612 537979 292672
rect 536359 292592 537979 292612
rect 538059 292612 538069 292672
rect 538139 292612 538149 292672
rect 538059 292592 538149 292612
rect 538229 292612 538239 292672
rect 540449 292612 540459 292682
rect 538229 292602 540459 292612
rect 540539 292612 540549 292682
rect 540619 292612 540629 292682
rect 540539 292602 540629 292612
rect 540709 292612 540719 292682
rect 542909 292612 542919 292672
rect 540709 292602 542919 292612
rect 538229 292592 542919 292602
rect 542999 292612 543009 292672
rect 543079 292612 543089 292672
rect 542999 292592 543089 292612
rect 543169 292612 543179 292672
rect 543169 292592 544799 292612
rect 536359 292584 544799 292592
rect 536359 292572 536380 292584
rect 536368 292550 536380 292572
rect 537356 292572 537616 292584
rect 537356 292550 537368 292572
rect 536368 292544 537368 292550
rect 537604 292550 537616 292572
rect 538592 292572 538852 292584
rect 538592 292550 538604 292572
rect 537604 292544 538604 292550
rect 538840 292550 538852 292572
rect 539828 292572 540088 292584
rect 539828 292550 539840 292572
rect 538840 292544 539840 292550
rect 540076 292550 540088 292572
rect 541064 292572 541324 292584
rect 541064 292550 541076 292572
rect 540076 292544 541076 292550
rect 541312 292550 541324 292572
rect 542300 292572 542560 292584
rect 542300 292550 542312 292572
rect 541312 292544 542312 292550
rect 542548 292550 542560 292572
rect 543536 292572 543796 292584
rect 543536 292550 543548 292572
rect 542548 292544 543548 292550
rect 543784 292550 543796 292572
rect 544772 292572 544799 292584
rect 544772 292550 544784 292572
rect 543784 292544 544784 292550
rect 536281 292522 536327 292534
rect 536281 292454 536287 292522
rect 536321 292512 536327 292522
rect 537409 292522 537455 292534
rect 537517 292522 537563 292534
rect 537409 292512 537415 292522
rect 536321 292462 537415 292512
rect 536321 292454 536327 292462
rect 536281 292442 536327 292454
rect 537409 292454 537415 292462
rect 537557 292512 537563 292522
rect 538645 292522 538691 292534
rect 538753 292522 538799 292534
rect 538645 292512 538651 292522
rect 537557 292462 538651 292512
rect 537557 292454 537563 292462
rect 537409 292452 537419 292454
rect 537549 292452 537563 292454
rect 537409 292442 537455 292452
rect 537517 292442 537563 292452
rect 538645 292454 538651 292462
rect 538793 292512 538799 292522
rect 539881 292522 539927 292534
rect 539989 292522 540035 292534
rect 541117 292522 541163 292534
rect 541225 292522 541271 292534
rect 542353 292522 542399 292534
rect 542461 292522 542507 292534
rect 539881 292512 539887 292522
rect 538793 292462 539887 292512
rect 538793 292454 538799 292462
rect 538645 292452 538659 292454
rect 538789 292452 538799 292454
rect 538645 292442 538691 292452
rect 538753 292442 538799 292452
rect 539881 292454 539887 292462
rect 540029 292512 540039 292522
rect 541117 292512 541123 292522
rect 540029 292462 541123 292512
rect 539881 292452 539899 292454
rect 540029 292452 540039 292462
rect 541117 292454 541123 292462
rect 541265 292512 541271 292522
rect 542349 292512 542359 292522
rect 541265 292462 542359 292512
rect 541265 292454 541271 292462
rect 541117 292452 541129 292454
rect 541259 292452 541271 292454
rect 542349 292452 542359 292462
rect 542501 292512 542507 292522
rect 543589 292522 543635 292534
rect 543697 292522 543743 292534
rect 543589 292512 543595 292522
rect 542501 292462 543595 292512
rect 542501 292454 542507 292462
rect 542489 292452 542507 292454
rect 539881 292442 539927 292452
rect 539989 292442 540035 292452
rect 541117 292442 541163 292452
rect 541225 292442 541271 292452
rect 542353 292442 542399 292452
rect 542461 292442 542507 292452
rect 543589 292454 543595 292462
rect 543737 292512 543743 292522
rect 544825 292522 544871 292534
rect 544825 292512 544831 292522
rect 543737 292462 544831 292512
rect 543737 292454 543743 292462
rect 543589 292452 543599 292454
rect 543729 292452 543743 292454
rect 543589 292442 543635 292452
rect 543697 292442 543743 292452
rect 544825 292454 544831 292462
rect 544865 292454 544871 292522
rect 544825 292442 544871 292454
rect 536368 292426 537368 292432
rect 536368 292412 536380 292426
rect 537356 292412 537368 292426
rect 537604 292426 538604 292432
rect 537604 292412 537616 292426
rect 536359 292392 536380 292412
rect 537356 292392 537616 292412
rect 538592 292412 538604 292426
rect 538840 292426 539840 292432
rect 538840 292412 538852 292426
rect 539828 292412 539840 292426
rect 540076 292426 541076 292432
rect 540076 292412 540088 292426
rect 541064 292412 541076 292426
rect 541312 292426 542312 292432
rect 541312 292412 541324 292426
rect 538592 292392 538852 292412
rect 539828 292392 540088 292412
rect 541064 292392 541324 292412
rect 542300 292412 542312 292426
rect 542548 292426 543548 292432
rect 542548 292412 542560 292426
rect 543536 292412 543548 292426
rect 543784 292426 544784 292432
rect 543784 292412 543796 292426
rect 544772 292412 544784 292426
rect 542300 292392 542560 292412
rect 543536 292392 543796 292412
rect 544772 292392 544799 292412
rect 536359 292372 536699 292392
rect 536689 292332 536699 292372
rect 536779 292372 536869 292392
rect 536779 292332 536789 292372
rect 536859 292332 536869 292372
rect 536949 292372 538379 292392
rect 536949 292332 536959 292372
rect 538359 292312 538379 292372
rect 538459 292312 538489 292392
rect 538569 292372 539209 292392
rect 538569 292312 538589 292372
rect 539199 292332 539209 292372
rect 539289 292372 539379 292392
rect 539289 292332 539299 292372
rect 539369 292332 539379 292372
rect 539459 292372 540789 292392
rect 539459 292332 539469 292372
rect 540769 292332 540789 292372
rect 540869 292332 540899 292392
rect 540979 292372 541699 292392
rect 540979 292332 540999 292372
rect 540769 292312 540999 292332
rect 541689 292322 541699 292372
rect 541779 292372 541869 292392
rect 541779 292322 541789 292372
rect 541859 292322 541869 292372
rect 541949 292372 543249 292392
rect 541949 292322 541959 292372
rect 543229 292332 543249 292372
rect 543329 292332 543359 292392
rect 543439 292372 544189 292392
rect 543439 292332 543459 292372
rect 544179 292332 544189 292372
rect 544269 292372 544359 292392
rect 544269 292332 544279 292372
rect 544349 292332 544359 292372
rect 544439 292372 544799 292392
rect 544439 292332 544449 292372
rect 543229 292312 543459 292332
rect 538359 292302 538589 292312
rect 550109 292302 550539 292422
rect 530609 292132 531039 292252
rect 537967 292222 538081 292228
rect 537967 292142 537979 292222
rect 538069 292142 538081 292222
rect 537967 292136 538081 292142
rect 538127 292222 538241 292228
rect 538127 292142 538139 292222
rect 538229 292142 538241 292222
rect 538127 292136 538241 292142
rect 540447 292212 540551 292218
rect 540447 292142 540459 292212
rect 540539 292142 540551 292212
rect 540447 292136 540551 292142
rect 540617 292212 540721 292218
rect 540617 292142 540629 292212
rect 540709 292142 540721 292212
rect 540617 292136 540721 292142
rect 542907 292212 543011 292218
rect 542907 292142 542919 292212
rect 542999 292142 543011 292212
rect 542907 292136 543011 292142
rect 543077 292212 543181 292218
rect 543077 292142 543089 292212
rect 543169 292142 543181 292212
rect 543077 292136 543181 292142
rect 550109 292162 550129 292302
rect 550259 292162 550389 292302
rect 550519 292162 550539 292302
rect 530609 291992 530629 292132
rect 530759 291992 530879 292132
rect 531009 291992 531039 292132
rect 537969 292032 537979 292092
rect 536359 292012 537979 292032
rect 538059 292032 538069 292092
rect 538139 292032 538149 292092
rect 538059 292012 538149 292032
rect 538229 292032 538239 292092
rect 540449 292032 540459 292102
rect 538229 292022 540459 292032
rect 540539 292032 540549 292102
rect 540619 292032 540629 292102
rect 540539 292022 540629 292032
rect 540709 292032 540719 292102
rect 542909 292032 542919 292092
rect 540709 292022 542919 292032
rect 538229 292012 542919 292022
rect 542999 292032 543009 292092
rect 543079 292032 543089 292092
rect 542999 292012 543089 292032
rect 543169 292032 543179 292092
rect 543169 292012 544799 292032
rect 536359 292004 544799 292012
rect 536359 291992 536380 292004
rect 530609 291967 531039 291992
rect 536368 291970 536380 291992
rect 537356 291992 537616 292004
rect 537356 291970 537368 291992
rect 530609 291955 531143 291967
rect 530609 290841 530740 291955
rect 531137 290841 531143 291955
rect 533165 291955 533574 291967
rect 536368 291964 537368 291970
rect 537604 291970 537616 291992
rect 538592 291992 538852 292004
rect 538592 291970 538604 291992
rect 537604 291964 538604 291970
rect 538840 291970 538852 291992
rect 539828 291992 540088 292004
rect 539828 291970 539840 291992
rect 538840 291964 539840 291970
rect 540076 291970 540088 291992
rect 541064 291992 541324 292004
rect 541064 291970 541076 291992
rect 540076 291964 541076 291970
rect 541312 291970 541324 291992
rect 542300 291992 542560 292004
rect 542300 291970 542312 291992
rect 541312 291964 542312 291970
rect 542548 291970 542560 291992
rect 543536 291992 543796 292004
rect 543536 291970 543548 291992
rect 542548 291964 543548 291970
rect 543784 291970 543796 291992
rect 544772 291992 544799 292004
rect 544772 291970 544784 291992
rect 543784 291964 544784 291970
rect 550109 291967 550539 292162
rect 533165 291862 533171 291955
rect 530609 290829 531143 290841
rect 533039 290940 533171 291862
rect 533568 291422 533574 291955
rect 547794 291955 548203 291967
rect 536281 291942 536327 291954
rect 536281 291874 536287 291942
rect 536321 291932 536327 291942
rect 537409 291942 537455 291954
rect 537517 291942 537563 291954
rect 537409 291932 537415 291942
rect 536321 291882 537415 291932
rect 536321 291874 536327 291882
rect 536281 291862 536327 291874
rect 537409 291874 537415 291882
rect 537557 291932 537563 291942
rect 538645 291942 538691 291954
rect 538753 291942 538799 291954
rect 539881 291942 539927 291954
rect 539989 291942 540035 291954
rect 538645 291932 538651 291942
rect 537557 291882 538651 291932
rect 537557 291874 537563 291882
rect 537409 291872 537419 291874
rect 537549 291872 537563 291874
rect 537409 291862 537455 291872
rect 537517 291862 537563 291872
rect 538645 291874 538651 291882
rect 538793 291932 538799 291942
rect 539879 291932 539887 291942
rect 538793 291882 539887 291932
rect 538793 291874 538799 291882
rect 538645 291872 538659 291874
rect 538789 291872 538799 291874
rect 539879 291874 539887 291882
rect 540029 291932 540035 291942
rect 541117 291942 541163 291954
rect 541225 291942 541271 291954
rect 542353 291942 542399 291954
rect 542461 291942 542507 291954
rect 541117 291932 541123 291942
rect 540029 291882 541123 291932
rect 540029 291874 540035 291882
rect 539879 291872 539889 291874
rect 540019 291872 540035 291874
rect 538645 291862 538691 291872
rect 538753 291862 538799 291872
rect 539881 291862 539927 291872
rect 539989 291862 540035 291872
rect 541117 291874 541123 291882
rect 541265 291932 541271 291942
rect 542349 291932 542359 291942
rect 541265 291882 542359 291932
rect 541265 291874 541271 291882
rect 541117 291872 541129 291874
rect 541259 291872 541271 291874
rect 542349 291872 542359 291882
rect 542501 291932 542507 291942
rect 543589 291942 543635 291954
rect 543697 291942 543743 291954
rect 543589 291932 543595 291942
rect 542501 291882 543595 291932
rect 542501 291874 542507 291882
rect 542489 291872 542507 291874
rect 541117 291862 541163 291872
rect 541225 291862 541271 291872
rect 542353 291862 542399 291872
rect 542461 291862 542507 291872
rect 543589 291874 543595 291882
rect 543737 291932 543743 291942
rect 544825 291942 544871 291954
rect 544825 291932 544831 291942
rect 543737 291882 544831 291932
rect 543737 291874 543743 291882
rect 543589 291872 543599 291874
rect 543729 291872 543743 291874
rect 543589 291862 543635 291872
rect 543697 291862 543743 291872
rect 544825 291874 544831 291882
rect 544865 291874 544871 291942
rect 544825 291862 544871 291874
rect 547794 291862 547800 291955
rect 536368 291846 537368 291852
rect 536368 291822 536380 291846
rect 536359 291812 536380 291822
rect 537356 291822 537368 291846
rect 537604 291846 538604 291852
rect 537604 291822 537616 291846
rect 537356 291812 537616 291822
rect 538592 291822 538604 291846
rect 538840 291846 539840 291852
rect 538840 291822 538852 291846
rect 538592 291812 538852 291822
rect 539828 291822 539840 291846
rect 540076 291846 541076 291852
rect 540076 291822 540088 291846
rect 539828 291812 540088 291822
rect 541064 291822 541076 291846
rect 541312 291846 542312 291852
rect 541312 291822 541324 291846
rect 541064 291812 541324 291822
rect 542300 291822 542312 291846
rect 542548 291846 543548 291852
rect 542548 291822 542560 291846
rect 542300 291812 542560 291822
rect 543536 291822 543548 291846
rect 543784 291846 544784 291852
rect 543784 291822 543796 291846
rect 543536 291812 543796 291822
rect 544772 291822 544784 291846
rect 544772 291812 544799 291822
rect 536359 291802 539209 291812
rect 536359 291782 536679 291802
rect 536669 291722 536679 291782
rect 536759 291782 536889 291802
rect 536759 291722 536769 291782
rect 536879 291722 536889 291782
rect 536969 291782 539209 291802
rect 536969 291722 536979 291782
rect 538359 291732 538589 291782
rect 539199 291752 539209 291782
rect 539289 291782 539379 291812
rect 539289 291752 539299 291782
rect 539369 291752 539379 291782
rect 539459 291782 540789 291812
rect 539459 291752 539469 291782
rect 540769 291752 540789 291782
rect 540869 291752 540899 291812
rect 540979 291782 541699 291812
rect 540979 291752 540999 291782
rect 541689 291752 541699 291782
rect 541779 291782 541869 291812
rect 541779 291752 541789 291782
rect 541859 291752 541869 291782
rect 541949 291782 543249 291812
rect 541949 291752 541959 291782
rect 543229 291752 543249 291782
rect 543329 291752 543359 291812
rect 543439 291782 544189 291812
rect 543439 291752 543459 291782
rect 544179 291752 544189 291782
rect 544269 291782 544359 291812
rect 544269 291752 544279 291782
rect 544349 291752 544359 291782
rect 544439 291782 544799 291812
rect 544439 291752 544449 291782
rect 540769 291732 540999 291752
rect 543229 291732 543459 291752
rect 536089 291492 536099 291562
rect 534519 291482 536099 291492
rect 536179 291492 536189 291562
rect 536319 291492 536329 291562
rect 536179 291482 536329 291492
rect 536409 291492 536419 291562
rect 538639 291492 538649 291552
rect 536409 291482 538649 291492
rect 534519 291472 538649 291482
rect 538729 291492 538739 291552
rect 538809 291492 538819 291552
rect 538729 291472 538819 291492
rect 538899 291492 538909 291552
rect 541099 291492 541109 291552
rect 538899 291472 541109 291492
rect 541189 291492 541199 291552
rect 541289 291492 541299 291552
rect 541189 291472 541299 291492
rect 541379 291492 541389 291552
rect 543549 291492 543559 291552
rect 541379 291472 543559 291492
rect 543639 291492 543649 291552
rect 543739 291492 543749 291552
rect 543639 291472 543749 291492
rect 543829 291492 543839 291552
rect 546059 291492 546069 291552
rect 543829 291472 546069 291492
rect 546149 291492 546159 291552
rect 546229 291492 546239 291552
rect 546149 291472 546239 291492
rect 546319 291492 546329 291552
rect 546319 291472 546669 291492
rect 534519 291464 546669 291472
rect 534519 291442 534540 291464
rect 534528 291430 534540 291442
rect 535516 291442 535776 291464
rect 535516 291430 535528 291442
rect 534528 291424 535528 291430
rect 535764 291430 535776 291442
rect 536752 291442 537012 291464
rect 536752 291430 536764 291442
rect 535764 291424 536764 291430
rect 537000 291430 537012 291442
rect 537988 291442 538248 291464
rect 537988 291430 538000 291442
rect 537000 291424 538000 291430
rect 538236 291430 538248 291442
rect 539224 291442 539484 291464
rect 539224 291430 539236 291442
rect 538236 291424 539236 291430
rect 539472 291430 539484 291442
rect 540460 291442 540720 291464
rect 540460 291430 540472 291442
rect 539472 291424 540472 291430
rect 540708 291430 540720 291442
rect 541696 291442 541956 291464
rect 541696 291430 541708 291442
rect 540708 291424 541708 291430
rect 541944 291430 541956 291442
rect 542932 291442 543192 291464
rect 542932 291430 542944 291442
rect 541944 291424 542944 291430
rect 543180 291430 543192 291442
rect 544168 291442 544428 291464
rect 544168 291430 544180 291442
rect 543180 291424 544180 291430
rect 544416 291430 544428 291442
rect 545404 291442 545664 291464
rect 545404 291430 545416 291442
rect 544416 291424 545416 291430
rect 545652 291430 545664 291442
rect 546640 291442 546669 291464
rect 546640 291430 546652 291442
rect 545652 291424 546652 291430
rect 547669 291422 547800 291862
rect 533568 291414 534479 291422
rect 546699 291414 547800 291422
rect 533568 291402 534487 291414
rect 533568 291334 534447 291402
rect 534481 291392 534487 291402
rect 535569 291402 535615 291414
rect 535677 291402 535723 291414
rect 535569 291392 535575 291402
rect 534481 291352 535575 291392
rect 534481 291334 534487 291352
rect 533568 291322 534487 291334
rect 535569 291334 535575 291352
rect 535717 291392 535723 291402
rect 536805 291402 536851 291414
rect 536913 291402 536959 291414
rect 538041 291402 538087 291414
rect 538149 291402 538195 291414
rect 536805 291392 536811 291402
rect 535717 291352 536811 291392
rect 535717 291334 535723 291352
rect 535569 291332 535579 291334
rect 535709 291332 535723 291334
rect 535569 291322 535615 291332
rect 535677 291322 535723 291332
rect 536805 291334 536811 291352
rect 536953 291392 536959 291402
rect 538039 291392 538047 291402
rect 536953 291352 538047 291392
rect 536953 291334 536959 291352
rect 536805 291332 536819 291334
rect 536949 291332 536959 291334
rect 538039 291334 538047 291352
rect 538189 291392 538195 291402
rect 539277 291402 539323 291414
rect 539385 291402 539431 291414
rect 539277 291392 539283 291402
rect 538189 291352 539283 291392
rect 538189 291334 538195 291352
rect 538039 291332 538049 291334
rect 538179 291332 538195 291334
rect 536805 291322 536851 291332
rect 536913 291322 536959 291332
rect 538041 291322 538087 291332
rect 538149 291322 538195 291332
rect 539277 291334 539283 291352
rect 539425 291392 539431 291402
rect 540513 291402 540559 291414
rect 540621 291402 540667 291414
rect 541749 291402 541795 291414
rect 541857 291402 541903 291414
rect 540513 291392 540519 291402
rect 539425 291352 540519 291392
rect 539425 291334 539431 291352
rect 539277 291332 539289 291334
rect 539419 291332 539431 291334
rect 539277 291322 539323 291332
rect 539385 291322 539431 291332
rect 540513 291334 540519 291352
rect 540661 291392 540669 291402
rect 541749 291392 541755 291402
rect 540661 291352 541755 291392
rect 540661 291334 540669 291352
rect 540513 291332 540529 291334
rect 540659 291332 540669 291334
rect 541749 291334 541755 291352
rect 541897 291392 541903 291402
rect 542985 291402 543031 291414
rect 543093 291402 543139 291414
rect 544221 291402 544267 291414
rect 544329 291402 544375 291414
rect 542985 291392 542991 291402
rect 541897 291352 542991 291392
rect 541897 291334 541903 291352
rect 541749 291332 541759 291334
rect 541889 291332 541903 291334
rect 540513 291322 540559 291332
rect 540621 291322 540667 291332
rect 541749 291322 541795 291332
rect 541857 291322 541903 291332
rect 542985 291334 542991 291352
rect 543133 291392 543139 291402
rect 544219 291392 544227 291402
rect 543133 291352 544227 291392
rect 543133 291334 543139 291352
rect 542985 291332 542999 291334
rect 543129 291332 543139 291334
rect 544219 291334 544227 291352
rect 544369 291392 544375 291402
rect 545457 291402 545503 291414
rect 545565 291402 545611 291414
rect 545457 291392 545463 291402
rect 544369 291352 545463 291392
rect 544369 291334 544375 291352
rect 544219 291332 544229 291334
rect 544359 291332 544375 291334
rect 542985 291322 543031 291332
rect 543093 291322 543139 291332
rect 544221 291322 544267 291332
rect 544329 291322 544375 291332
rect 545457 291334 545463 291352
rect 545605 291392 545611 291402
rect 546693 291402 547800 291414
rect 546693 291392 546699 291402
rect 545605 291352 546699 291392
rect 545605 291334 545611 291352
rect 545457 291332 545469 291334
rect 545599 291332 545611 291334
rect 545457 291322 545503 291332
rect 545565 291322 545611 291332
rect 546693 291334 546699 291352
rect 546733 291334 547800 291402
rect 546693 291322 547800 291334
rect 533039 290880 533080 290940
rect 533140 290880 533171 290940
rect 533568 290882 533574 291322
rect 534528 291306 535528 291312
rect 534528 291292 534540 291306
rect 534519 291272 534540 291292
rect 535516 291292 535528 291306
rect 535764 291306 536764 291312
rect 535764 291292 535776 291306
rect 535516 291272 535776 291292
rect 536752 291292 536764 291306
rect 537000 291306 538000 291312
rect 537000 291292 537012 291306
rect 536752 291272 537012 291292
rect 537988 291292 538000 291306
rect 538236 291306 539236 291312
rect 538236 291292 538248 291306
rect 537988 291272 538248 291292
rect 539224 291292 539236 291306
rect 539472 291306 540472 291312
rect 539472 291292 539484 291306
rect 539224 291272 539484 291292
rect 540460 291292 540472 291306
rect 540708 291306 541708 291312
rect 540708 291292 540720 291306
rect 540460 291272 540720 291292
rect 541696 291292 541708 291306
rect 541944 291306 542944 291312
rect 541944 291292 541956 291306
rect 541696 291272 541956 291292
rect 542932 291292 542944 291306
rect 543180 291306 544180 291312
rect 543180 291292 543192 291306
rect 542932 291272 543192 291292
rect 544168 291292 544180 291306
rect 544416 291306 545416 291312
rect 544416 291292 544428 291306
rect 544168 291272 544428 291292
rect 545404 291292 545416 291306
rect 545652 291306 546652 291312
rect 545652 291292 545664 291306
rect 545404 291272 545664 291292
rect 546640 291292 546652 291306
rect 546640 291272 546669 291292
rect 534519 291242 534849 291272
rect 534839 291202 534849 291242
rect 534929 291242 535059 291272
rect 534929 291202 534939 291242
rect 535049 291202 535059 291242
rect 535139 291242 537329 291272
rect 535139 291202 535149 291242
rect 537319 291202 537329 291242
rect 537409 291242 537549 291272
rect 537409 291202 537419 291242
rect 537539 291202 537549 291242
rect 537629 291242 539859 291272
rect 537629 291202 537639 291242
rect 539849 291202 539859 291242
rect 539939 291242 540039 291272
rect 539939 291202 539949 291242
rect 540029 291202 540039 291242
rect 540119 291242 542319 291272
rect 540119 291202 540129 291242
rect 542309 291192 542319 291242
rect 542399 291242 542499 291272
rect 542399 291192 542409 291242
rect 542489 291192 542499 291242
rect 542579 291242 544799 291272
rect 542579 291192 542589 291242
rect 544789 291192 544799 291242
rect 544879 291242 544969 291272
rect 544879 291192 544889 291242
rect 544959 291192 544969 291242
rect 545049 291242 546669 291272
rect 545049 291192 545059 291242
rect 536107 291142 536221 291148
rect 536107 291062 536119 291142
rect 536209 291062 536221 291142
rect 536107 291056 536221 291062
rect 536287 291142 536401 291148
rect 536287 291062 536299 291142
rect 536389 291062 536401 291142
rect 536287 291056 536401 291062
rect 538637 291142 538751 291148
rect 538637 291062 538649 291142
rect 538739 291062 538751 291142
rect 538637 291056 538751 291062
rect 538797 291142 538911 291148
rect 538797 291062 538809 291142
rect 538899 291062 538911 291142
rect 538797 291056 538911 291062
rect 541107 291142 541221 291148
rect 541107 291062 541119 291142
rect 541209 291062 541221 291142
rect 541107 291056 541221 291062
rect 541267 291142 541381 291148
rect 541267 291062 541279 291142
rect 541369 291062 541381 291142
rect 541267 291056 541381 291062
rect 543557 291142 543671 291148
rect 543557 291062 543569 291142
rect 543659 291062 543671 291142
rect 543557 291056 543671 291062
rect 543717 291142 543831 291148
rect 543717 291062 543729 291142
rect 543819 291062 543831 291142
rect 543717 291056 543831 291062
rect 546057 291142 546171 291148
rect 546057 291062 546069 291142
rect 546159 291062 546171 291142
rect 546057 291056 546171 291062
rect 546217 291142 546331 291148
rect 546217 291062 546229 291142
rect 546319 291062 546331 291142
rect 546217 291056 546331 291062
rect 536089 290962 536099 291022
rect 534519 290942 536099 290962
rect 536179 290962 536189 291022
rect 536319 290962 536329 291022
rect 536179 290942 536329 290962
rect 536409 290962 536419 291022
rect 538639 290962 538649 291012
rect 536409 290942 538649 290962
rect 534519 290932 538649 290942
rect 538729 290962 538739 291012
rect 538809 290962 538819 291022
rect 538729 290942 538819 290962
rect 538899 290962 538909 291022
rect 541099 290962 541109 291022
rect 538899 290942 541109 290962
rect 541189 290962 541199 291022
rect 541289 290962 541299 291022
rect 541189 290942 541299 290962
rect 541379 290962 541389 291022
rect 543549 290962 543559 291012
rect 541379 290942 543559 290962
rect 538729 290932 543559 290942
rect 543639 290962 543649 291012
rect 543739 290962 543749 291012
rect 543639 290932 543749 290962
rect 543829 290962 543839 291012
rect 546059 290962 546069 291012
rect 543829 290932 546069 290962
rect 546149 290962 546159 291012
rect 546229 290962 546239 291012
rect 546149 290932 546239 290962
rect 546319 290962 546329 291012
rect 546319 290932 546669 290962
rect 534519 290924 546669 290932
rect 534519 290912 534540 290924
rect 534528 290890 534540 290912
rect 535516 290912 535776 290924
rect 535516 290890 535528 290912
rect 534528 290884 535528 290890
rect 535764 290890 535776 290912
rect 536752 290912 537012 290924
rect 536752 290890 536764 290912
rect 535764 290884 536764 290890
rect 537000 290890 537012 290912
rect 537988 290912 538248 290924
rect 537988 290890 538000 290912
rect 537000 290884 538000 290890
rect 538236 290890 538248 290912
rect 539224 290912 539484 290924
rect 539224 290890 539236 290912
rect 538236 290884 539236 290890
rect 539472 290890 539484 290912
rect 540460 290912 540720 290924
rect 540460 290890 540472 290912
rect 539472 290884 540472 290890
rect 540708 290890 540720 290912
rect 541696 290912 541956 290924
rect 541696 290890 541708 290912
rect 540708 290884 541708 290890
rect 541944 290890 541956 290912
rect 542932 290912 543192 290924
rect 542932 290890 542944 290912
rect 541944 290884 542944 290890
rect 543180 290890 543192 290912
rect 544168 290912 544428 290924
rect 544168 290890 544180 290912
rect 543180 290884 544180 290890
rect 544416 290890 544428 290912
rect 545404 290912 545664 290924
rect 545404 290890 545416 290912
rect 544416 290884 545416 290890
rect 545652 290890 545664 290912
rect 546640 290912 546669 290924
rect 546640 290890 546652 290912
rect 545652 290884 546652 290890
rect 533039 290841 533171 290880
rect 533568 290874 534479 290882
rect 533568 290862 534487 290874
rect 533568 290841 534447 290862
rect 530609 290497 531039 290829
rect 533039 290820 534447 290841
rect 533039 290760 533080 290820
rect 533140 290760 533180 290820
rect 533240 290760 533280 290820
rect 533340 290794 534447 290820
rect 534481 290852 534487 290862
rect 535569 290872 535615 290874
rect 535677 290872 535723 290874
rect 535569 290862 535579 290872
rect 535709 290862 535723 290872
rect 535569 290852 535575 290862
rect 534481 290812 535575 290852
rect 534481 290794 534487 290812
rect 533340 290782 534487 290794
rect 535569 290794 535575 290812
rect 535717 290852 535723 290862
rect 536805 290862 536851 290874
rect 536913 290862 536959 290874
rect 538041 290862 538087 290874
rect 538149 290862 538195 290874
rect 536805 290852 536811 290862
rect 535717 290812 536811 290852
rect 535609 290794 535615 290802
rect 535569 290782 535615 290794
rect 535677 290794 535683 290802
rect 535717 290794 535723 290812
rect 535677 290782 535723 290794
rect 536805 290794 536811 290812
rect 536953 290852 536959 290862
rect 538039 290852 538047 290862
rect 536953 290812 538047 290852
rect 536953 290794 536959 290812
rect 536805 290792 536819 290794
rect 536949 290792 536959 290794
rect 538039 290794 538047 290812
rect 538189 290852 538195 290862
rect 539277 290862 539323 290874
rect 539385 290862 539431 290874
rect 539277 290852 539283 290862
rect 538189 290812 539283 290852
rect 538189 290794 538195 290812
rect 538039 290792 538049 290794
rect 538179 290792 538195 290794
rect 536805 290782 536851 290792
rect 536913 290782 536959 290792
rect 538041 290782 538087 290792
rect 538149 290782 538195 290792
rect 539277 290794 539283 290812
rect 539425 290852 539431 290862
rect 540513 290862 540559 290874
rect 540621 290862 540667 290874
rect 541749 290862 541795 290874
rect 541857 290862 541903 290874
rect 540513 290852 540519 290862
rect 539425 290812 540519 290852
rect 539425 290794 539431 290812
rect 539277 290792 539289 290794
rect 539419 290792 539431 290794
rect 539277 290782 539323 290792
rect 539385 290782 539431 290792
rect 540513 290794 540519 290812
rect 540661 290852 540669 290862
rect 541749 290852 541755 290862
rect 540661 290812 541755 290852
rect 540661 290794 540669 290812
rect 540513 290792 540529 290794
rect 540659 290792 540669 290794
rect 541749 290794 541755 290812
rect 541897 290852 541903 290862
rect 542985 290862 543031 290874
rect 543093 290862 543139 290874
rect 544221 290862 544267 290874
rect 544329 290862 544375 290874
rect 542985 290852 542991 290862
rect 541897 290812 542991 290852
rect 541897 290794 541903 290812
rect 541749 290792 541759 290794
rect 541889 290792 541903 290794
rect 540513 290782 540559 290792
rect 540621 290782 540667 290792
rect 541749 290782 541795 290792
rect 541857 290782 541903 290792
rect 542985 290794 542991 290812
rect 543133 290852 543139 290862
rect 544219 290852 544227 290862
rect 543133 290812 544227 290852
rect 543133 290794 543139 290812
rect 542985 290792 542999 290794
rect 543129 290792 543139 290794
rect 544219 290794 544227 290812
rect 544369 290852 544375 290862
rect 545457 290862 545503 290874
rect 545565 290862 545611 290874
rect 545457 290852 545463 290862
rect 544369 290812 545463 290852
rect 544369 290794 544375 290812
rect 544219 290792 544229 290794
rect 544359 290792 544375 290794
rect 542985 290782 543031 290792
rect 543093 290782 543139 290792
rect 544221 290782 544267 290792
rect 544329 290782 544375 290792
rect 545457 290794 545463 290812
rect 545605 290852 545611 290862
rect 546693 290872 546739 290874
rect 547669 290872 547800 291322
rect 546693 290862 547800 290872
rect 546693 290852 546699 290862
rect 545605 290812 546699 290852
rect 545605 290794 545611 290812
rect 545457 290792 545469 290794
rect 545599 290792 545611 290794
rect 545457 290782 545503 290792
rect 545565 290782 545611 290792
rect 546693 290794 546699 290812
rect 546733 290841 547800 290862
rect 548197 290841 548203 291955
rect 546733 290829 548203 290841
rect 550109 291955 550634 291967
rect 550109 290841 550231 291955
rect 550628 290841 550634 291955
rect 550109 290829 550634 290841
rect 546733 290794 548099 290829
rect 546693 290782 548099 290794
rect 533340 290772 534479 290782
rect 546699 290772 548099 290782
rect 533340 290760 533469 290772
rect 533039 290720 533469 290760
rect 534528 290766 535528 290772
rect 534528 290752 534540 290766
rect 533039 290660 533080 290720
rect 533140 290660 533180 290720
rect 533240 290660 533280 290720
rect 533340 290660 533469 290720
rect 534519 290732 534540 290752
rect 535516 290752 535528 290766
rect 535764 290766 536764 290772
rect 535764 290752 535776 290766
rect 535516 290732 535776 290752
rect 536752 290752 536764 290766
rect 537000 290766 538000 290772
rect 537000 290752 537012 290766
rect 536752 290732 537012 290752
rect 537988 290752 538000 290766
rect 538236 290766 539236 290772
rect 538236 290752 538248 290766
rect 537988 290732 538248 290752
rect 539224 290752 539236 290766
rect 539472 290766 540472 290772
rect 539472 290752 539484 290766
rect 539224 290732 539484 290752
rect 540460 290752 540472 290766
rect 540708 290766 541708 290772
rect 540708 290752 540720 290766
rect 540460 290732 540720 290752
rect 541696 290752 541708 290766
rect 541944 290766 542944 290772
rect 541944 290752 541956 290766
rect 541696 290732 541956 290752
rect 542932 290752 542944 290766
rect 543180 290766 544180 290772
rect 543180 290752 543192 290766
rect 542932 290732 543192 290752
rect 544168 290752 544180 290766
rect 544416 290766 545416 290772
rect 544416 290752 544428 290766
rect 544168 290732 544428 290752
rect 545404 290752 545416 290766
rect 545652 290766 546652 290772
rect 545652 290752 545664 290766
rect 545404 290732 545664 290752
rect 546640 290752 546652 290766
rect 546640 290732 546669 290752
rect 534519 290702 534849 290732
rect 534839 290662 534849 290702
rect 534929 290702 535059 290732
rect 534929 290662 534939 290702
rect 535049 290662 535059 290702
rect 535139 290702 537329 290732
rect 535139 290662 535149 290702
rect 537319 290662 537329 290702
rect 537409 290702 537549 290732
rect 537409 290662 537419 290702
rect 537539 290662 537549 290702
rect 537629 290702 539859 290732
rect 537629 290662 537639 290702
rect 539849 290662 539859 290702
rect 539939 290702 540049 290732
rect 539939 290662 539949 290702
rect 540039 290662 540049 290702
rect 540129 290702 542319 290732
rect 540129 290662 540139 290702
rect 533039 290580 533469 290660
rect 542309 290652 542319 290702
rect 542399 290702 542499 290732
rect 542399 290652 542409 290702
rect 542489 290652 542499 290702
rect 542579 290702 544799 290732
rect 542579 290652 542589 290702
rect 544789 290652 544799 290702
rect 544879 290702 544969 290732
rect 544879 290652 544889 290702
rect 544959 290652 544969 290702
rect 545049 290702 546669 290732
rect 545049 290652 545059 290702
rect 533039 290520 533080 290580
rect 533140 290520 533180 290580
rect 533240 290520 533280 290580
rect 533340 290520 533469 290580
rect 533039 290497 533469 290520
rect 547669 290497 548099 290772
rect 550109 290497 550539 290829
rect 530609 290485 531143 290497
rect 530609 289392 530740 290485
rect 530734 289371 530740 289392
rect 531137 289371 531143 290485
rect 533039 290485 533574 290497
rect 533039 290480 533171 290485
rect 533039 290420 533080 290480
rect 533140 290420 533171 290480
rect 533039 290380 533171 290420
rect 533039 290320 533080 290380
rect 533140 290320 533171 290380
rect 533568 290342 533574 290485
rect 547669 290485 548203 290497
rect 536089 290422 536099 290482
rect 534519 290402 536099 290422
rect 536179 290422 536189 290482
rect 536319 290422 536329 290482
rect 536179 290402 536329 290422
rect 536409 290422 536419 290482
rect 538629 290422 538639 290472
rect 536409 290402 538639 290422
rect 534519 290392 538639 290402
rect 538719 290422 538729 290472
rect 538799 290422 538809 290472
rect 538719 290392 538809 290422
rect 538889 290422 538899 290472
rect 541099 290422 541109 290472
rect 538889 290392 541109 290422
rect 541189 290422 541199 290472
rect 541279 290422 541289 290472
rect 541189 290392 541289 290422
rect 541369 290422 541379 290472
rect 543549 290422 543559 290472
rect 541369 290392 543559 290422
rect 543639 290422 543649 290472
rect 543739 290422 543749 290472
rect 543639 290392 543749 290422
rect 543829 290422 543839 290472
rect 546059 290422 546069 290472
rect 543829 290392 546069 290422
rect 546149 290422 546159 290472
rect 546229 290422 546239 290472
rect 546149 290392 546239 290422
rect 546319 290422 546329 290472
rect 546319 290392 546669 290422
rect 534519 290384 546669 290392
rect 534519 290372 534540 290384
rect 534528 290350 534540 290372
rect 535516 290372 535776 290384
rect 535516 290350 535528 290372
rect 534528 290344 535528 290350
rect 535764 290350 535776 290372
rect 536752 290372 537012 290384
rect 536752 290350 536764 290372
rect 535764 290344 536764 290350
rect 537000 290350 537012 290372
rect 537988 290372 538248 290384
rect 537988 290350 538000 290372
rect 537000 290344 538000 290350
rect 538236 290350 538248 290372
rect 539224 290372 539484 290384
rect 539224 290350 539236 290372
rect 538236 290344 539236 290350
rect 539472 290350 539484 290372
rect 540460 290372 540720 290384
rect 540460 290350 540472 290372
rect 539472 290344 540472 290350
rect 540708 290350 540720 290372
rect 541696 290372 541956 290384
rect 541696 290350 541708 290372
rect 540708 290344 541708 290350
rect 541944 290350 541956 290372
rect 542932 290372 543192 290384
rect 542932 290350 542944 290372
rect 541944 290344 542944 290350
rect 543180 290350 543192 290372
rect 544168 290372 544428 290384
rect 544168 290350 544180 290372
rect 543180 290344 544180 290350
rect 544416 290350 544428 290372
rect 545404 290372 545664 290384
rect 545404 290350 545416 290372
rect 544416 290344 545416 290350
rect 545652 290350 545664 290372
rect 546640 290372 546669 290384
rect 546640 290350 546652 290372
rect 545652 290344 546652 290350
rect 547669 290342 547800 290485
rect 533568 290322 534499 290342
rect 546699 290334 547800 290342
rect 533039 290280 533171 290320
rect 533039 290220 533080 290280
rect 533140 290220 533171 290280
rect 533568 290254 534447 290322
rect 534481 290312 534499 290322
rect 535569 290322 535615 290334
rect 535677 290322 535723 290334
rect 535569 290312 535575 290322
rect 534481 290272 535575 290312
rect 534481 290254 534499 290272
rect 533568 290232 534499 290254
rect 535569 290254 535575 290272
rect 535717 290312 535723 290322
rect 536805 290322 536851 290334
rect 536913 290322 536959 290334
rect 538041 290322 538087 290334
rect 538149 290322 538195 290334
rect 536805 290312 536811 290322
rect 535717 290272 536811 290312
rect 535717 290254 535723 290272
rect 535569 290252 535579 290254
rect 535709 290252 535723 290254
rect 535569 290242 535615 290252
rect 535677 290242 535723 290252
rect 536805 290254 536811 290272
rect 536953 290312 536959 290322
rect 538039 290312 538047 290322
rect 536953 290272 538047 290312
rect 536953 290254 536959 290272
rect 536805 290252 536819 290254
rect 536949 290252 536959 290254
rect 538039 290254 538047 290272
rect 538189 290312 538195 290322
rect 539277 290322 539323 290334
rect 539385 290322 539431 290334
rect 539277 290312 539283 290322
rect 538189 290272 539283 290312
rect 538189 290254 538195 290272
rect 538039 290252 538049 290254
rect 538179 290252 538195 290254
rect 536805 290242 536851 290252
rect 536913 290242 536959 290252
rect 538041 290242 538087 290252
rect 538149 290242 538195 290252
rect 539277 290254 539283 290272
rect 539425 290312 539431 290322
rect 540513 290322 540559 290334
rect 540621 290322 540667 290334
rect 541749 290322 541795 290334
rect 541857 290322 541903 290334
rect 540513 290312 540519 290322
rect 539425 290272 540519 290312
rect 539425 290254 539431 290272
rect 539277 290252 539289 290254
rect 539419 290252 539431 290254
rect 539277 290242 539323 290252
rect 539385 290242 539431 290252
rect 540513 290254 540519 290272
rect 540661 290312 540669 290322
rect 541749 290312 541755 290322
rect 540661 290272 541755 290312
rect 540661 290254 540669 290272
rect 540513 290252 540529 290254
rect 540659 290252 540669 290254
rect 541749 290254 541755 290272
rect 541897 290312 541903 290322
rect 542985 290322 543031 290334
rect 543093 290322 543139 290334
rect 544221 290322 544267 290334
rect 544329 290322 544375 290334
rect 542985 290312 542991 290322
rect 541897 290272 542991 290312
rect 541897 290254 541903 290272
rect 541749 290252 541759 290254
rect 541889 290252 541903 290254
rect 540513 290242 540559 290252
rect 540621 290242 540667 290252
rect 541749 290242 541795 290252
rect 541857 290242 541903 290252
rect 542985 290254 542991 290272
rect 543133 290312 543139 290322
rect 544219 290312 544227 290322
rect 543133 290272 544227 290312
rect 543133 290254 543139 290272
rect 542985 290252 542999 290254
rect 543129 290252 543139 290254
rect 544219 290254 544227 290272
rect 544369 290312 544375 290322
rect 545457 290322 545503 290334
rect 545565 290322 545611 290334
rect 545457 290312 545463 290322
rect 544369 290272 545463 290312
rect 544369 290254 544375 290272
rect 544219 290252 544229 290254
rect 544359 290252 544375 290254
rect 542985 290242 543031 290252
rect 543093 290242 543139 290252
rect 544221 290242 544267 290252
rect 544329 290242 544375 290252
rect 545457 290254 545463 290272
rect 545605 290312 545611 290322
rect 546693 290322 547800 290334
rect 546693 290312 546699 290322
rect 545605 290272 546699 290312
rect 545605 290254 545611 290272
rect 545457 290252 545469 290254
rect 545599 290252 545611 290254
rect 545457 290242 545503 290252
rect 545565 290242 545611 290252
rect 546693 290254 546699 290272
rect 546733 290254 547800 290322
rect 546693 290242 547800 290254
rect 533039 289382 533171 290220
rect 530734 289359 531143 289371
rect 533165 289371 533171 289382
rect 533568 289802 533574 290232
rect 534528 290226 535528 290232
rect 534528 290212 534540 290226
rect 534519 290192 534540 290212
rect 535516 290212 535528 290226
rect 535764 290226 536764 290232
rect 535764 290212 535776 290226
rect 535516 290192 535776 290212
rect 536752 290212 536764 290226
rect 537000 290226 538000 290232
rect 537000 290212 537012 290226
rect 536752 290192 537012 290212
rect 537988 290212 538000 290226
rect 538236 290226 539236 290232
rect 538236 290212 538248 290226
rect 537988 290192 538248 290212
rect 539224 290212 539236 290226
rect 539472 290226 540472 290232
rect 539472 290212 539484 290226
rect 539224 290192 539484 290212
rect 540460 290212 540472 290226
rect 540708 290226 541708 290232
rect 540708 290212 540720 290226
rect 540460 290192 540720 290212
rect 541696 290212 541708 290226
rect 541944 290226 542944 290232
rect 541944 290212 541956 290226
rect 541696 290192 541956 290212
rect 542932 290212 542944 290226
rect 543180 290226 544180 290232
rect 543180 290212 543192 290226
rect 542932 290192 543192 290212
rect 544168 290212 544180 290226
rect 544416 290226 545416 290232
rect 544416 290212 544428 290226
rect 544168 290192 544428 290212
rect 545404 290212 545416 290226
rect 545652 290226 546652 290232
rect 545652 290212 545664 290226
rect 545404 290192 545664 290212
rect 546640 290212 546652 290226
rect 546640 290192 546669 290212
rect 534519 290162 534849 290192
rect 534839 290122 534849 290162
rect 534929 290162 535059 290192
rect 534929 290122 534939 290162
rect 535049 290122 535059 290162
rect 535139 290162 537319 290192
rect 535139 290122 535149 290162
rect 537309 290122 537319 290162
rect 537399 290162 537559 290192
rect 537399 290122 537409 290162
rect 537549 290122 537559 290162
rect 537639 290162 539859 290192
rect 537639 290122 537649 290162
rect 539849 290122 539859 290162
rect 539939 290162 540039 290192
rect 539939 290122 539949 290162
rect 540029 290122 540039 290162
rect 540119 290162 542329 290192
rect 540119 290122 540129 290162
rect 542319 290112 542329 290162
rect 542409 290162 542499 290192
rect 542409 290112 542419 290162
rect 542489 290112 542499 290162
rect 542579 290162 544799 290192
rect 542579 290112 542589 290162
rect 544789 290112 544799 290162
rect 544879 290162 544969 290192
rect 544879 290112 544889 290162
rect 544959 290112 544969 290162
rect 545049 290162 546669 290192
rect 545049 290112 545059 290162
rect 536287 290072 536401 290078
rect 536107 290062 536221 290068
rect 536107 289982 536119 290062
rect 536209 289982 536221 290062
rect 536287 289992 536299 290072
rect 536389 289992 536401 290072
rect 536287 289986 536401 289992
rect 538637 290062 538751 290068
rect 536107 289976 536221 289982
rect 538637 289982 538649 290062
rect 538739 289982 538751 290062
rect 538637 289976 538751 289982
rect 538797 290062 538911 290068
rect 538797 289982 538809 290062
rect 538899 289982 538911 290062
rect 538797 289976 538911 289982
rect 541107 290062 541221 290068
rect 541107 289982 541119 290062
rect 541209 289982 541221 290062
rect 541107 289976 541221 289982
rect 541267 290062 541381 290068
rect 541267 289982 541279 290062
rect 541369 289982 541381 290062
rect 541267 289976 541381 289982
rect 543557 290062 543671 290068
rect 543557 289982 543569 290062
rect 543659 289982 543671 290062
rect 543557 289976 543671 289982
rect 543717 290062 543831 290068
rect 543717 289982 543729 290062
rect 543819 289982 543831 290062
rect 543717 289976 543831 289982
rect 546057 290062 546171 290068
rect 546057 289982 546069 290062
rect 546159 289982 546171 290062
rect 546057 289976 546171 289982
rect 546217 290062 546331 290068
rect 546217 289982 546229 290062
rect 546319 289982 546331 290062
rect 546217 289976 546331 289982
rect 536089 289882 536099 289932
rect 534519 289852 536099 289882
rect 536179 289882 536189 289932
rect 536319 289882 536329 289932
rect 536179 289852 536329 289882
rect 536409 289882 536419 289932
rect 538619 289882 538629 289942
rect 536409 289862 538629 289882
rect 538709 289882 538719 289942
rect 538809 289882 538819 289942
rect 538709 289862 538819 289882
rect 538899 289882 538909 289942
rect 541099 289882 541109 289932
rect 538899 289862 541109 289882
rect 536409 289852 541109 289862
rect 541189 289882 541199 289932
rect 541289 289882 541299 289932
rect 541189 289852 541299 289882
rect 541379 289882 541389 289932
rect 543549 289882 543559 289932
rect 541379 289852 543559 289882
rect 543639 289882 543649 289932
rect 543739 289882 543749 289932
rect 543639 289852 543749 289882
rect 543829 289882 543839 289932
rect 546059 289882 546069 289922
rect 543829 289852 546069 289882
rect 534519 289844 546069 289852
rect 546149 289882 546159 289922
rect 546229 289882 546239 289922
rect 546149 289844 546239 289882
rect 546319 289882 546329 289922
rect 546319 289844 546669 289882
rect 534519 289832 534540 289844
rect 534528 289810 534540 289832
rect 535516 289832 535776 289844
rect 535516 289810 535528 289832
rect 534528 289804 535528 289810
rect 535764 289810 535776 289832
rect 536752 289832 537012 289844
rect 536752 289810 536764 289832
rect 535764 289804 536764 289810
rect 537000 289810 537012 289832
rect 537988 289832 538248 289844
rect 537988 289810 538000 289832
rect 537000 289804 538000 289810
rect 538236 289810 538248 289832
rect 539224 289832 539484 289844
rect 539224 289810 539236 289832
rect 538236 289804 539236 289810
rect 539472 289810 539484 289832
rect 540460 289832 540720 289844
rect 540460 289810 540472 289832
rect 539472 289804 540472 289810
rect 540708 289810 540720 289832
rect 541696 289832 541956 289844
rect 541696 289810 541708 289832
rect 540708 289804 541708 289810
rect 541944 289810 541956 289832
rect 542932 289832 543192 289844
rect 542932 289810 542944 289832
rect 541944 289804 542944 289810
rect 543180 289810 543192 289832
rect 544168 289832 544428 289844
rect 544168 289810 544180 289832
rect 543180 289804 544180 289810
rect 544416 289810 544428 289832
rect 545404 289832 545664 289844
rect 545404 289810 545416 289832
rect 544416 289804 545416 289810
rect 545652 289810 545664 289832
rect 546640 289832 546669 289844
rect 546640 289810 546652 289832
rect 545652 289804 546652 289810
rect 547669 289802 547800 290242
rect 533568 289782 534489 289802
rect 546699 289794 547800 289802
rect 533568 289714 534447 289782
rect 534481 289772 534489 289782
rect 535569 289782 535615 289794
rect 535677 289782 535723 289794
rect 535569 289772 535575 289782
rect 534481 289732 535575 289772
rect 534481 289714 534489 289732
rect 533568 289692 534489 289714
rect 535569 289714 535575 289732
rect 535717 289772 535723 289782
rect 536805 289782 536851 289794
rect 536913 289782 536959 289794
rect 538041 289782 538087 289794
rect 538149 289782 538195 289794
rect 536805 289772 536811 289782
rect 535717 289732 536811 289772
rect 535717 289714 535723 289732
rect 535569 289712 535579 289714
rect 535709 289712 535723 289714
rect 535569 289702 535615 289712
rect 535677 289702 535723 289712
rect 536805 289714 536811 289732
rect 536953 289772 536959 289782
rect 538039 289772 538047 289782
rect 536953 289732 538047 289772
rect 536953 289714 536959 289732
rect 536805 289712 536819 289714
rect 536949 289712 536959 289714
rect 538039 289714 538047 289732
rect 538189 289772 538195 289782
rect 539277 289782 539323 289794
rect 539385 289782 539431 289794
rect 539277 289772 539283 289782
rect 538189 289732 539283 289772
rect 538189 289714 538195 289732
rect 538039 289712 538049 289714
rect 538179 289712 538195 289714
rect 536805 289702 536851 289712
rect 536913 289702 536959 289712
rect 538041 289702 538087 289712
rect 538149 289702 538195 289712
rect 539277 289714 539283 289732
rect 539425 289772 539431 289782
rect 540513 289782 540559 289794
rect 540621 289782 540667 289794
rect 541749 289782 541795 289794
rect 541857 289782 541903 289794
rect 540513 289772 540519 289782
rect 539425 289732 540519 289772
rect 539425 289714 539431 289732
rect 539277 289712 539289 289714
rect 539419 289712 539431 289714
rect 539277 289702 539323 289712
rect 539385 289702 539431 289712
rect 540513 289714 540519 289732
rect 540661 289772 540669 289782
rect 541749 289772 541755 289782
rect 540661 289732 541755 289772
rect 540661 289714 540669 289732
rect 540513 289712 540529 289714
rect 540659 289712 540669 289714
rect 541749 289714 541755 289732
rect 541897 289772 541903 289782
rect 542985 289782 543031 289794
rect 543093 289782 543139 289794
rect 544221 289782 544267 289794
rect 544329 289782 544375 289794
rect 542985 289772 542991 289782
rect 541897 289732 542991 289772
rect 541897 289714 541903 289732
rect 541749 289712 541759 289714
rect 541889 289712 541903 289714
rect 540513 289702 540559 289712
rect 540621 289702 540667 289712
rect 541749 289702 541795 289712
rect 541857 289702 541903 289712
rect 542985 289714 542991 289732
rect 543133 289772 543139 289782
rect 544219 289772 544227 289782
rect 543133 289732 544227 289772
rect 543133 289714 543139 289732
rect 542985 289712 542999 289714
rect 543129 289712 543139 289714
rect 544219 289714 544227 289732
rect 544369 289772 544375 289782
rect 545457 289782 545503 289794
rect 545565 289782 545611 289794
rect 545457 289772 545463 289782
rect 544369 289732 545463 289772
rect 544369 289714 544375 289732
rect 544219 289712 544229 289714
rect 544359 289712 544375 289714
rect 542985 289702 543031 289712
rect 543093 289702 543139 289712
rect 544221 289702 544267 289712
rect 544329 289702 544375 289712
rect 545457 289714 545463 289732
rect 545605 289772 545611 289782
rect 546693 289782 547800 289794
rect 546693 289772 546699 289782
rect 545605 289732 546699 289772
rect 545605 289714 545611 289732
rect 545457 289712 545469 289714
rect 545599 289712 545611 289714
rect 545457 289702 545503 289712
rect 545565 289702 545611 289712
rect 546693 289714 546699 289732
rect 546733 289714 547800 289782
rect 546693 289702 547800 289714
rect 533568 289371 533574 289692
rect 534528 289686 535528 289692
rect 534528 289672 534540 289686
rect 534519 289652 534540 289672
rect 535516 289672 535528 289686
rect 535764 289686 536764 289692
rect 535764 289672 535776 289686
rect 535516 289652 535776 289672
rect 536752 289672 536764 289686
rect 537000 289686 538000 289692
rect 537000 289672 537012 289686
rect 536752 289652 537012 289672
rect 537988 289672 538000 289686
rect 538236 289686 539236 289692
rect 538236 289672 538248 289686
rect 537988 289652 538248 289672
rect 539224 289672 539236 289686
rect 539472 289686 540472 289692
rect 539472 289672 539484 289686
rect 539224 289652 539484 289672
rect 540460 289672 540472 289686
rect 540708 289686 541708 289692
rect 540708 289672 540720 289686
rect 540460 289652 540720 289672
rect 541696 289672 541708 289686
rect 541944 289686 542944 289692
rect 541944 289672 541956 289686
rect 541696 289652 541956 289672
rect 542932 289672 542944 289686
rect 543180 289686 544180 289692
rect 543180 289672 543192 289686
rect 542932 289652 543192 289672
rect 544168 289672 544180 289686
rect 544416 289686 545416 289692
rect 544416 289672 544428 289686
rect 544168 289652 544428 289672
rect 545404 289672 545416 289686
rect 545652 289686 546652 289692
rect 545652 289672 545664 289686
rect 545404 289652 545664 289672
rect 546640 289672 546652 289686
rect 546640 289652 546669 289672
rect 534519 289622 534849 289652
rect 534839 289582 534849 289622
rect 534929 289622 535059 289652
rect 534929 289582 534939 289622
rect 535049 289582 535059 289622
rect 535139 289622 537319 289652
rect 535139 289582 535149 289622
rect 537309 289572 537319 289622
rect 537399 289622 537559 289652
rect 537399 289572 537409 289622
rect 537549 289572 537559 289622
rect 537639 289622 539859 289652
rect 537639 289572 537649 289622
rect 539849 289582 539859 289622
rect 539939 289622 540049 289652
rect 539939 289582 539949 289622
rect 540039 289582 540049 289622
rect 540129 289622 542319 289652
rect 540129 289582 540139 289622
rect 542309 289572 542319 289622
rect 542399 289622 542509 289652
rect 542399 289572 542409 289622
rect 542499 289572 542509 289622
rect 542589 289642 546669 289652
rect 542589 289622 544799 289642
rect 542589 289572 542599 289622
rect 544789 289562 544799 289622
rect 544879 289622 544969 289642
rect 544879 289562 544889 289622
rect 544959 289562 544969 289622
rect 545049 289622 546669 289642
rect 545049 289562 545059 289622
rect 547669 289382 547800 289702
rect 533165 289359 533574 289371
rect 547794 289371 547800 289382
rect 548197 289371 548203 290485
rect 547794 289359 548203 289371
rect 550109 290485 550634 290497
rect 550109 289371 550231 290485
rect 550628 289371 550634 290485
rect 550109 289362 550634 289371
rect 550225 289359 550634 289362
rect 531753 289252 531855 289264
rect 531963 289252 532065 289264
rect 531749 289122 531759 289252
rect 531849 289122 531859 289252
rect 531959 289122 531969 289252
rect 532059 289122 532069 289252
rect 549063 289242 549145 289254
rect 549223 289242 549305 289254
rect 549059 289152 549069 289242
rect 549139 289152 549149 289242
rect 549219 289152 549229 289242
rect 549299 289152 549309 289242
rect 538359 289132 538589 289142
rect 531753 289110 531855 289122
rect 531963 289110 532065 289122
rect 536809 289082 536819 289132
rect 536449 289064 536819 289082
rect 536949 289082 536959 289132
rect 538129 289122 538229 289132
rect 538039 289082 538049 289122
rect 536949 289064 538049 289082
rect 538179 289082 538229 289122
rect 538359 289082 538379 289132
rect 538179 289064 538379 289082
rect 538459 289064 538489 289132
rect 538569 289082 538589 289132
rect 540549 289122 540649 289152
rect 540769 289132 540999 289152
rect 543229 289142 543459 289152
rect 539279 289082 539289 289122
rect 538569 289064 539289 289082
rect 539419 289082 539429 289122
rect 540519 289082 540529 289122
rect 539419 289064 540529 289082
rect 540659 289082 540669 289122
rect 540769 289082 540789 289132
rect 540659 289064 540789 289082
rect 540869 289064 540899 289132
rect 540979 289082 540999 289132
rect 541749 289082 541759 289122
rect 540979 289064 541759 289082
rect 541889 289082 541899 289122
rect 542979 289082 542999 289142
rect 541889 289072 542999 289082
rect 543129 289082 543139 289142
rect 543229 289082 543249 289142
rect 543129 289072 543249 289082
rect 541889 289064 543249 289072
rect 543329 289064 543359 289142
rect 543439 289082 543459 289142
rect 549063 289140 549145 289152
rect 549223 289140 549305 289152
rect 544219 289082 544229 289122
rect 543439 289064 544229 289082
rect 544359 289082 544369 289122
rect 544359 289064 544779 289082
rect 562260 289080 567820 293300
rect 536449 289042 536471 289064
rect 536459 289030 536471 289042
rect 537447 289042 537689 289064
rect 537447 289030 537459 289042
rect 536459 289024 537459 289030
rect 537677 289030 537689 289042
rect 538665 289042 538907 289064
rect 538665 289030 538677 289042
rect 537677 289024 538677 289030
rect 538895 289030 538907 289042
rect 539883 289042 540125 289064
rect 539883 289030 539895 289042
rect 538895 289024 539895 289030
rect 540113 289030 540125 289042
rect 541101 289042 541343 289064
rect 541101 289030 541113 289042
rect 540113 289024 541113 289030
rect 541331 289030 541343 289042
rect 542319 289042 542561 289064
rect 542319 289030 542331 289042
rect 541331 289024 542331 289030
rect 542549 289030 542561 289042
rect 543537 289042 543779 289064
rect 543537 289030 543549 289042
rect 542549 289024 543549 289030
rect 543767 289030 543779 289042
rect 544755 289042 544779 289064
rect 544755 289030 544767 289042
rect 543767 289024 544767 289030
rect 544820 289014 567820 289080
rect 536381 289002 536427 289014
rect 536381 288992 536387 289002
rect 536379 288952 536387 288992
rect 536381 288934 536387 288952
rect 536421 288992 536427 289002
rect 537491 289002 537537 289014
rect 537491 288992 537497 289002
rect 536421 288952 537497 288992
rect 536421 288934 536427 288952
rect 536381 288922 536427 288934
rect 537491 288934 537497 288952
rect 537531 288992 537537 289002
rect 537599 289002 537645 289014
rect 537599 288992 537605 289002
rect 537531 288952 537605 288992
rect 537531 288934 537537 288952
rect 537491 288922 537537 288934
rect 537599 288934 537605 288952
rect 537639 288992 537645 289002
rect 538709 289002 538755 289014
rect 538817 289002 538863 289014
rect 538709 288992 538715 289002
rect 537639 288952 538715 288992
rect 537639 288934 537645 288952
rect 537599 288922 537645 288934
rect 538709 288934 538715 288952
rect 538749 288934 538823 289002
rect 538857 288992 538863 289002
rect 539927 289002 539973 289014
rect 540035 289002 540081 289014
rect 539927 288992 539933 289002
rect 538857 288952 539933 288992
rect 538857 288934 538863 288952
rect 538709 288932 538863 288934
rect 538709 288922 538755 288932
rect 538817 288922 538863 288932
rect 539927 288934 539933 288952
rect 539967 288934 540041 289002
rect 540075 288992 540081 289002
rect 541145 289002 541191 289014
rect 541253 289002 541299 289014
rect 541145 288992 541151 289002
rect 540075 288952 541151 288992
rect 540075 288934 540081 288952
rect 539927 288932 540081 288934
rect 539927 288922 539973 288932
rect 540035 288922 540081 288932
rect 541145 288934 541151 288952
rect 541185 288934 541259 289002
rect 541293 288992 541299 289002
rect 542363 289002 542409 289014
rect 542471 289002 542517 289014
rect 543581 289002 543627 289014
rect 543689 289002 543735 289014
rect 542363 288992 542369 289002
rect 541293 288952 542369 288992
rect 541293 288934 541299 288952
rect 541145 288932 541299 288934
rect 541145 288922 541191 288932
rect 541253 288922 541299 288932
rect 542363 288934 542369 288952
rect 542403 288934 542477 289002
rect 542511 288992 542519 289002
rect 543579 288992 543587 289002
rect 542511 288952 543587 288992
rect 542511 288934 542519 288952
rect 542363 288932 542519 288934
rect 543579 288934 543587 288952
rect 543621 288934 543695 289002
rect 543729 288992 543735 289002
rect 544799 289002 567820 289014
rect 544799 288992 544805 289002
rect 543729 288952 544805 288992
rect 543729 288934 543735 288952
rect 543579 288932 543735 288934
rect 542363 288922 542409 288932
rect 542471 288922 542517 288932
rect 543581 288922 543627 288932
rect 543689 288922 543735 288932
rect 544799 288934 544805 288952
rect 544839 288934 567820 289002
rect 544799 288922 567820 288934
rect 536459 288906 537459 288912
rect 536459 288892 536471 288906
rect 536449 288872 536471 288892
rect 537447 288892 537459 288906
rect 537677 288906 538677 288912
rect 537677 288892 537689 288906
rect 537447 288872 537689 288892
rect 538665 288892 538677 288906
rect 538895 288906 539895 288912
rect 538895 288892 538907 288906
rect 538665 288872 538907 288892
rect 539883 288892 539895 288906
rect 540113 288906 541113 288912
rect 540113 288892 540125 288906
rect 539883 288872 540125 288892
rect 541101 288892 541113 288906
rect 541331 288906 542331 288912
rect 541331 288892 541343 288906
rect 541101 288872 541343 288892
rect 542319 288892 542331 288906
rect 542549 288906 543549 288912
rect 542549 288892 542561 288906
rect 542319 288872 542561 288892
rect 543537 288892 543549 288906
rect 543767 288906 544767 288912
rect 543767 288892 543779 288906
rect 543537 288872 543779 288892
rect 544755 288892 544767 288906
rect 544755 288872 544779 288892
rect 536449 288862 541769 288872
rect 536449 288852 536759 288862
rect 536749 288782 536759 288852
rect 536849 288782 536899 288862
rect 536989 288852 541769 288862
rect 536989 288782 536999 288852
rect 539339 288802 539439 288852
rect 541759 288802 541769 288852
rect 541859 288802 541909 288872
rect 541999 288852 544779 288872
rect 544820 288860 567820 288922
rect 568110 288858 578380 288864
rect 541999 288802 542009 288852
rect 536759 288632 536989 288782
rect 538267 288772 538401 288778
rect 538267 288662 538279 288772
rect 538389 288662 538401 288772
rect 538267 288656 538401 288662
rect 539127 288772 539261 288778
rect 539127 288662 539139 288772
rect 539249 288662 539261 288772
rect 539127 288656 539261 288662
rect 540337 288772 540471 288778
rect 540337 288662 540349 288772
rect 540459 288662 540471 288772
rect 540337 288656 540471 288662
rect 541187 288772 541321 288778
rect 541187 288662 541199 288772
rect 541309 288662 541321 288772
rect 541187 288656 541321 288662
rect 536749 288582 536759 288632
rect 536449 288564 536759 288582
rect 536849 288564 536899 288632
rect 536989 288582 536999 288632
rect 538129 288582 538229 288632
rect 540549 288582 540649 288652
rect 541769 288622 541999 288802
rect 544219 288792 544319 288852
rect 568110 288824 570720 288858
rect 575860 288824 578380 288858
rect 568110 288814 578380 288824
rect 542757 288772 542891 288778
rect 542757 288662 542769 288772
rect 542879 288662 542891 288772
rect 542757 288656 542891 288662
rect 543637 288772 543771 288778
rect 543637 288662 543649 288772
rect 543759 288662 543771 288772
rect 543637 288656 543771 288662
rect 541759 288582 541769 288622
rect 536989 288564 541769 288582
rect 541859 288564 541909 288622
rect 541999 288582 542009 288622
rect 542979 288582 543079 288642
rect 541999 288564 544779 288582
rect 536449 288542 536471 288564
rect 536459 288530 536471 288542
rect 537447 288542 537689 288564
rect 537447 288530 537459 288542
rect 536459 288524 537459 288530
rect 537677 288530 537689 288542
rect 538665 288542 538907 288564
rect 538665 288530 538677 288542
rect 537677 288524 538677 288530
rect 538895 288530 538907 288542
rect 539883 288542 540125 288564
rect 539883 288530 539895 288542
rect 538895 288524 539895 288530
rect 540113 288530 540125 288542
rect 541101 288542 541343 288564
rect 542319 288542 542561 288564
rect 541101 288530 541113 288542
rect 540113 288524 541113 288530
rect 541331 288530 541343 288542
rect 542319 288530 542331 288542
rect 541331 288524 542331 288530
rect 542549 288530 542561 288542
rect 543537 288542 543779 288564
rect 543537 288530 543549 288542
rect 542549 288524 543549 288530
rect 543767 288530 543779 288542
rect 544755 288542 544779 288564
rect 544755 288530 544767 288542
rect 543767 288524 544767 288530
rect 544820 288514 550960 288580
rect 536381 288502 536427 288514
rect 536381 288434 536387 288502
rect 536421 288492 536427 288502
rect 537491 288502 537537 288514
rect 537491 288492 537497 288502
rect 536421 288452 537497 288492
rect 536421 288434 536427 288452
rect 536381 288422 536427 288434
rect 537491 288434 537497 288452
rect 537531 288492 537537 288502
rect 537599 288502 537645 288514
rect 537599 288492 537605 288502
rect 537531 288452 537605 288492
rect 537531 288434 537537 288452
rect 537491 288422 537537 288434
rect 537599 288434 537605 288452
rect 537639 288492 537645 288502
rect 538709 288502 538755 288514
rect 538817 288502 538863 288514
rect 538709 288492 538715 288502
rect 537639 288452 538715 288492
rect 537639 288434 537645 288452
rect 537599 288422 537645 288434
rect 538709 288434 538715 288452
rect 538749 288434 538823 288502
rect 538857 288492 538863 288502
rect 539927 288502 539973 288514
rect 540035 288502 540081 288514
rect 539927 288492 539933 288502
rect 538857 288452 539933 288492
rect 538857 288434 538863 288452
rect 538709 288432 538863 288434
rect 538709 288422 538755 288432
rect 538817 288422 538863 288432
rect 539927 288434 539933 288452
rect 539967 288434 540041 288502
rect 540075 288492 540081 288502
rect 541145 288502 541191 288514
rect 541253 288502 541299 288514
rect 541145 288492 541151 288502
rect 540075 288452 541151 288492
rect 540075 288434 540081 288452
rect 539927 288432 540081 288434
rect 539927 288422 539973 288432
rect 540035 288422 540081 288432
rect 541145 288434 541151 288452
rect 541185 288434 541259 288502
rect 541293 288492 541299 288502
rect 542363 288502 542409 288514
rect 542471 288502 542517 288514
rect 543581 288502 543627 288514
rect 543689 288502 543735 288514
rect 542363 288492 542369 288502
rect 541293 288452 542369 288492
rect 541293 288434 541299 288452
rect 541145 288432 541299 288434
rect 541145 288422 541191 288432
rect 541253 288422 541299 288432
rect 542363 288434 542369 288452
rect 542403 288434 542477 288502
rect 542511 288492 542519 288502
rect 543579 288492 543587 288502
rect 542511 288452 543587 288492
rect 542511 288434 542519 288452
rect 542363 288432 542519 288434
rect 543579 288434 543587 288452
rect 543621 288434 543695 288502
rect 543729 288492 543735 288502
rect 544799 288502 550960 288514
rect 544799 288492 544805 288502
rect 543729 288452 544805 288492
rect 543729 288434 543735 288452
rect 543579 288432 543735 288434
rect 542363 288422 542409 288432
rect 542471 288422 542517 288432
rect 543581 288422 543627 288432
rect 543689 288422 543735 288432
rect 544799 288434 544805 288452
rect 544839 288434 550960 288502
rect 544799 288422 550960 288434
rect 536459 288406 537459 288412
rect 536459 288392 536471 288406
rect 536449 288372 536471 288392
rect 537447 288392 537459 288406
rect 537677 288406 538677 288412
rect 537677 288392 537689 288406
rect 537447 288372 537689 288392
rect 538665 288392 538677 288406
rect 538895 288406 539895 288412
rect 538895 288392 538907 288406
rect 539883 288392 539895 288406
rect 540113 288406 541113 288412
rect 540113 288392 540125 288406
rect 538665 288372 538907 288392
rect 539883 288372 540125 288392
rect 541101 288392 541113 288406
rect 541331 288406 542331 288412
rect 541331 288392 541343 288406
rect 542319 288392 542331 288406
rect 542549 288406 543549 288412
rect 542549 288392 542561 288406
rect 541101 288372 541343 288392
rect 542319 288372 542561 288392
rect 543537 288392 543549 288406
rect 543767 288406 544767 288412
rect 543767 288392 543779 288406
rect 543537 288372 543779 288392
rect 544755 288392 544767 288406
rect 544755 288372 544779 288392
rect 536449 288352 537089 288372
rect 536889 288302 536989 288352
rect 537079 288292 537089 288352
rect 537169 288352 537239 288372
rect 537169 288292 537179 288352
rect 537229 288292 537239 288352
rect 537319 288352 539579 288372
rect 537319 288292 537329 288352
rect 538039 288332 538189 288352
rect 539279 288322 539439 288352
rect 539339 288302 539439 288322
rect 539569 288312 539579 288352
rect 539659 288352 539729 288372
rect 539659 288312 539669 288352
rect 539719 288312 539729 288352
rect 539809 288352 542059 288372
rect 539809 288312 539819 288352
rect 540519 288322 540669 288352
rect 541779 288292 541879 288352
rect 542049 288312 542059 288352
rect 542139 288352 542199 288372
rect 542139 288312 542149 288352
rect 542189 288312 542199 288352
rect 542279 288352 544779 288372
rect 544820 288360 550960 288422
rect 542279 288312 542289 288352
rect 542989 288322 543139 288352
rect 544219 288322 544369 288352
rect 544219 288292 544319 288322
rect 537449 288142 537759 288172
rect 537329 288082 537539 288142
rect 537009 288064 537539 288082
rect 537619 288064 537649 288142
rect 537729 288082 537759 288142
rect 542389 288132 542609 288142
rect 539939 288082 539949 288112
rect 537729 288064 539949 288082
rect 540029 288082 540039 288112
rect 542389 288082 542399 288132
rect 540029 288064 542399 288082
rect 542479 288064 542519 288132
rect 542599 288082 542609 288132
rect 543589 288082 543599 288122
rect 542599 288064 543599 288082
rect 543679 288082 543689 288122
rect 543679 288064 544129 288082
rect 537009 288042 537031 288064
rect 537019 288030 537031 288042
rect 538007 288042 538249 288064
rect 538007 288030 538019 288042
rect 537019 288024 538019 288030
rect 538237 288030 538249 288042
rect 539225 288042 539467 288064
rect 539225 288030 539237 288042
rect 538237 288024 539237 288030
rect 539455 288030 539467 288042
rect 540443 288042 540685 288064
rect 540443 288030 540455 288042
rect 539455 288024 540455 288030
rect 540673 288030 540685 288042
rect 541661 288042 541903 288064
rect 541661 288030 541673 288042
rect 540673 288024 541673 288030
rect 541891 288030 541903 288042
rect 542879 288042 543121 288064
rect 544097 288042 544129 288064
rect 542879 288030 542891 288042
rect 541891 288024 542891 288030
rect 543109 288030 543121 288042
rect 544097 288030 544109 288042
rect 543109 288024 544109 288030
rect 536941 288002 536987 288014
rect 536941 287982 536947 288002
rect 536929 287862 536947 287982
rect 536941 287834 536947 287862
rect 536981 287982 536987 288002
rect 538051 288002 538097 288014
rect 538051 287982 538057 288002
rect 536981 287862 538057 287982
rect 536981 287834 536987 287862
rect 536941 287822 536987 287834
rect 538051 287834 538057 287862
rect 538091 287982 538097 288002
rect 538159 288002 538205 288014
rect 538159 287982 538165 288002
rect 538091 287862 538165 287982
rect 538091 287834 538097 287862
rect 538051 287822 538097 287834
rect 538159 287834 538165 287862
rect 538199 287982 538205 288002
rect 539269 288002 539315 288014
rect 539269 287982 539275 288002
rect 538199 287962 539275 287982
rect 538199 287882 538719 287962
rect 538799 287882 539275 287962
rect 538199 287862 539275 287882
rect 538199 287834 538205 287862
rect 538159 287822 538205 287834
rect 539269 287834 539275 287862
rect 539309 287982 539315 288002
rect 539377 288002 539423 288014
rect 539377 287982 539383 288002
rect 539309 287862 539383 287982
rect 539309 287834 539315 287862
rect 539269 287822 539315 287834
rect 539377 287834 539383 287862
rect 539417 287982 539423 288002
rect 540487 288002 540533 288014
rect 540487 287982 540493 288002
rect 539417 287862 540493 287982
rect 539417 287834 539423 287862
rect 539377 287822 539423 287834
rect 540487 287834 540493 287862
rect 540527 287982 540533 288002
rect 540595 288002 540641 288014
rect 540595 287982 540601 288002
rect 540527 287862 540601 287982
rect 540527 287834 540533 287862
rect 540487 287822 540533 287834
rect 540595 287834 540601 287862
rect 540635 287982 540641 288002
rect 541705 288002 541751 288014
rect 541705 287982 541711 288002
rect 540635 287962 541711 287982
rect 540635 287882 541129 287962
rect 541209 287882 541711 287962
rect 540635 287862 541711 287882
rect 540635 287834 540641 287862
rect 540595 287822 540641 287834
rect 541705 287834 541711 287862
rect 541745 287982 541751 288002
rect 541813 288002 541859 288014
rect 541813 287982 541819 288002
rect 541745 287862 541819 287982
rect 541745 287834 541751 287862
rect 541705 287822 541751 287834
rect 541813 287834 541819 287862
rect 541853 287982 541859 288002
rect 542923 288002 542969 288014
rect 542923 287982 542929 288002
rect 541853 287862 542929 287982
rect 541853 287834 541859 287862
rect 541813 287822 541859 287834
rect 542923 287834 542929 287862
rect 542963 287982 542969 288002
rect 543031 288002 543077 288014
rect 543031 287982 543037 288002
rect 542963 287862 543037 287982
rect 542963 287834 542969 287862
rect 542923 287822 542969 287834
rect 543031 287834 543037 287862
rect 543071 287982 543077 288002
rect 544141 288002 544187 288014
rect 544141 287982 544147 288002
rect 543071 287862 544147 287982
rect 543071 287834 543077 287862
rect 543031 287822 543077 287834
rect 544141 287834 544147 287862
rect 544181 287834 544187 288002
rect 544141 287822 544187 287834
rect 537019 287806 538019 287812
rect 537019 287782 537031 287806
rect 538007 287782 538019 287806
rect 538237 287806 539237 287812
rect 538237 287782 538249 287806
rect 537009 287772 537031 287782
rect 538007 287772 538249 287782
rect 539225 287782 539237 287806
rect 539455 287806 540455 287812
rect 539455 287782 539467 287806
rect 539225 287772 539467 287782
rect 540443 287782 540455 287806
rect 540673 287806 541673 287812
rect 540673 287782 540685 287806
rect 540443 287772 540685 287782
rect 541661 287782 541673 287806
rect 541891 287806 542891 287812
rect 541891 287782 541903 287806
rect 542879 287782 542891 287806
rect 543109 287806 544109 287812
rect 543109 287782 543121 287806
rect 541661 287772 541903 287782
rect 542879 287772 543121 287782
rect 544097 287782 544109 287806
rect 544097 287772 544129 287782
rect 537009 287742 537459 287772
rect 537449 287702 537459 287742
rect 537539 287742 542349 287772
rect 537539 287702 537549 287742
rect 542339 287702 542349 287742
rect 542429 287742 544129 287772
rect 542429 287702 542439 287742
rect 537557 287652 537691 287658
rect 537557 287562 537569 287652
rect 537679 287562 537691 287652
rect 537557 287556 537691 287562
rect 542467 287652 542601 287658
rect 542467 287562 542479 287652
rect 542589 287562 542601 287652
rect 542467 287556 542601 287562
rect 539939 287462 539949 287492
rect 537009 287444 539949 287462
rect 540029 287462 540039 287492
rect 543589 287462 543599 287502
rect 540029 287444 543599 287462
rect 543679 287462 543689 287502
rect 543679 287444 544129 287462
rect 537009 287422 537031 287444
rect 537019 287410 537031 287422
rect 538007 287422 538249 287444
rect 538007 287410 538019 287422
rect 537019 287404 538019 287410
rect 538237 287410 538249 287422
rect 539225 287422 539467 287444
rect 539225 287410 539237 287422
rect 538237 287404 539237 287410
rect 539455 287410 539467 287422
rect 540443 287422 540685 287444
rect 540443 287410 540455 287422
rect 539455 287404 540455 287410
rect 540673 287410 540685 287422
rect 541661 287422 541903 287444
rect 541661 287410 541673 287422
rect 540673 287404 541673 287410
rect 541891 287410 541903 287422
rect 542879 287422 543121 287444
rect 544097 287422 544129 287444
rect 542879 287410 542891 287422
rect 541891 287404 542891 287410
rect 543109 287410 543121 287422
rect 544097 287410 544109 287422
rect 543109 287404 544109 287410
rect 536941 287382 536987 287394
rect 536941 287352 536947 287382
rect 536909 287252 536947 287352
rect 536941 287214 536947 287252
rect 536981 287362 536987 287382
rect 538051 287382 538097 287394
rect 538051 287362 538057 287382
rect 536981 287242 538057 287362
rect 536981 287214 536987 287242
rect 536941 287202 536987 287214
rect 538051 287214 538057 287242
rect 538091 287362 538097 287382
rect 538159 287382 538205 287394
rect 538159 287362 538165 287382
rect 538091 287342 538165 287362
rect 538199 287362 538205 287382
rect 539269 287382 539315 287394
rect 539269 287362 539275 287382
rect 538199 287342 539275 287362
rect 538091 287262 538109 287342
rect 538199 287262 538229 287342
rect 538319 287262 538719 287342
rect 538799 287262 539275 287342
rect 538091 287242 538165 287262
rect 538091 287214 538097 287242
rect 538051 287202 538097 287214
rect 538159 287214 538165 287242
rect 538199 287242 539275 287262
rect 538199 287214 538205 287242
rect 538159 287202 538205 287214
rect 539269 287214 539275 287242
rect 539309 287362 539315 287382
rect 539377 287382 539423 287394
rect 539377 287362 539383 287382
rect 539309 287242 539383 287362
rect 539309 287214 539315 287242
rect 539269 287202 539315 287214
rect 539377 287214 539383 287242
rect 539417 287362 539423 287382
rect 540487 287382 540533 287394
rect 540487 287362 540493 287382
rect 539417 287242 540493 287362
rect 539417 287214 539423 287242
rect 539377 287202 539423 287214
rect 540487 287214 540493 287242
rect 540527 287362 540533 287382
rect 540595 287382 540641 287394
rect 540595 287362 540601 287382
rect 540527 287342 540601 287362
rect 540635 287362 540641 287382
rect 541705 287382 541751 287394
rect 541705 287362 541711 287382
rect 540635 287342 541711 287362
rect 540527 287262 540559 287342
rect 540649 287262 540679 287342
rect 540769 287262 541129 287342
rect 541209 287262 541711 287342
rect 540527 287242 540601 287262
rect 540527 287214 540533 287242
rect 540487 287202 540533 287214
rect 540595 287214 540601 287242
rect 540635 287242 541711 287262
rect 540635 287214 540641 287242
rect 540595 287202 540641 287214
rect 541705 287214 541711 287242
rect 541745 287362 541751 287382
rect 541813 287382 541859 287394
rect 541813 287362 541819 287382
rect 541745 287242 541819 287362
rect 541745 287214 541751 287242
rect 541705 287202 541751 287214
rect 541813 287214 541819 287242
rect 541853 287362 541859 287382
rect 542923 287382 542969 287394
rect 542923 287362 542929 287382
rect 541853 287242 542929 287362
rect 541853 287214 541859 287242
rect 541813 287202 541859 287214
rect 542923 287214 542929 287242
rect 542963 287362 542969 287382
rect 543031 287382 543077 287394
rect 543031 287362 543037 287382
rect 542963 287342 543037 287362
rect 543071 287362 543077 287382
rect 544141 287382 544187 287394
rect 544141 287362 544147 287382
rect 543071 287342 544147 287362
rect 542963 287262 542989 287342
rect 543079 287262 543109 287342
rect 543199 287262 544147 287342
rect 542963 287242 543037 287262
rect 542963 287214 542969 287242
rect 542923 287202 542969 287214
rect 543031 287214 543037 287242
rect 543071 287242 544147 287262
rect 543071 287214 543077 287242
rect 543031 287202 543077 287214
rect 544141 287214 544147 287242
rect 544181 287362 544187 287382
rect 544181 287242 544189 287362
rect 544181 287214 544187 287242
rect 544141 287202 544187 287214
rect 537019 287186 538019 287192
rect 537019 287162 537031 287186
rect 538007 287162 538019 287186
rect 538237 287186 539237 287192
rect 538237 287162 538249 287186
rect 537009 287152 537031 287162
rect 538007 287152 538249 287162
rect 539225 287162 539237 287186
rect 539455 287186 540455 287192
rect 539455 287162 539467 287186
rect 539225 287152 539467 287162
rect 540443 287162 540455 287186
rect 540673 287186 541673 287192
rect 540673 287162 540685 287186
rect 540443 287152 540685 287162
rect 541661 287162 541673 287186
rect 541891 287186 542891 287192
rect 541891 287162 541903 287186
rect 542879 287162 542891 287186
rect 543109 287186 544109 287192
rect 543109 287162 543121 287186
rect 541661 287152 541903 287162
rect 542879 287152 543121 287162
rect 544097 287162 544109 287186
rect 544097 287152 544129 287162
rect 537009 287122 537459 287152
rect 537449 287082 537459 287122
rect 537539 287122 542349 287152
rect 537539 287082 537549 287122
rect 542339 287082 542349 287122
rect 542429 287122 544129 287152
rect 542429 287082 542439 287122
rect 539329 286882 539339 286912
rect 536449 286844 539339 286882
rect 539429 286882 539439 286912
rect 544209 286882 544219 286932
rect 539429 286852 544219 286882
rect 544309 286882 544319 286932
rect 544309 286852 544769 286882
rect 539429 286844 544769 286852
rect 536449 286842 536471 286844
rect 536459 286810 536471 286842
rect 537447 286842 537689 286844
rect 537447 286810 537459 286842
rect 536459 286804 537459 286810
rect 537677 286810 537689 286842
rect 538665 286842 538907 286844
rect 538665 286810 538677 286842
rect 537677 286804 538677 286810
rect 538895 286810 538907 286842
rect 539883 286842 540125 286844
rect 539883 286810 539895 286842
rect 538895 286804 539895 286810
rect 540113 286810 540125 286842
rect 541101 286842 541343 286844
rect 541101 286810 541113 286842
rect 540113 286804 541113 286810
rect 541331 286810 541343 286842
rect 542319 286842 542561 286844
rect 542319 286810 542331 286842
rect 541331 286804 542331 286810
rect 542549 286810 542561 286842
rect 543537 286842 543779 286844
rect 543537 286810 543549 286842
rect 542549 286804 543549 286810
rect 543767 286810 543779 286842
rect 544755 286842 544769 286844
rect 544755 286810 544767 286842
rect 543767 286804 544767 286810
rect 536381 286782 536427 286794
rect 536381 286762 536387 286782
rect 536369 286642 536387 286762
rect 536381 286614 536387 286642
rect 536421 286762 536427 286782
rect 537491 286782 537537 286794
rect 537491 286762 537497 286782
rect 536421 286642 537497 286762
rect 536421 286614 536427 286642
rect 536381 286602 536427 286614
rect 537491 286614 537497 286642
rect 537531 286762 537537 286782
rect 537599 286782 537645 286794
rect 537599 286762 537605 286782
rect 537531 286642 537605 286762
rect 537531 286614 537537 286642
rect 537491 286602 537537 286614
rect 537599 286614 537605 286642
rect 537639 286762 537645 286782
rect 538709 286782 538755 286794
rect 538709 286762 538715 286782
rect 537639 286742 538715 286762
rect 537639 286662 538109 286742
rect 538199 286662 538229 286742
rect 538319 286662 538715 286742
rect 537639 286642 538715 286662
rect 537639 286614 537645 286642
rect 537599 286602 537645 286614
rect 538709 286614 538715 286642
rect 538749 286762 538755 286782
rect 538817 286782 538863 286794
rect 538817 286762 538823 286782
rect 538749 286642 538823 286762
rect 538749 286614 538755 286642
rect 538709 286602 538755 286614
rect 538817 286614 538823 286642
rect 538857 286762 538863 286782
rect 539927 286782 539973 286794
rect 539927 286762 539933 286782
rect 538857 286642 539933 286762
rect 538857 286614 538863 286642
rect 538817 286602 538863 286614
rect 539927 286614 539933 286642
rect 539967 286762 539973 286782
rect 540035 286782 540081 286794
rect 540035 286762 540041 286782
rect 539967 286642 540041 286762
rect 539967 286614 539973 286642
rect 539927 286602 539973 286614
rect 540035 286614 540041 286642
rect 540075 286762 540081 286782
rect 541145 286782 541191 286794
rect 541145 286762 541151 286782
rect 540075 286742 541151 286762
rect 540075 286662 540559 286742
rect 540649 286662 540679 286742
rect 540769 286662 541151 286742
rect 540075 286642 541151 286662
rect 540075 286614 540081 286642
rect 540035 286602 540081 286614
rect 541145 286614 541151 286642
rect 541185 286762 541191 286782
rect 541253 286782 541299 286794
rect 541253 286762 541259 286782
rect 541185 286642 541259 286762
rect 541185 286614 541191 286642
rect 541145 286602 541191 286614
rect 541253 286614 541259 286642
rect 541293 286762 541299 286782
rect 542363 286782 542409 286794
rect 542363 286762 542369 286782
rect 541293 286642 542369 286762
rect 541293 286614 541299 286642
rect 541253 286602 541299 286614
rect 542363 286614 542369 286642
rect 542403 286762 542409 286782
rect 542471 286782 542517 286794
rect 542471 286762 542477 286782
rect 542403 286642 542477 286762
rect 542403 286614 542409 286642
rect 542363 286602 542409 286614
rect 542471 286614 542477 286642
rect 542511 286762 542517 286782
rect 543581 286782 543627 286794
rect 543581 286762 543587 286782
rect 542511 286742 543587 286762
rect 542511 286662 542989 286742
rect 543079 286662 543109 286742
rect 543199 286662 543587 286742
rect 542511 286642 543587 286662
rect 542511 286614 542517 286642
rect 542471 286602 542517 286614
rect 543581 286614 543587 286642
rect 543621 286762 543627 286782
rect 543689 286782 543735 286794
rect 543689 286762 543695 286782
rect 543621 286642 543695 286762
rect 543621 286614 543627 286642
rect 543581 286602 543627 286614
rect 543689 286614 543695 286642
rect 543729 286762 543735 286782
rect 544799 286782 544845 286794
rect 544799 286762 544805 286782
rect 543729 286642 544805 286762
rect 543729 286614 543735 286642
rect 543689 286602 543735 286614
rect 544799 286614 544805 286642
rect 544839 286762 544845 286782
rect 544839 286642 544849 286762
rect 544839 286614 544845 286642
rect 544799 286602 544845 286614
rect 536459 286586 537459 286592
rect 536459 286562 536471 286586
rect 536449 286552 536471 286562
rect 537447 286562 537459 286586
rect 537677 286586 538677 286592
rect 537677 286562 537689 286586
rect 537447 286552 537689 286562
rect 538665 286562 538677 286586
rect 538895 286586 539895 286592
rect 538895 286562 538907 286586
rect 538665 286552 538907 286562
rect 539883 286562 539895 286586
rect 540113 286586 541113 286592
rect 540113 286562 540125 286586
rect 539883 286552 540125 286562
rect 541101 286562 541113 286586
rect 541331 286586 542331 286592
rect 541331 286562 541343 286586
rect 541101 286552 541343 286562
rect 542319 286562 542331 286586
rect 542549 286586 543549 286592
rect 542549 286562 542561 286586
rect 542319 286552 542561 286562
rect 543537 286562 543549 286586
rect 543767 286586 544767 286592
rect 543767 286562 543779 286586
rect 543537 286552 543779 286562
rect 544755 286562 544767 286586
rect 544755 286552 544769 286562
rect 536449 286522 536759 286552
rect 536749 286502 536759 286522
rect 536849 286522 536899 286552
rect 536849 286502 536859 286522
rect 536889 286502 536899 286522
rect 536989 286522 541769 286552
rect 536989 286502 536999 286522
rect 541759 286502 541769 286522
rect 541859 286522 541909 286552
rect 541859 286502 541869 286522
rect 541899 286502 541909 286522
rect 541999 286522 544769 286552
rect 541999 286502 542009 286522
rect 537489 286452 537649 286462
rect 537489 286352 537509 286452
rect 537629 286352 537649 286452
rect 537489 286282 537649 286352
rect 538709 286452 538869 286462
rect 538709 286352 538729 286452
rect 538849 286352 538869 286452
rect 538709 286282 538869 286352
rect 539919 286452 540079 286462
rect 541147 286452 541291 286458
rect 543587 286452 543731 286458
rect 539919 286352 539939 286452
rect 540059 286352 540079 286452
rect 539329 286282 539339 286312
rect 536449 286244 539339 286282
rect 539429 286282 539439 286312
rect 539919 286282 540079 286352
rect 541139 286352 541159 286452
rect 541279 286352 541299 286452
rect 542377 286442 542521 286448
rect 541139 286282 541299 286352
rect 542369 286342 542389 286442
rect 542509 286342 542529 286442
rect 542369 286282 542529 286342
rect 543579 286352 543599 286452
rect 543719 286352 543739 286452
rect 543579 286282 543739 286352
rect 544209 286282 544219 286332
rect 539429 286252 544219 286282
rect 544309 286282 544319 286332
rect 550420 286300 550960 288360
rect 568110 288530 568160 288814
rect 572750 288764 572810 288774
rect 568290 288744 572750 288750
rect 572890 288764 572950 288774
rect 572810 288744 572890 288750
rect 573065 288764 573125 288774
rect 572950 288744 573065 288750
rect 573255 288764 573315 288774
rect 573125 288744 573255 288750
rect 573415 288764 573475 288774
rect 573315 288744 573415 288750
rect 573605 288764 573665 288774
rect 573475 288744 573605 288750
rect 573805 288764 573865 288774
rect 573665 288744 573805 288750
rect 573985 288764 574045 288774
rect 573865 288744 573985 288750
rect 574175 288764 574235 288774
rect 574045 288744 574175 288750
rect 574375 288764 574435 288774
rect 574235 288744 574375 288750
rect 574540 288754 574600 288764
rect 574435 288744 574540 288750
rect 574600 288744 578290 288750
rect 568220 288707 568260 288714
rect 568212 288695 568260 288707
rect 568290 288710 568302 288744
rect 578278 288710 578290 288744
rect 568290 288704 572750 288710
rect 572810 288704 572890 288710
rect 572950 288704 573065 288710
rect 573125 288704 573255 288710
rect 573315 288704 573415 288710
rect 573475 288704 573605 288710
rect 573665 288704 573805 288710
rect 573865 288704 573985 288710
rect 574045 288704 574175 288710
rect 574235 288704 574375 288710
rect 574435 288704 574540 288710
rect 568212 288661 568218 288695
rect 568252 288661 568260 288695
rect 572750 288694 572810 288704
rect 572890 288694 572950 288704
rect 573065 288694 573125 288704
rect 573255 288694 573315 288704
rect 573415 288694 573475 288704
rect 573605 288694 573665 288704
rect 573805 288694 573865 288704
rect 573985 288694 574045 288704
rect 574175 288694 574235 288704
rect 574375 288694 574435 288704
rect 574600 288704 578290 288710
rect 574540 288684 574600 288694
rect 568212 288654 568260 288661
rect 578320 288654 578660 288660
rect 568212 288652 568310 288654
rect 578280 288652 578660 288654
rect 568212 288649 578660 288652
rect 568110 287944 568116 288530
rect 568150 287944 568160 288530
rect 568220 288646 578660 288649
rect 568220 288612 568302 288646
rect 578278 288612 578660 288646
rect 568220 288606 578660 288612
rect 568220 288604 568310 288606
rect 578280 288604 578660 288606
rect 568220 288511 568260 288604
rect 578320 288600 578660 288604
rect 578320 288597 578360 288600
rect 572750 288564 572810 288574
rect 568212 288499 568260 288511
rect 568290 288548 572750 288554
rect 572890 288564 572950 288574
rect 572810 288548 572890 288554
rect 573065 288564 573125 288574
rect 572950 288548 573065 288554
rect 573255 288564 573315 288574
rect 573125 288548 573255 288554
rect 573415 288564 573475 288574
rect 573315 288548 573415 288554
rect 573605 288564 573665 288574
rect 573475 288548 573605 288554
rect 573805 288564 573865 288574
rect 573665 288548 573805 288554
rect 573985 288564 574045 288574
rect 573865 288548 573985 288554
rect 574175 288564 574235 288574
rect 574045 288548 574175 288554
rect 574375 288564 574435 288574
rect 574235 288548 574375 288554
rect 574540 288564 574600 288574
rect 574435 288548 574540 288554
rect 578320 288563 578328 288597
rect 574600 288548 578290 288554
rect 568290 288514 568302 288548
rect 578278 288514 578290 288548
rect 568290 288508 572750 288514
rect 568212 288465 568218 288499
rect 568252 288465 568260 288499
rect 572810 288508 572890 288514
rect 572750 288494 572810 288504
rect 572950 288508 573065 288514
rect 572890 288494 572950 288504
rect 573125 288508 573255 288514
rect 573065 288494 573125 288504
rect 573315 288508 573415 288514
rect 573255 288494 573315 288504
rect 573475 288508 573605 288514
rect 573415 288494 573475 288504
rect 573665 288508 573805 288514
rect 573605 288494 573665 288504
rect 573865 288508 573985 288514
rect 573805 288494 573865 288504
rect 574045 288508 574175 288514
rect 573985 288494 574045 288504
rect 574235 288508 574375 288514
rect 574175 288494 574235 288504
rect 574435 288508 574540 288514
rect 574375 288494 574435 288504
rect 574600 288508 578290 288514
rect 578320 288520 578360 288563
rect 578440 288520 578540 288600
rect 578620 288520 578660 288600
rect 574540 288494 574600 288504
rect 568212 288464 568260 288465
rect 568212 288456 568310 288464
rect 568212 288454 578290 288456
rect 578320 288454 578660 288520
rect 568212 288453 578660 288454
rect 568220 288450 578660 288453
rect 568220 288416 568302 288450
rect 578278 288440 578660 288450
rect 578278 288416 578360 288440
rect 568220 288410 578360 288416
rect 568220 288404 568310 288410
rect 578280 288404 578360 288410
rect 568220 288315 568260 288404
rect 578320 288401 578360 288404
rect 572750 288364 572810 288374
rect 568212 288303 568260 288315
rect 568290 288352 572750 288358
rect 572890 288364 572950 288374
rect 572810 288352 572890 288358
rect 573065 288364 573125 288374
rect 572950 288352 573065 288358
rect 573255 288364 573315 288374
rect 573125 288352 573255 288358
rect 573415 288364 573475 288374
rect 573315 288352 573415 288358
rect 573605 288364 573665 288374
rect 573475 288352 573605 288358
rect 573805 288364 573865 288374
rect 573665 288352 573805 288358
rect 573985 288364 574045 288374
rect 573865 288352 573985 288358
rect 574175 288364 574235 288374
rect 574045 288352 574175 288358
rect 574375 288364 574435 288374
rect 574235 288352 574375 288358
rect 574540 288364 574600 288374
rect 574435 288352 574540 288358
rect 578320 288367 578328 288401
rect 578320 288360 578360 288367
rect 578440 288360 578540 288440
rect 578620 288360 578660 288440
rect 574600 288352 578290 288358
rect 568290 288318 568302 288352
rect 578278 288318 578290 288352
rect 568290 288312 572750 288318
rect 568212 288269 568218 288303
rect 568252 288269 568260 288303
rect 572810 288312 572890 288318
rect 572750 288294 572810 288304
rect 572950 288312 573065 288318
rect 572890 288294 572950 288304
rect 573125 288312 573255 288318
rect 573065 288294 573125 288304
rect 573315 288312 573415 288318
rect 573255 288294 573315 288304
rect 573475 288312 573605 288318
rect 573415 288294 573475 288304
rect 573665 288312 573805 288318
rect 573605 288294 573665 288304
rect 573865 288312 573985 288318
rect 573805 288294 573865 288304
rect 574045 288312 574175 288318
rect 573985 288294 574045 288304
rect 574235 288312 574375 288318
rect 574175 288294 574235 288304
rect 574435 288312 574540 288318
rect 574375 288294 574435 288304
rect 574600 288312 578290 288318
rect 574540 288294 574600 288304
rect 568212 288264 568260 288269
rect 578320 288280 578660 288360
rect 578320 288264 578360 288280
rect 568212 288260 568310 288264
rect 578280 288260 578360 288264
rect 568212 288257 578360 288260
rect 568220 288254 578360 288257
rect 568220 288220 568302 288254
rect 578278 288220 578360 288254
rect 568220 288214 578360 288220
rect 568220 288204 568310 288214
rect 578320 288205 578360 288214
rect 568220 288119 568260 288204
rect 572750 288174 572810 288184
rect 568212 288107 568260 288119
rect 568290 288156 572750 288162
rect 572890 288174 572950 288184
rect 572810 288156 572890 288162
rect 573065 288174 573125 288184
rect 572950 288156 573065 288162
rect 573255 288174 573315 288184
rect 573125 288156 573255 288162
rect 573415 288174 573475 288184
rect 573315 288156 573415 288162
rect 573605 288174 573665 288184
rect 573475 288156 573605 288162
rect 573805 288174 573865 288184
rect 573665 288156 573805 288162
rect 573985 288174 574045 288184
rect 573865 288156 573985 288162
rect 574175 288174 574235 288184
rect 574045 288156 574175 288162
rect 574375 288174 574435 288184
rect 574235 288156 574375 288162
rect 574540 288174 574600 288184
rect 574435 288156 574540 288162
rect 578320 288171 578328 288205
rect 578440 288200 578540 288280
rect 578620 288200 578660 288280
rect 578362 288171 578660 288200
rect 574600 288156 578290 288162
rect 568290 288122 568302 288156
rect 578278 288122 578290 288156
rect 568290 288116 572750 288122
rect 568212 288073 568218 288107
rect 568252 288074 568260 288107
rect 572810 288116 572890 288122
rect 572750 288104 572810 288114
rect 572950 288116 573065 288122
rect 572890 288104 572950 288114
rect 573125 288116 573255 288122
rect 573065 288104 573125 288114
rect 573315 288116 573415 288122
rect 573255 288104 573315 288114
rect 573475 288116 573605 288122
rect 573415 288104 573475 288114
rect 573665 288116 573805 288122
rect 573605 288104 573665 288114
rect 573865 288116 573985 288122
rect 573805 288104 573865 288114
rect 574045 288116 574175 288122
rect 573985 288104 574045 288114
rect 574235 288116 574375 288122
rect 574175 288104 574235 288114
rect 574435 288116 574540 288122
rect 574375 288104 574435 288114
rect 574600 288116 578290 288122
rect 574540 288104 574600 288114
rect 578320 288100 578660 288171
rect 568252 288073 568310 288074
rect 568212 288064 568310 288073
rect 578320 288064 578360 288100
rect 568212 288061 578360 288064
rect 568110 287654 568160 287944
rect 568220 288058 578360 288061
rect 568220 288024 568302 288058
rect 578278 288024 578360 288058
rect 568220 288020 578360 288024
rect 578440 288020 578540 288100
rect 578620 288020 578660 288100
rect 568220 288018 578660 288020
rect 568220 288014 568310 288018
rect 578280 288014 578660 288018
rect 568220 287923 568260 288014
rect 578320 288009 578660 288014
rect 572750 287974 572810 287984
rect 568212 287911 568260 287923
rect 568290 287960 572750 287966
rect 572890 287974 572950 287984
rect 572810 287960 572890 287966
rect 573065 287974 573125 287984
rect 572950 287960 573065 287966
rect 573255 287974 573315 287984
rect 573125 287960 573255 287966
rect 573415 287974 573475 287984
rect 573315 287960 573415 287966
rect 573605 287974 573665 287984
rect 573475 287960 573605 287966
rect 573805 287974 573865 287984
rect 573665 287960 573805 287966
rect 573985 287974 574045 287984
rect 573865 287960 573985 287966
rect 574175 287974 574235 287984
rect 574045 287960 574175 287966
rect 574375 287974 574435 287984
rect 574235 287960 574375 287966
rect 574540 287974 574600 287984
rect 574435 287960 574540 287966
rect 578320 287975 578328 288009
rect 578362 287975 578660 288009
rect 574600 287960 578290 287966
rect 568290 287926 568302 287960
rect 578278 287926 578290 287960
rect 568290 287920 572750 287926
rect 568212 287877 568218 287911
rect 568252 287877 568260 287911
rect 572810 287920 572890 287926
rect 572750 287904 572810 287914
rect 572950 287920 573065 287926
rect 572890 287904 572950 287914
rect 573125 287920 573255 287926
rect 573065 287904 573125 287914
rect 573315 287920 573415 287926
rect 573255 287904 573315 287914
rect 573475 287920 573605 287926
rect 573415 287904 573475 287914
rect 573665 287920 573805 287926
rect 573605 287904 573665 287914
rect 573865 287920 573985 287926
rect 573805 287904 573865 287914
rect 574045 287920 574175 287926
rect 573985 287904 574045 287914
rect 574235 287920 574375 287926
rect 574175 287904 574235 287914
rect 574435 287920 574540 287926
rect 574375 287904 574435 287914
rect 574600 287920 578290 287926
rect 578320 287940 578660 287975
rect 574540 287904 574600 287914
rect 568212 287874 568260 287877
rect 578320 287874 578360 287940
rect 568212 287868 568310 287874
rect 578280 287868 578360 287874
rect 568212 287865 578360 287868
rect 568220 287862 578360 287865
rect 568220 287828 568302 287862
rect 578278 287860 578360 287862
rect 578440 287860 578540 287940
rect 578620 287860 578660 287940
rect 578278 287828 578660 287860
rect 568220 287824 578660 287828
rect 568220 287822 578290 287824
rect 568220 287814 568310 287822
rect 578320 287813 578660 287824
rect 572750 287774 572810 287784
rect 568290 287764 572750 287770
rect 572890 287774 572950 287784
rect 572810 287764 572890 287770
rect 573065 287774 573125 287784
rect 572950 287764 573065 287770
rect 573255 287774 573315 287784
rect 573125 287764 573255 287770
rect 573415 287774 573475 287784
rect 573315 287764 573415 287770
rect 573605 287774 573665 287784
rect 573475 287764 573605 287770
rect 573805 287774 573865 287784
rect 573665 287764 573805 287770
rect 573985 287774 574045 287784
rect 573865 287764 573985 287770
rect 574175 287774 574235 287784
rect 574045 287764 574175 287770
rect 574375 287774 574435 287784
rect 574235 287764 574375 287770
rect 574540 287774 574600 287784
rect 574435 287764 574540 287770
rect 578320 287779 578328 287813
rect 578362 287779 578660 287813
rect 574600 287764 578290 287770
rect 568290 287730 568302 287764
rect 578278 287730 578290 287764
rect 578320 287740 578660 287779
rect 568290 287724 572750 287730
rect 572810 287724 572890 287730
rect 572750 287704 572810 287714
rect 572950 287724 573065 287730
rect 572890 287704 572950 287714
rect 573125 287724 573255 287730
rect 573065 287704 573125 287714
rect 573315 287724 573415 287730
rect 573255 287704 573315 287714
rect 573475 287724 573605 287730
rect 573415 287704 573475 287714
rect 573665 287724 573805 287730
rect 573605 287704 573665 287714
rect 573865 287724 573985 287730
rect 573805 287704 573865 287714
rect 574045 287724 574175 287730
rect 573985 287704 574045 287714
rect 574235 287724 574375 287730
rect 574175 287704 574235 287714
rect 574435 287724 574540 287730
rect 574375 287704 574435 287714
rect 574600 287724 578290 287730
rect 574540 287704 574600 287714
rect 570708 287654 575872 287656
rect 568110 287650 578380 287654
rect 567800 287616 570720 287650
rect 575860 287616 578380 287650
rect 567800 287604 578380 287616
rect 544309 286252 544769 286282
rect 539429 286244 544769 286252
rect 536449 286242 536471 286244
rect 536459 286210 536471 286242
rect 537447 286242 537689 286244
rect 537447 286210 537459 286242
rect 536459 286204 537459 286210
rect 537677 286210 537689 286242
rect 538665 286242 538907 286244
rect 538665 286210 538677 286242
rect 537677 286204 538677 286210
rect 538895 286210 538907 286242
rect 539883 286242 540125 286244
rect 539883 286210 539895 286242
rect 538895 286204 539895 286210
rect 540113 286210 540125 286242
rect 541101 286242 541343 286244
rect 541101 286210 541113 286242
rect 540113 286204 541113 286210
rect 541331 286210 541343 286242
rect 542319 286242 542561 286244
rect 542319 286210 542331 286242
rect 541331 286204 542331 286210
rect 542549 286210 542561 286242
rect 543537 286242 543779 286244
rect 543537 286210 543549 286242
rect 542549 286204 543549 286210
rect 543767 286210 543779 286242
rect 544755 286242 544769 286244
rect 544755 286210 544767 286242
rect 543767 286204 544767 286210
rect 550420 286200 559740 286300
rect 536381 286182 536427 286194
rect 536381 286014 536387 286182
rect 536421 286162 536427 286182
rect 537491 286182 537537 286194
rect 537491 286162 537497 286182
rect 536421 286042 537497 286162
rect 536421 286014 536427 286042
rect 536381 286002 536427 286014
rect 537491 286014 537497 286042
rect 537531 286162 537537 286182
rect 537599 286182 537645 286194
rect 537599 286162 537605 286182
rect 537531 286042 537605 286162
rect 537531 286014 537537 286042
rect 537491 286002 537537 286014
rect 537599 286014 537605 286042
rect 537639 286162 537645 286182
rect 538709 286182 538755 286194
rect 538709 286162 538715 286182
rect 537639 286142 538715 286162
rect 537639 286062 538109 286142
rect 538199 286062 538229 286142
rect 538319 286062 538715 286142
rect 537639 286042 538715 286062
rect 537639 286014 537645 286042
rect 537599 286002 537645 286014
rect 538709 286014 538715 286042
rect 538749 286162 538755 286182
rect 538817 286182 538863 286194
rect 538817 286162 538823 286182
rect 538749 286042 538823 286162
rect 538749 286014 538755 286042
rect 538709 286002 538755 286014
rect 538817 286014 538823 286042
rect 538857 286162 538863 286182
rect 539927 286182 539973 286194
rect 539927 286162 539933 286182
rect 538857 286042 539933 286162
rect 538857 286014 538863 286042
rect 538817 286002 538863 286014
rect 539927 286014 539933 286042
rect 539967 286162 539973 286182
rect 540035 286182 540081 286194
rect 540035 286162 540041 286182
rect 539967 286042 540041 286162
rect 539967 286014 539973 286042
rect 539927 286002 539973 286014
rect 540035 286014 540041 286042
rect 540075 286162 540081 286182
rect 541145 286182 541191 286194
rect 541145 286162 541151 286182
rect 540075 286146 541151 286162
rect 540075 286056 540420 286146
rect 540508 286142 541151 286146
rect 540508 286062 540559 286142
rect 540649 286062 540679 286142
rect 540769 286062 541151 286142
rect 540508 286056 541151 286062
rect 540075 286042 541151 286056
rect 540075 286014 540081 286042
rect 540035 286002 540081 286014
rect 541145 286014 541151 286042
rect 541185 286162 541191 286182
rect 541253 286182 541299 286194
rect 541253 286162 541259 286182
rect 541185 286042 541259 286162
rect 541185 286014 541191 286042
rect 541145 286002 541191 286014
rect 541253 286014 541259 286042
rect 541293 286162 541299 286182
rect 542363 286182 542409 286194
rect 542363 286162 542369 286182
rect 541293 286042 542369 286162
rect 541293 286014 541299 286042
rect 541253 286002 541299 286014
rect 542363 286014 542369 286042
rect 542403 286162 542409 286182
rect 542471 286182 542517 286194
rect 542471 286162 542477 286182
rect 542403 286042 542477 286162
rect 542403 286014 542409 286042
rect 542363 286002 542409 286014
rect 542471 286014 542477 286042
rect 542511 286162 542517 286182
rect 543581 286182 543627 286194
rect 543581 286162 543587 286182
rect 542511 286142 543587 286162
rect 542511 286062 542989 286142
rect 543079 286062 543109 286142
rect 543199 286062 543587 286142
rect 542511 286042 543587 286062
rect 542511 286014 542517 286042
rect 542471 286002 542517 286014
rect 543581 286014 543587 286042
rect 543621 286162 543627 286182
rect 543689 286182 543735 286194
rect 543689 286162 543695 286182
rect 543621 286042 543695 286162
rect 543621 286014 543627 286042
rect 543581 286002 543627 286014
rect 543689 286014 543695 286042
rect 543729 286162 543735 286182
rect 544799 286182 544845 286194
rect 544799 286162 544805 286182
rect 543729 286042 544805 286162
rect 543729 286014 543735 286042
rect 543689 286002 543735 286014
rect 544799 286014 544805 286042
rect 544839 286162 544845 286182
rect 544839 286042 544849 286162
rect 544839 286014 544845 286042
rect 544799 286002 544845 286014
rect 550420 286000 557700 286200
rect 557900 286000 558100 286200
rect 558300 286000 558500 286200
rect 558700 286000 558900 286200
rect 559100 286000 559300 286200
rect 559500 286000 559740 286200
rect 536459 285986 537459 285992
rect 536459 285962 536471 285986
rect 537447 285962 537459 285986
rect 537677 285986 538677 285992
rect 537677 285962 537689 285986
rect 536449 285952 536471 285962
rect 537447 285952 537689 285962
rect 538665 285962 538677 285986
rect 538895 285986 539895 285992
rect 538895 285962 538907 285986
rect 538665 285952 538907 285962
rect 539883 285962 539895 285986
rect 540113 285986 541113 285992
rect 540113 285962 540125 285986
rect 539883 285952 540125 285962
rect 541101 285962 541113 285986
rect 541331 285986 542331 285992
rect 541331 285962 541343 285986
rect 541101 285952 541343 285962
rect 542319 285962 542331 285986
rect 542549 285986 543549 285992
rect 542549 285962 542561 285986
rect 542319 285952 542561 285962
rect 543537 285962 543549 285986
rect 543767 285986 544767 285992
rect 543767 285962 543779 285986
rect 543537 285952 543779 285962
rect 544755 285962 544767 285986
rect 544755 285952 544769 285962
rect 536449 285922 536759 285952
rect 536749 285882 536759 285922
rect 536849 285922 536899 285952
rect 536849 285882 536859 285922
rect 536889 285882 536899 285922
rect 536989 285922 541769 285952
rect 536989 285882 536999 285922
rect 541759 285902 541769 285922
rect 541859 285922 541909 285952
rect 541859 285902 541869 285922
rect 541899 285902 541909 285922
rect 541999 285922 544769 285952
rect 541999 285902 542009 285922
rect 550420 285800 559740 286000
rect 550420 285600 557700 285800
rect 557900 285600 558100 285800
rect 558300 285600 558500 285800
rect 558700 285600 558900 285800
rect 559100 285600 559300 285800
rect 559500 285600 559740 285800
rect 537372 285478 537556 285484
rect 538432 285478 538616 285484
rect 539892 285478 540076 285484
rect 541112 285478 541296 285484
rect 542592 285478 542776 285484
rect 543592 285478 543776 285484
rect 537004 285318 537384 285478
rect 537544 285318 538444 285478
rect 538604 285318 539904 285478
rect 540064 285318 541124 285478
rect 541284 285318 542604 285478
rect 542764 285318 543604 285478
rect 543764 285318 544204 285478
rect 537004 285270 544204 285318
rect 537004 285236 537025 285270
rect 538001 285258 538261 285270
rect 538001 285236 538024 285258
rect 536926 285208 536972 285220
rect 537004 285218 538024 285236
rect 538244 285236 538261 285258
rect 539237 285258 539497 285270
rect 539237 285236 539249 285258
rect 538244 285230 539249 285236
rect 539484 285236 539497 285258
rect 540473 285258 540733 285270
rect 540473 285236 540485 285258
rect 539484 285230 540485 285236
rect 540721 285236 540733 285258
rect 541709 285258 541969 285270
rect 541709 285236 541724 285258
rect 540721 285230 541724 285236
rect 536926 285040 536932 285208
rect 536966 285168 536972 285208
rect 538054 285208 538100 285220
rect 538054 285168 538060 285208
rect 536966 285040 538060 285168
rect 538094 285168 538100 285208
rect 538162 285208 538208 285220
rect 538244 285218 539244 285230
rect 538162 285168 538168 285208
rect 538094 285040 538168 285168
rect 538202 285168 538208 285208
rect 539290 285208 539336 285220
rect 539290 285168 539296 285208
rect 538202 285158 539296 285168
rect 538202 285088 538884 285158
rect 538954 285088 539104 285158
rect 539174 285088 539296 285158
rect 538202 285040 539296 285088
rect 539330 285168 539336 285208
rect 539398 285208 539444 285220
rect 539484 285218 540484 285230
rect 539398 285168 539404 285208
rect 539330 285040 539404 285168
rect 539438 285168 539444 285208
rect 540526 285208 540572 285220
rect 540526 285168 540532 285208
rect 539438 285040 540532 285168
rect 540566 285168 540572 285208
rect 540634 285208 540680 285220
rect 540724 285218 541724 285230
rect 541944 285236 541969 285258
rect 542945 285258 543205 285270
rect 542945 285236 542964 285258
rect 540634 285168 540640 285208
rect 540566 285040 540640 285168
rect 540674 285168 540680 285208
rect 541762 285208 541808 285220
rect 541762 285168 541768 285208
rect 540674 285040 541768 285168
rect 541802 285168 541808 285208
rect 541870 285208 541916 285220
rect 541944 285218 542964 285236
rect 543184 285236 543205 285258
rect 544181 285236 544204 285270
rect 541870 285168 541876 285208
rect 541802 285040 541876 285168
rect 541910 285168 541916 285208
rect 542998 285208 543044 285220
rect 542998 285168 543004 285208
rect 541910 285158 543004 285168
rect 541910 285088 542064 285158
rect 542134 285088 542304 285158
rect 542374 285088 543004 285158
rect 541910 285040 543004 285088
rect 543038 285168 543044 285208
rect 543106 285208 543152 285220
rect 543184 285218 544204 285236
rect 550420 285400 559740 285600
rect 543106 285168 543112 285208
rect 543038 285040 543112 285168
rect 543146 285168 543152 285208
rect 544234 285208 544280 285220
rect 544234 285168 544240 285208
rect 543146 285040 544240 285168
rect 544274 285040 544280 285208
rect 536926 285028 544280 285040
rect 550420 285200 557700 285400
rect 557900 285200 558100 285400
rect 558300 285200 558500 285400
rect 558700 285200 558900 285400
rect 559100 285200 559300 285400
rect 559500 285200 559740 285400
rect 536926 285012 544274 285028
rect 536926 284978 537025 285012
rect 538001 284978 538261 285012
rect 539237 284978 539497 285012
rect 540473 284978 540733 285012
rect 541709 284978 541969 285012
rect 542945 284978 543205 285012
rect 544181 284978 544274 285012
rect 536926 284956 544274 284978
rect 550420 285000 559740 285200
rect 537372 284898 537556 284904
rect 538432 284898 538616 284904
rect 539892 284898 540076 284904
rect 541112 284898 541296 284904
rect 542592 284898 542776 284904
rect 543592 284898 543776 284904
rect 537004 284738 537384 284898
rect 537544 284738 538444 284898
rect 538604 284738 539904 284898
rect 540064 284738 541124 284898
rect 541284 284738 542604 284898
rect 542764 284738 543604 284898
rect 543764 284738 544204 284898
rect 537004 284680 544204 284738
rect 537004 284658 537025 284680
rect 537013 284646 537025 284658
rect 538001 284668 538261 284680
rect 538001 284646 538013 284668
rect 537013 284640 538013 284646
rect 538249 284646 538261 284668
rect 539237 284668 539497 284680
rect 539237 284646 539249 284668
rect 538249 284640 539249 284646
rect 539485 284646 539497 284668
rect 540473 284668 540733 284680
rect 540473 284646 540485 284668
rect 539485 284640 540485 284646
rect 540721 284646 540733 284668
rect 541709 284668 541969 284680
rect 541709 284646 541721 284668
rect 540721 284640 541721 284646
rect 541957 284646 541969 284668
rect 542945 284668 543205 284680
rect 542945 284646 542957 284668
rect 541957 284640 542957 284646
rect 543193 284646 543205 284668
rect 544181 284658 544204 284680
rect 550420 284800 557700 285000
rect 557900 284800 558100 285000
rect 558300 284800 558500 285000
rect 558700 284800 558900 285000
rect 559100 284800 559300 285000
rect 559500 284800 559740 285000
rect 544181 284646 544193 284658
rect 543193 284640 544193 284646
rect 536926 284618 536972 284630
rect 536926 284578 536932 284618
rect 536924 284488 536932 284578
rect 536926 284450 536932 284488
rect 536966 284578 536972 284618
rect 538054 284618 538100 284630
rect 538054 284578 538060 284618
rect 536966 284488 538060 284578
rect 536966 284450 536972 284488
rect 536926 284438 536972 284450
rect 538054 284450 538060 284488
rect 538094 284578 538100 284618
rect 538162 284618 538208 284630
rect 538162 284578 538168 284618
rect 538094 284488 538168 284578
rect 538094 284450 538100 284488
rect 538054 284438 538100 284450
rect 538162 284450 538168 284488
rect 538202 284578 538208 284618
rect 539290 284618 539336 284630
rect 539290 284578 539296 284618
rect 538202 284568 539296 284578
rect 538202 284498 538884 284568
rect 538954 284498 539104 284568
rect 539174 284498 539296 284568
rect 538202 284488 539296 284498
rect 538202 284450 538208 284488
rect 538162 284438 538208 284450
rect 539290 284450 539296 284488
rect 539330 284578 539336 284618
rect 539398 284618 539444 284630
rect 539398 284578 539404 284618
rect 539330 284488 539404 284578
rect 539330 284450 539336 284488
rect 539290 284438 539336 284450
rect 539398 284450 539404 284488
rect 539438 284578 539444 284618
rect 540526 284618 540572 284630
rect 540526 284578 540532 284618
rect 539438 284488 540532 284578
rect 539438 284450 539444 284488
rect 539398 284438 539444 284450
rect 540526 284450 540532 284488
rect 540566 284578 540572 284618
rect 540634 284618 540680 284630
rect 540634 284578 540640 284618
rect 540566 284488 540640 284578
rect 540566 284450 540572 284488
rect 540526 284438 540572 284450
rect 540634 284450 540640 284488
rect 540674 284578 540680 284618
rect 541762 284618 541808 284630
rect 541762 284578 541768 284618
rect 540674 284488 541768 284578
rect 540674 284450 540680 284488
rect 540634 284438 540680 284450
rect 541762 284450 541768 284488
rect 541802 284578 541808 284618
rect 541870 284618 541916 284630
rect 541870 284578 541876 284618
rect 541802 284488 541876 284578
rect 541802 284450 541808 284488
rect 541762 284438 541808 284450
rect 541870 284450 541876 284488
rect 541910 284578 541916 284618
rect 542998 284618 543044 284630
rect 542998 284578 543004 284618
rect 541910 284568 543004 284578
rect 541910 284498 542064 284568
rect 542134 284498 542304 284568
rect 542374 284498 543004 284568
rect 541910 284488 543004 284498
rect 541910 284450 541916 284488
rect 541870 284438 541916 284450
rect 542998 284450 543004 284488
rect 543038 284578 543044 284618
rect 543106 284618 543152 284630
rect 543106 284578 543112 284618
rect 543038 284488 543112 284578
rect 543038 284450 543044 284488
rect 542998 284438 543044 284450
rect 543106 284450 543112 284488
rect 543146 284578 543152 284618
rect 544234 284618 544280 284630
rect 544234 284578 544240 284618
rect 543146 284488 544240 284578
rect 543146 284450 543152 284488
rect 543106 284438 543152 284450
rect 544234 284450 544240 284488
rect 544274 284450 544280 284618
rect 544234 284438 544280 284450
rect 550420 284600 559740 284800
rect 537004 284422 538013 284428
rect 537004 284388 537025 284422
rect 538001 284408 538013 284422
rect 538249 284422 539249 284428
rect 538249 284408 538261 284422
rect 538001 284388 538261 284408
rect 539237 284408 539249 284422
rect 539485 284422 540485 284428
rect 539485 284408 539497 284422
rect 540473 284408 540485 284422
rect 540721 284422 541721 284428
rect 540721 284408 540733 284422
rect 541709 284408 541721 284422
rect 541957 284422 542957 284428
rect 541957 284408 541969 284422
rect 539237 284388 539497 284408
rect 540473 284388 540733 284408
rect 541709 284388 541969 284408
rect 542945 284408 542957 284422
rect 543193 284422 544198 284428
rect 543193 284408 543205 284422
rect 542945 284388 543205 284408
rect 544181 284388 544198 284422
rect 537004 284338 540044 284388
rect 540114 284338 540154 284388
rect 540224 284338 540984 284388
rect 541054 284338 541094 284388
rect 541164 284338 544198 284388
rect 537004 284328 544198 284338
rect 550420 284400 557700 284600
rect 557900 284400 558100 284600
rect 558300 284400 558500 284600
rect 558700 284400 558900 284600
rect 559100 284400 559300 284600
rect 559500 284400 559740 284600
rect 550420 284200 559740 284400
rect 550420 284000 557700 284200
rect 557900 284000 558100 284200
rect 558300 284000 558500 284200
rect 558700 284000 558900 284200
rect 559100 284000 559300 284200
rect 559500 284000 559740 284200
rect 540400 283918 540410 283926
rect 539684 283890 540410 283918
rect 540470 283890 540510 283926
rect 539684 283856 539786 283890
rect 540012 283856 540254 283890
rect 540480 283866 540510 283890
rect 540570 283866 540610 283926
rect 540670 283866 540710 283926
rect 540770 283918 540780 283926
rect 540770 283890 541504 283918
rect 540480 283856 540722 283866
rect 540948 283856 541190 283890
rect 541416 283856 541504 283890
rect 539684 283848 541504 283856
rect 539684 283838 540984 283848
rect 539684 283828 540044 283838
rect 539684 283768 539702 283828
rect 539696 283660 539702 283768
rect 539736 283768 540044 283828
rect 540114 283768 540154 283838
rect 540224 283828 540984 283838
rect 540224 283768 540530 283828
rect 539736 283688 540062 283768
rect 539736 283660 539742 283688
rect 539696 283648 539742 283660
rect 540054 283660 540062 283688
rect 540096 283660 540170 283768
rect 540204 283688 540530 283768
rect 540204 283660 540214 283688
rect 540054 283648 540214 283660
rect 540524 283660 540530 283688
rect 540564 283660 540638 283828
rect 540672 283778 540984 283828
rect 541054 283778 541094 283848
rect 541164 283840 541504 283848
rect 541164 283828 541506 283840
rect 541164 283778 541466 283828
rect 540672 283688 540998 283778
rect 540672 283660 540679 283688
rect 540524 283648 540679 283660
rect 540992 283660 540998 283688
rect 541032 283660 541106 283778
rect 541140 283688 541466 283778
rect 541140 283660 541149 283688
rect 540992 283648 541149 283660
rect 541460 283660 541466 283688
rect 541500 283660 541506 283828
rect 541460 283648 541506 283660
rect 550420 283800 559740 284000
rect 539774 283632 540024 283638
rect 539774 283618 539786 283632
rect 539764 283598 539786 283618
rect 540012 283618 540024 283632
rect 540242 283632 540492 283638
rect 540242 283618 540254 283632
rect 540012 283598 540254 283618
rect 540480 283618 540492 283632
rect 540710 283632 540960 283638
rect 540710 283618 540722 283632
rect 540480 283598 540722 283618
rect 540948 283618 540960 283632
rect 541178 283632 541428 283638
rect 541178 283618 541190 283632
rect 540948 283598 541190 283618
rect 541416 283618 541428 283632
rect 541416 283598 541434 283618
rect 539764 283578 541434 283598
rect 550420 283600 557700 283800
rect 557900 283600 558100 283800
rect 558300 283600 558500 283800
rect 558700 283600 558900 283800
rect 559100 283600 559300 283800
rect 559500 283600 559740 283800
rect 539764 283524 541474 283578
rect 539752 283518 541486 283524
rect 539752 283368 539764 283518
rect 539984 283508 540284 283518
rect 539984 283368 539996 283508
rect 539752 283362 539996 283368
rect 540272 283368 540284 283508
rect 540504 283508 540704 283518
rect 540504 283368 540516 283508
rect 540272 283362 540516 283368
rect 540692 283368 540704 283508
rect 540924 283508 541254 283518
rect 540924 283368 540936 283508
rect 540692 283362 540936 283368
rect 541242 283368 541254 283508
rect 541474 283368 541486 283518
rect 541242 283362 541486 283368
rect 550420 283400 559740 283600
rect 542044 283328 542394 283348
rect 538864 283308 542064 283328
rect 538864 283238 538884 283308
rect 538954 283238 539094 283308
rect 539164 283265 542064 283308
rect 539164 283238 540006 283265
rect 538864 283231 540006 283238
rect 540482 283231 540724 283265
rect 541200 283258 542064 283265
rect 542134 283258 542304 283328
rect 542374 283258 542394 283328
rect 541200 283238 542394 283258
rect 541200 283231 542064 283238
rect 538864 283218 542064 283231
rect 538864 283148 538884 283218
rect 538954 283148 539094 283218
rect 539164 283203 542064 283218
rect 539164 283148 539922 283203
rect 538864 283118 539194 283148
rect 539916 283135 539922 283148
rect 539956 283148 540532 283203
rect 539956 283135 539962 283148
rect 539916 283123 539962 283135
rect 540526 283135 540532 283148
rect 540566 283148 540640 283203
rect 540566 283135 540572 283148
rect 540526 283123 540572 283135
rect 540634 283135 540640 283148
rect 540674 283148 541250 283203
rect 540674 283135 540680 283148
rect 540634 283123 540680 283135
rect 541244 283135 541250 283148
rect 541284 283168 542064 283203
rect 542134 283168 542304 283238
rect 542374 283168 542394 283238
rect 541284 283148 542394 283168
rect 550420 283200 557700 283400
rect 557900 283200 558100 283400
rect 558300 283200 558500 283400
rect 558700 283200 558900 283400
rect 559100 283200 559300 283400
rect 559500 283200 559740 283400
rect 541284 283135 541290 283148
rect 541244 283123 541290 283135
rect 539994 283107 540494 283113
rect 539994 283093 540006 283107
rect 539989 283078 540006 283093
rect 540482 283093 540494 283107
rect 540712 283107 541212 283113
rect 540712 283093 540724 283107
rect 539984 283073 540006 283078
rect 540482 283073 540724 283093
rect 541200 283093 541212 283107
rect 541200 283078 541224 283093
rect 541200 283073 541234 283078
rect 539984 283018 540044 283073
rect 540114 283018 540154 283073
rect 540224 283018 540984 283073
rect 541054 283018 541094 283073
rect 541164 283018 541234 283073
rect 539984 283008 541234 283018
rect 550420 283000 559740 283200
rect 539512 282968 539716 282974
rect 537392 282958 537596 282964
rect 537392 282828 537404 282958
rect 537584 282828 537596 282958
rect 537392 282822 537596 282828
rect 538532 282958 538736 282964
rect 538532 282828 538544 282958
rect 538724 282828 538736 282958
rect 539512 282838 539524 282968
rect 539704 282838 539716 282968
rect 539512 282832 539716 282838
rect 540282 282968 540486 282974
rect 540282 282838 540294 282968
rect 540474 282838 540486 282968
rect 540282 282832 540486 282838
rect 540722 282968 540926 282974
rect 540722 282838 540734 282968
rect 540914 282838 540926 282968
rect 542512 282968 542716 282974
rect 540722 282832 540926 282838
rect 541442 282958 541646 282964
rect 538532 282822 538736 282828
rect 541442 282828 541454 282958
rect 541634 282828 541646 282958
rect 542512 282838 542524 282968
rect 542704 282838 542716 282968
rect 542512 282832 542716 282838
rect 543512 282968 543716 282974
rect 543512 282838 543524 282968
rect 543704 282838 543716 282968
rect 543512 282832 543716 282838
rect 541442 282822 541646 282828
rect 550420 282800 557700 283000
rect 557900 282800 558100 283000
rect 558300 282800 558500 283000
rect 558700 282800 558900 283000
rect 559100 282800 559300 283000
rect 559500 282800 559740 283000
rect 537054 282788 544144 282793
rect 537054 282740 538884 282788
rect 538954 282740 539104 282788
rect 539174 282740 542064 282788
rect 542134 282740 542304 282788
rect 542374 282746 544144 282788
rect 542374 282740 544149 282746
rect 537054 282718 537071 282740
rect 537059 282706 537071 282718
rect 538047 282718 538289 282740
rect 539265 282718 539507 282740
rect 538047 282706 538059 282718
rect 537059 282700 538059 282706
rect 538277 282706 538289 282718
rect 539265 282706 539277 282718
rect 538277 282700 539277 282706
rect 539495 282706 539507 282718
rect 540483 282718 540725 282740
rect 540483 282706 540495 282718
rect 539495 282700 540495 282706
rect 540713 282706 540725 282718
rect 541701 282718 541943 282740
rect 542919 282718 543161 282740
rect 541701 282706 541713 282718
rect 540713 282700 541713 282706
rect 541931 282706 541943 282718
rect 542919 282706 542931 282718
rect 541931 282700 542931 282706
rect 543149 282706 543161 282718
rect 544137 282706 544149 282740
rect 543149 282700 544149 282706
rect 536981 282678 537027 282690
rect 536981 282510 536987 282678
rect 537021 282643 537027 282678
rect 538091 282678 538137 282690
rect 538091 282643 538097 282678
rect 537021 282558 538097 282643
rect 537021 282510 537027 282558
rect 536981 282498 537027 282510
rect 538091 282510 538097 282558
rect 538131 282643 538137 282678
rect 538199 282678 538245 282690
rect 538199 282643 538205 282678
rect 538131 282558 538205 282643
rect 538131 282510 538137 282558
rect 538091 282498 538137 282510
rect 538199 282510 538205 282558
rect 538239 282643 538245 282678
rect 539309 282678 539355 282690
rect 539309 282643 539315 282678
rect 538239 282558 539315 282643
rect 538239 282510 538245 282558
rect 538199 282498 538245 282510
rect 539309 282510 539315 282558
rect 539349 282643 539355 282678
rect 539417 282678 539463 282690
rect 539417 282643 539423 282678
rect 539349 282558 539423 282643
rect 539349 282510 539355 282558
rect 539309 282498 539355 282510
rect 539417 282510 539423 282558
rect 539457 282643 539463 282678
rect 540527 282678 540573 282690
rect 540527 282643 540533 282678
rect 539457 282638 540533 282643
rect 539457 282568 540044 282638
rect 540114 282568 540154 282638
rect 540224 282568 540533 282638
rect 539457 282558 540533 282568
rect 539457 282510 539463 282558
rect 539417 282498 539463 282510
rect 540527 282510 540533 282558
rect 540567 282643 540573 282678
rect 540635 282678 540681 282690
rect 540635 282643 540641 282678
rect 540567 282558 540641 282643
rect 540567 282510 540573 282558
rect 540527 282498 540573 282510
rect 540635 282510 540641 282558
rect 540675 282643 540681 282678
rect 541745 282678 541791 282690
rect 541745 282643 541751 282678
rect 540675 282638 541751 282643
rect 540675 282568 540984 282638
rect 541054 282568 541094 282638
rect 541164 282568 541751 282638
rect 540675 282558 541751 282568
rect 540675 282510 540681 282558
rect 540635 282498 540681 282510
rect 541745 282510 541751 282558
rect 541785 282643 541791 282678
rect 541853 282678 541899 282690
rect 541853 282643 541859 282678
rect 541785 282558 541859 282643
rect 541785 282510 541791 282558
rect 541745 282498 541791 282510
rect 541853 282510 541859 282558
rect 541893 282643 541899 282678
rect 542963 282678 543009 282690
rect 542963 282643 542969 282678
rect 541893 282558 542969 282643
rect 541893 282510 541899 282558
rect 541853 282498 541899 282510
rect 542963 282510 542969 282558
rect 543003 282643 543009 282678
rect 543071 282678 543117 282690
rect 543071 282643 543077 282678
rect 543003 282558 543077 282643
rect 543003 282510 543009 282558
rect 542963 282498 543009 282510
rect 543071 282510 543077 282558
rect 543111 282643 543117 282678
rect 544181 282678 544227 282690
rect 544181 282643 544187 282678
rect 543111 282558 544187 282643
rect 543111 282510 543117 282558
rect 543071 282498 543117 282510
rect 544181 282510 544187 282558
rect 544221 282510 544227 282678
rect 544181 282498 544227 282510
rect 550420 282600 559740 282800
rect 537059 282482 538059 282488
rect 537059 282468 537071 282482
rect 537054 282448 537071 282468
rect 538047 282468 538059 282482
rect 538277 282482 539277 282488
rect 538277 282468 538289 282482
rect 538047 282448 538289 282468
rect 539265 282468 539277 282482
rect 539495 282482 540495 282488
rect 539495 282468 539507 282482
rect 539265 282448 539507 282468
rect 540483 282468 540495 282482
rect 540713 282482 541713 282488
rect 540713 282468 540725 282482
rect 540483 282448 540725 282468
rect 541701 282468 541713 282482
rect 541931 282482 542931 282488
rect 541931 282468 541943 282482
rect 541701 282448 541943 282468
rect 542919 282468 542931 282482
rect 543149 282482 544149 282488
rect 543149 282468 543161 282482
rect 542919 282448 543161 282468
rect 544137 282448 544149 282482
rect 537054 282442 544149 282448
rect 537054 282393 544144 282442
rect 550420 282400 557700 282600
rect 557900 282400 558100 282600
rect 558300 282400 558500 282600
rect 558700 282400 558900 282600
rect 559100 282400 559300 282600
rect 559500 282400 559740 282600
rect 538404 282098 538804 282393
rect 539804 282098 540204 282393
rect 541104 282098 541504 282393
rect 542394 282098 542804 282393
rect 550420 282340 559740 282400
rect 537604 281990 543604 282098
rect 537604 281984 540807 281990
rect 537604 281587 537777 281984
rect 538891 281587 539297 281984
rect 540411 281593 540807 281984
rect 541921 281593 542317 281990
rect 543431 281593 543604 281990
rect 540411 281587 543604 281593
rect 537604 281498 543604 281587
rect 567800 281384 568390 287604
rect 567800 281378 578400 281384
rect 567800 281344 570740 281378
rect 575880 281344 578400 281378
rect 567800 281334 578400 281344
rect 567800 281300 568280 281334
rect 567800 281100 567900 281300
rect 568100 281215 568280 281300
rect 572770 281284 572830 281294
rect 568310 281264 572770 281270
rect 572910 281284 572970 281294
rect 572830 281264 572910 281270
rect 573085 281284 573145 281294
rect 572970 281264 573085 281270
rect 573275 281284 573335 281294
rect 573145 281264 573275 281270
rect 573435 281284 573495 281294
rect 573335 281264 573435 281270
rect 573625 281284 573685 281294
rect 573495 281264 573625 281270
rect 573825 281284 573885 281294
rect 573685 281264 573825 281270
rect 574005 281284 574065 281294
rect 573885 281264 574005 281270
rect 574195 281284 574255 281294
rect 574065 281264 574195 281270
rect 574395 281284 574455 281294
rect 574255 281264 574395 281270
rect 574560 281274 574620 281284
rect 574455 281264 574560 281270
rect 574620 281264 578310 281270
rect 568310 281230 568322 281264
rect 578298 281230 578310 281264
rect 568310 281224 572770 281230
rect 572830 281224 572910 281230
rect 572970 281224 573085 281230
rect 573145 281224 573275 281230
rect 573335 281224 573435 281230
rect 573495 281224 573625 281230
rect 573685 281224 573825 281230
rect 573885 281224 574005 281230
rect 574065 281224 574195 281230
rect 574255 281224 574395 281230
rect 574455 281224 574560 281230
rect 568100 281181 568238 281215
rect 568272 281181 568280 281215
rect 572770 281214 572830 281224
rect 572910 281214 572970 281224
rect 573085 281214 573145 281224
rect 573275 281214 573335 281224
rect 573435 281214 573495 281224
rect 573625 281214 573685 281224
rect 573825 281214 573885 281224
rect 574005 281214 574065 281224
rect 574195 281214 574255 281224
rect 574395 281214 574455 281224
rect 574620 281224 578310 281230
rect 574560 281204 574620 281214
rect 568100 281174 568280 281181
rect 568100 281172 568330 281174
rect 578300 281172 578390 281174
rect 568100 281166 578390 281172
rect 568100 281132 568322 281166
rect 578298 281132 578390 281166
rect 568100 281126 578390 281132
rect 568100 281124 568330 281126
rect 578300 281124 578390 281126
rect 568100 281100 568280 281124
rect 537352 281058 537496 281064
rect 537352 280938 537364 281058
rect 537484 280938 537496 281058
rect 537352 280932 537496 280938
rect 543722 281058 543866 281064
rect 543722 280938 543734 281058
rect 543854 280938 543866 281058
rect 543722 280932 543866 280938
rect 567800 281050 568280 281100
rect 578342 281117 578390 281124
rect 572770 281084 572830 281094
rect 567800 281000 568136 281050
rect 567800 280800 567900 281000
rect 568100 280800 568136 281000
rect 567800 280700 568136 280800
rect 13060 280500 13280 280520
rect 13060 280430 13190 280500
rect 13260 280430 13280 280500
rect 13060 280390 13280 280430
rect 13060 280320 13080 280390
rect 13150 280320 13280 280390
rect 13060 279630 13280 280320
rect 567800 280500 567900 280700
rect 568100 280500 568136 280700
rect 567800 280464 568136 280500
rect 568170 281019 568280 281050
rect 568310 281068 572770 281074
rect 572910 281084 572970 281094
rect 572830 281068 572910 281074
rect 573085 281084 573145 281094
rect 572970 281068 573085 281074
rect 573275 281084 573335 281094
rect 573145 281068 573275 281074
rect 573435 281084 573495 281094
rect 573335 281068 573435 281074
rect 573625 281084 573685 281094
rect 573495 281068 573625 281074
rect 573825 281084 573885 281094
rect 573685 281068 573825 281074
rect 574005 281084 574065 281094
rect 573885 281068 574005 281074
rect 574195 281084 574255 281094
rect 574065 281068 574195 281074
rect 574395 281084 574455 281094
rect 574255 281068 574395 281074
rect 574560 281084 574620 281094
rect 574455 281068 574560 281074
rect 578342 281083 578348 281117
rect 578382 281083 578390 281117
rect 574620 281068 578310 281074
rect 578342 281071 578390 281083
rect 568310 281034 568322 281068
rect 578298 281034 578310 281068
rect 568310 281028 572770 281034
rect 568170 280985 568238 281019
rect 568272 280985 568280 281019
rect 572830 281028 572910 281034
rect 572770 281014 572830 281024
rect 572970 281028 573085 281034
rect 572910 281014 572970 281024
rect 573145 281028 573275 281034
rect 573085 281014 573145 281024
rect 573335 281028 573435 281034
rect 573275 281014 573335 281024
rect 573495 281028 573625 281034
rect 573435 281014 573495 281024
rect 573685 281028 573825 281034
rect 573625 281014 573685 281024
rect 573885 281028 574005 281034
rect 573825 281014 573885 281024
rect 574065 281028 574195 281034
rect 574005 281014 574065 281024
rect 574255 281028 574395 281034
rect 574195 281014 574255 281024
rect 574455 281028 574560 281034
rect 574395 281014 574455 281024
rect 574620 281028 578310 281034
rect 574560 281014 574620 281024
rect 568170 280984 568280 280985
rect 568170 280976 568330 280984
rect 568170 280974 578310 280976
rect 578350 280974 578390 281071
rect 568170 280970 578390 280974
rect 568170 280936 568322 280970
rect 578298 280936 578390 280970
rect 568170 280930 578390 280936
rect 568170 280924 568330 280930
rect 578300 280924 578390 280930
rect 568170 280823 568280 280924
rect 578342 280921 578390 280924
rect 572770 280884 572830 280894
rect 568310 280872 572770 280878
rect 572910 280884 572970 280894
rect 572830 280872 572910 280878
rect 573085 280884 573145 280894
rect 572970 280872 573085 280878
rect 573275 280884 573335 280894
rect 573145 280872 573275 280878
rect 573435 280884 573495 280894
rect 573335 280872 573435 280878
rect 573625 280884 573685 280894
rect 573495 280872 573625 280878
rect 573825 280884 573885 280894
rect 573685 280872 573825 280878
rect 574005 280884 574065 280894
rect 573885 280872 574005 280878
rect 574195 280884 574255 280894
rect 574065 280872 574195 280878
rect 574395 280884 574455 280894
rect 574255 280872 574395 280878
rect 574560 280884 574620 280894
rect 574455 280872 574560 280878
rect 578342 280887 578348 280921
rect 578382 280887 578390 280921
rect 574620 280872 578310 280878
rect 578342 280875 578390 280887
rect 568310 280838 568322 280872
rect 578298 280838 578310 280872
rect 568310 280832 572770 280838
rect 568170 280789 568238 280823
rect 568272 280789 568280 280823
rect 572830 280832 572910 280838
rect 572770 280814 572830 280824
rect 572970 280832 573085 280838
rect 572910 280814 572970 280824
rect 573145 280832 573275 280838
rect 573085 280814 573145 280824
rect 573335 280832 573435 280838
rect 573275 280814 573335 280824
rect 573495 280832 573625 280838
rect 573435 280814 573495 280824
rect 573685 280832 573825 280838
rect 573625 280814 573685 280824
rect 573885 280832 574005 280838
rect 573825 280814 573885 280824
rect 574065 280832 574195 280838
rect 574005 280814 574065 280824
rect 574255 280832 574395 280838
rect 574195 280814 574255 280824
rect 574455 280832 574560 280838
rect 574395 280814 574455 280824
rect 574620 280832 578310 280838
rect 574560 280814 574620 280824
rect 568170 280784 568280 280789
rect 578350 280784 578390 280875
rect 568170 280780 568330 280784
rect 578300 280780 578390 280784
rect 568170 280774 578390 280780
rect 568170 280740 568322 280774
rect 578298 280740 578390 280774
rect 568170 280734 578390 280740
rect 568170 280724 568330 280734
rect 578342 280725 578390 280734
rect 568170 280627 568280 280724
rect 572770 280694 572830 280704
rect 568310 280676 572770 280682
rect 572910 280694 572970 280704
rect 572830 280676 572910 280682
rect 573085 280694 573145 280704
rect 572970 280676 573085 280682
rect 573275 280694 573335 280704
rect 573145 280676 573275 280682
rect 573435 280694 573495 280704
rect 573335 280676 573435 280682
rect 573625 280694 573685 280704
rect 573495 280676 573625 280682
rect 573825 280694 573885 280704
rect 573685 280676 573825 280682
rect 574005 280694 574065 280704
rect 573885 280676 574005 280682
rect 574195 280694 574255 280704
rect 574065 280676 574195 280682
rect 574395 280694 574455 280704
rect 574255 280676 574395 280682
rect 574560 280694 574620 280704
rect 574455 280676 574560 280682
rect 578342 280691 578348 280725
rect 578382 280691 578390 280725
rect 574620 280676 578310 280682
rect 578342 280679 578390 280691
rect 568310 280642 568322 280676
rect 578298 280642 578310 280676
rect 568310 280636 572770 280642
rect 568170 280593 568238 280627
rect 568272 280594 568280 280627
rect 572830 280636 572910 280642
rect 572770 280624 572830 280634
rect 572970 280636 573085 280642
rect 572910 280624 572970 280634
rect 573145 280636 573275 280642
rect 573085 280624 573145 280634
rect 573335 280636 573435 280642
rect 573275 280624 573335 280634
rect 573495 280636 573625 280642
rect 573435 280624 573495 280634
rect 573685 280636 573825 280642
rect 573625 280624 573685 280634
rect 573885 280636 574005 280642
rect 573825 280624 573885 280634
rect 574065 280636 574195 280642
rect 574005 280624 574065 280634
rect 574255 280636 574395 280642
rect 574195 280624 574255 280634
rect 574455 280636 574560 280642
rect 574395 280624 574455 280634
rect 574620 280636 578310 280642
rect 574560 280624 574620 280634
rect 568272 280593 568330 280594
rect 568170 280584 568330 280593
rect 578350 280584 578390 280679
rect 568170 280578 578390 280584
rect 568170 280544 568322 280578
rect 578298 280544 578390 280578
rect 568170 280538 578390 280544
rect 568170 280534 568330 280538
rect 578300 280534 578390 280538
rect 568170 280464 568280 280534
rect 578342 280529 578390 280534
rect 572770 280494 572830 280504
rect 567800 280431 568280 280464
rect 568310 280480 572770 280486
rect 572910 280494 572970 280504
rect 572830 280480 572910 280486
rect 573085 280494 573145 280504
rect 572970 280480 573085 280486
rect 573275 280494 573335 280504
rect 573145 280480 573275 280486
rect 573435 280494 573495 280504
rect 573335 280480 573435 280486
rect 573625 280494 573685 280504
rect 573495 280480 573625 280486
rect 573825 280494 573885 280504
rect 573685 280480 573825 280486
rect 574005 280494 574065 280504
rect 573885 280480 574005 280486
rect 574195 280494 574255 280504
rect 574065 280480 574195 280486
rect 574395 280494 574455 280504
rect 574255 280480 574395 280486
rect 574560 280494 574620 280504
rect 574455 280480 574560 280486
rect 578342 280495 578348 280529
rect 578382 280495 578390 280529
rect 574620 280480 578310 280486
rect 578342 280483 578390 280495
rect 568310 280446 568322 280480
rect 578298 280446 578310 280480
rect 568310 280440 572770 280446
rect 567800 280400 568238 280431
rect 567800 280200 567900 280400
rect 568100 280397 568238 280400
rect 568272 280397 568280 280431
rect 572830 280440 572910 280446
rect 572770 280424 572830 280434
rect 572970 280440 573085 280446
rect 572910 280424 572970 280434
rect 573145 280440 573275 280446
rect 573085 280424 573145 280434
rect 573335 280440 573435 280446
rect 573275 280424 573335 280434
rect 573495 280440 573625 280446
rect 573435 280424 573495 280434
rect 573685 280440 573825 280446
rect 573625 280424 573685 280434
rect 573885 280440 574005 280446
rect 573825 280424 573885 280434
rect 574065 280440 574195 280446
rect 574005 280424 574065 280434
rect 574255 280440 574395 280446
rect 574195 280424 574255 280434
rect 574455 280440 574560 280446
rect 574395 280424 574455 280434
rect 574620 280440 578310 280446
rect 574560 280424 574620 280434
rect 568100 280394 568280 280397
rect 578350 280394 578390 280483
rect 568100 280388 568330 280394
rect 578300 280388 578390 280394
rect 568100 280382 578390 280388
rect 568100 280348 568322 280382
rect 578298 280348 578390 280382
rect 568100 280344 578390 280348
rect 568100 280342 578310 280344
rect 568100 280334 568330 280342
rect 568100 280200 568280 280334
rect 578342 280333 578390 280344
rect 572770 280294 572830 280304
rect 568310 280284 572770 280290
rect 572910 280294 572970 280304
rect 572830 280284 572910 280290
rect 573085 280294 573145 280304
rect 572970 280284 573085 280290
rect 573275 280294 573335 280304
rect 573145 280284 573275 280290
rect 573435 280294 573495 280304
rect 573335 280284 573435 280290
rect 573625 280294 573685 280304
rect 573495 280284 573625 280290
rect 573825 280294 573885 280304
rect 573685 280284 573825 280290
rect 574005 280294 574065 280304
rect 573885 280284 574005 280290
rect 574195 280294 574255 280304
rect 574065 280284 574195 280290
rect 574395 280294 574455 280304
rect 574255 280284 574395 280290
rect 574560 280294 574620 280304
rect 574455 280284 574560 280290
rect 578342 280299 578348 280333
rect 578382 280299 578390 280333
rect 574620 280284 578310 280290
rect 578342 280287 578390 280299
rect 578350 280284 578390 280287
rect 568310 280250 568322 280284
rect 578298 280250 578310 280284
rect 568310 280244 572770 280250
rect 572830 280244 572910 280250
rect 572770 280224 572830 280234
rect 572970 280244 573085 280250
rect 572910 280224 572970 280234
rect 573145 280244 573275 280250
rect 573085 280224 573145 280234
rect 573335 280244 573435 280250
rect 573275 280224 573335 280234
rect 573495 280244 573625 280250
rect 573435 280224 573495 280234
rect 573685 280244 573825 280250
rect 573625 280224 573685 280234
rect 573885 280244 574005 280250
rect 573825 280224 573885 280234
rect 574065 280244 574195 280250
rect 574005 280224 574065 280234
rect 574255 280244 574395 280250
rect 574195 280224 574255 280234
rect 574455 280244 574560 280250
rect 574395 280224 574455 280234
rect 574620 280244 578310 280250
rect 574560 280224 574620 280234
rect 567800 280174 568280 280200
rect 570728 280174 575892 280176
rect 567800 280170 578400 280174
rect 567800 280136 570740 280170
rect 575880 280136 578400 280170
rect 567800 280124 578400 280136
rect 567800 280100 568280 280124
rect 11870 279609 14480 279630
rect 11870 279212 11887 279609
rect 13001 279212 13347 279609
rect 14461 279212 14480 279609
rect 11870 279190 14480 279212
rect 14534 278550 14646 278562
rect 14534 278370 14540 278550
rect 14640 278370 14646 278550
rect 14534 278358 14646 278370
rect 14534 278130 14646 278142
rect 14534 277950 14540 278130
rect 14640 277950 14646 278130
rect 14534 277938 14646 277950
rect 537352 278058 537496 278064
rect 537352 277938 537364 278058
rect 537484 277938 537496 278058
rect 537352 277932 537496 277938
rect 543722 278058 543866 278064
rect 543722 277938 543734 278058
rect 543854 277938 543866 278058
rect 543722 277932 543866 277938
rect 11870 277178 14480 277190
rect 11870 276781 11887 277178
rect 13001 276781 13347 277178
rect 14461 276781 14480 277178
rect 11870 276760 14480 276781
rect 13140 275990 13430 276760
rect 31014 276140 31266 276152
rect 12710 275910 13890 275990
rect 12710 275772 12760 275910
rect 12840 275850 12910 275860
rect 12801 275834 12840 275840
rect 13080 275850 13150 275860
rect 12910 275834 13080 275840
rect 13150 275834 13801 275840
rect 12801 275800 12813 275834
rect 13789 275800 13801 275834
rect 12801 275794 12840 275800
rect 12710 275704 12720 275772
rect 12754 275704 12760 275772
rect 12910 275794 13080 275800
rect 12840 275770 12910 275780
rect 13150 275794 13801 275800
rect 13080 275770 13150 275780
rect 13840 275772 13890 275910
rect 31014 275900 31020 276140
rect 31260 275900 31266 276140
rect 31014 275888 31266 275900
rect 32734 276140 32986 276152
rect 32734 275900 32740 276140
rect 32980 275900 32986 276140
rect 32734 275888 32986 275900
rect 34454 276140 34706 276152
rect 34454 275900 34460 276140
rect 34700 275900 34706 276140
rect 34454 275888 34706 275900
rect 35934 276140 36186 276152
rect 35934 275900 35940 276140
rect 36180 275900 36186 276140
rect 35934 275888 36186 275900
rect 37654 276140 37906 276152
rect 37654 275900 37660 276140
rect 37900 275900 37906 276140
rect 37654 275888 37906 275900
rect 39254 276140 39506 276152
rect 39254 275900 39260 276140
rect 39500 275900 39506 276140
rect 39254 275888 39506 275900
rect 40974 276140 41226 276152
rect 40974 275900 40980 276140
rect 41220 275900 41226 276140
rect 40974 275888 41226 275900
rect 42574 276140 42826 276152
rect 42574 275900 42580 276140
rect 42820 275900 42826 276140
rect 42574 275888 42826 275900
rect 44294 276140 44546 276152
rect 44294 275900 44300 276140
rect 44540 275900 44546 276140
rect 44294 275888 44546 275900
rect 44600 276140 45200 276300
rect 44600 275900 44780 276140
rect 45020 275900 45200 276140
rect 12710 275614 12760 275704
rect 13450 275700 13520 275710
rect 12801 275676 13450 275682
rect 13690 275700 13760 275710
rect 13520 275676 13690 275682
rect 13840 275704 13848 275772
rect 13882 275704 13890 275772
rect 13760 275676 13801 275682
rect 12801 275642 12813 275676
rect 13789 275642 13801 275676
rect 12801 275636 13450 275642
rect 13520 275636 13690 275642
rect 13450 275620 13520 275630
rect 13760 275636 13801 275642
rect 13690 275620 13760 275630
rect 12710 275546 12720 275614
rect 12754 275546 12760 275614
rect 13840 275614 13890 275704
rect 12710 275456 12760 275546
rect 12840 275540 12910 275550
rect 12801 275518 12840 275524
rect 13080 275540 13150 275550
rect 12910 275518 13080 275524
rect 13840 275546 13848 275614
rect 13882 275546 13890 275614
rect 13150 275518 13801 275524
rect 12801 275484 12813 275518
rect 13789 275484 13801 275518
rect 12801 275478 12840 275484
rect 12910 275478 13080 275484
rect 12840 275460 12910 275470
rect 13150 275478 13801 275484
rect 13080 275460 13150 275470
rect 12710 275388 12720 275456
rect 12754 275388 12760 275456
rect 13840 275456 13890 275546
rect 12710 275298 12760 275388
rect 13450 275380 13520 275390
rect 12801 275360 13450 275366
rect 13690 275380 13760 275390
rect 13520 275360 13690 275366
rect 13840 275388 13848 275456
rect 13882 275388 13890 275456
rect 13760 275360 13801 275366
rect 12801 275326 12813 275360
rect 13789 275326 13801 275360
rect 12801 275320 13450 275326
rect 13520 275320 13690 275326
rect 13450 275300 13520 275310
rect 13760 275320 13801 275326
rect 13690 275300 13760 275310
rect 12710 275230 12720 275298
rect 12754 275230 12760 275298
rect 13840 275298 13890 275388
rect 13840 275230 13848 275298
rect 13882 275230 13890 275298
rect 12710 275140 12760 275230
rect 12840 275220 12910 275230
rect 12801 275202 12840 275208
rect 13080 275220 13150 275230
rect 12910 275202 13080 275208
rect 13150 275202 13801 275208
rect 12801 275168 12813 275202
rect 13789 275168 13801 275202
rect 12801 275162 12840 275168
rect 12910 275162 13080 275168
rect 12840 275140 12910 275150
rect 13150 275162 13801 275168
rect 13080 275140 13150 275150
rect 13840 275140 13890 275230
rect 12710 275072 12720 275140
rect 12754 275072 12760 275140
rect 12710 274982 12760 275072
rect 13840 275072 13848 275140
rect 13882 275072 13890 275140
rect 17600 275300 18600 275400
rect 17600 275200 17700 275300
rect 17800 275200 18000 275300
rect 18200 275200 18400 275300
rect 18500 275200 18600 275300
rect 17600 275100 18600 275200
rect 13450 275060 13520 275070
rect 12801 275044 13450 275050
rect 13690 275060 13760 275070
rect 13520 275044 13690 275050
rect 13760 275044 13801 275050
rect 12801 275010 12813 275044
rect 13789 275010 13801 275044
rect 12801 275004 13450 275010
rect 12710 274914 12720 274982
rect 12754 274914 12760 274982
rect 13520 275004 13690 275010
rect 13450 274980 13520 274990
rect 13760 275004 13801 275010
rect 13690 274980 13760 274990
rect 13840 274982 13890 275072
rect 12710 274824 12760 274914
rect 13840 274914 13848 274982
rect 13882 274914 13890 274982
rect 12840 274900 12910 274910
rect 12801 274886 12840 274892
rect 13080 274900 13150 274910
rect 12910 274886 13080 274892
rect 13150 274886 13801 274892
rect 12801 274852 12813 274886
rect 13789 274852 13801 274886
rect 12801 274846 12840 274852
rect 12710 274756 12720 274824
rect 12754 274756 12760 274824
rect 12910 274846 13080 274852
rect 12840 274820 12910 274830
rect 13150 274846 13801 274852
rect 13080 274820 13150 274830
rect 13840 274824 13890 274914
rect 12710 274666 12760 274756
rect 13450 274750 13520 274760
rect 12801 274728 13450 274734
rect 13690 274750 13760 274760
rect 13520 274728 13690 274734
rect 13840 274756 13848 274824
rect 13882 274760 13890 274824
rect 13882 274756 13950 274760
rect 13760 274728 13801 274734
rect 12801 274694 12813 274728
rect 13789 274694 13801 274728
rect 12801 274688 13450 274694
rect 13520 274688 13690 274694
rect 13450 274670 13520 274680
rect 13760 274688 13801 274694
rect 13840 274720 13950 274756
rect 13690 274670 13760 274680
rect 12710 274598 12720 274666
rect 12754 274598 12760 274666
rect 13840 274666 13860 274720
rect 12710 274508 12760 274598
rect 12840 274590 12910 274600
rect 12801 274570 12840 274576
rect 13080 274590 13150 274600
rect 12910 274570 13080 274576
rect 13840 274598 13848 274666
rect 13940 274640 13950 274720
rect 13882 274600 13950 274640
rect 13882 274598 13890 274600
rect 13150 274570 13801 274576
rect 12801 274536 12813 274570
rect 13789 274536 13801 274570
rect 12801 274530 12840 274536
rect 12910 274530 13080 274536
rect 12840 274510 12910 274520
rect 13150 274530 13801 274536
rect 13080 274510 13150 274520
rect 12710 274440 12720 274508
rect 12754 274440 12760 274508
rect 13840 274508 13890 274598
rect 13840 274440 13848 274508
rect 13882 274440 13890 274508
rect 12710 274350 12760 274440
rect 13450 274430 13520 274440
rect 12801 274412 13450 274418
rect 13690 274430 13760 274440
rect 13520 274412 13690 274418
rect 13760 274412 13801 274418
rect 12801 274378 12813 274412
rect 13789 274378 13801 274412
rect 12801 274372 13450 274378
rect 13520 274372 13690 274378
rect 13450 274350 13520 274360
rect 13760 274372 13801 274378
rect 13690 274350 13760 274360
rect 13840 274350 13890 274440
rect 12612 274285 12658 274297
rect 12612 273360 12618 274285
rect 12310 273330 12618 273360
rect 12310 273060 12360 273330
rect 12310 272280 12618 273060
rect 12310 272010 12360 272280
rect 12310 271980 12618 272010
rect 12612 271029 12618 271980
rect 12652 271029 12658 274285
rect 12612 271017 12658 271029
rect 12710 274282 12720 274350
rect 12754 274282 12760 274350
rect 12710 274192 12760 274282
rect 13840 274282 13848 274350
rect 13882 274282 13890 274350
rect 14380 274400 15560 274480
rect 12840 274270 12910 274280
rect 12801 274254 12840 274260
rect 13080 274270 13150 274280
rect 12910 274254 13080 274260
rect 13150 274254 13801 274260
rect 12801 274220 12813 274254
rect 13789 274220 13801 274254
rect 12801 274214 12840 274220
rect 12710 274124 12720 274192
rect 12754 274124 12760 274192
rect 12910 274214 13080 274220
rect 12840 274190 12910 274200
rect 13150 274214 13801 274220
rect 13080 274190 13150 274200
rect 13840 274192 13890 274282
rect 12710 274034 12760 274124
rect 13840 274124 13848 274192
rect 13882 274124 13890 274192
rect 13450 274110 13520 274120
rect 12801 274096 13450 274102
rect 13690 274110 13760 274120
rect 13520 274096 13690 274102
rect 13760 274096 13801 274102
rect 12801 274062 12813 274096
rect 13789 274062 13801 274096
rect 12801 274056 13450 274062
rect 12710 273966 12720 274034
rect 12754 273966 12760 274034
rect 13520 274056 13690 274062
rect 13450 274030 13520 274040
rect 13760 274056 13801 274062
rect 13690 274030 13760 274040
rect 13840 274034 13890 274124
rect 12710 273876 12760 273966
rect 12840 273960 12910 273970
rect 12801 273938 12840 273944
rect 13080 273960 13150 273970
rect 12910 273938 13080 273944
rect 13840 273966 13848 274034
rect 13882 273966 13890 274034
rect 13150 273938 13801 273944
rect 12801 273904 12813 273938
rect 13789 273904 13801 273938
rect 12801 273898 12840 273904
rect 12910 273898 13080 273904
rect 12840 273880 12910 273890
rect 13150 273898 13801 273904
rect 13080 273880 13150 273890
rect 12710 273808 12720 273876
rect 12754 273808 12760 273876
rect 13840 273876 13890 273966
rect 12710 273718 12760 273808
rect 13450 273800 13520 273810
rect 12801 273780 13450 273786
rect 13690 273800 13760 273810
rect 13520 273780 13690 273786
rect 13840 273808 13848 273876
rect 13882 273808 13890 273876
rect 13760 273780 13801 273786
rect 12801 273746 12813 273780
rect 13789 273746 13801 273780
rect 12801 273740 13450 273746
rect 13520 273740 13690 273746
rect 13450 273720 13520 273730
rect 13760 273740 13801 273746
rect 13690 273720 13760 273730
rect 12710 273650 12720 273718
rect 12754 273650 12760 273718
rect 13840 273718 13890 273808
rect 13840 273650 13848 273718
rect 13882 273650 13890 273718
rect 12710 273560 12760 273650
rect 12840 273640 12910 273650
rect 12801 273622 12840 273628
rect 13080 273640 13150 273650
rect 12910 273622 13080 273628
rect 13150 273622 13801 273628
rect 12801 273588 12813 273622
rect 13789 273588 13801 273622
rect 12801 273582 12840 273588
rect 12910 273582 13080 273588
rect 12840 273560 12910 273570
rect 13150 273582 13801 273588
rect 13080 273560 13150 273570
rect 13840 273560 13890 273650
rect 12710 273492 12720 273560
rect 12754 273492 12760 273560
rect 12710 273402 12760 273492
rect 13840 273492 13848 273560
rect 13882 273492 13890 273560
rect 13944 274285 13990 274297
rect 13944 273550 13950 274285
rect 13450 273480 13520 273490
rect 12801 273464 13450 273470
rect 13690 273480 13760 273490
rect 13520 273464 13690 273470
rect 13760 273464 13801 273470
rect 12801 273430 12813 273464
rect 13789 273430 13801 273464
rect 12801 273424 13450 273430
rect 12710 273334 12720 273402
rect 12754 273334 12760 273402
rect 13520 273424 13690 273430
rect 13450 273400 13520 273410
rect 13760 273424 13801 273430
rect 13690 273400 13760 273410
rect 13840 273402 13890 273492
rect 12710 273244 12760 273334
rect 13840 273334 13848 273402
rect 13882 273334 13890 273402
rect 12840 273320 12910 273330
rect 12801 273306 12840 273312
rect 13080 273320 13150 273330
rect 12910 273306 13080 273312
rect 13150 273306 13801 273312
rect 12801 273272 12813 273306
rect 13789 273272 13801 273306
rect 12801 273266 12840 273272
rect 12710 273176 12720 273244
rect 12754 273176 12760 273244
rect 12910 273266 13080 273272
rect 12840 273240 12910 273250
rect 13150 273266 13801 273272
rect 13080 273240 13150 273250
rect 13840 273244 13890 273334
rect 12710 273086 12760 273176
rect 13450 273170 13520 273180
rect 12801 273148 13450 273154
rect 13690 273170 13760 273180
rect 13520 273148 13690 273154
rect 13840 273176 13848 273244
rect 13882 273176 13890 273244
rect 13760 273148 13801 273154
rect 12801 273114 12813 273148
rect 13789 273114 13801 273148
rect 12801 273108 13450 273114
rect 13520 273108 13690 273114
rect 13450 273090 13520 273100
rect 13760 273108 13801 273114
rect 13690 273090 13760 273100
rect 12710 273018 12720 273086
rect 12754 273018 12760 273086
rect 13840 273086 13890 273176
rect 12710 272928 12760 273018
rect 12840 273010 12910 273020
rect 12801 272990 12840 272996
rect 13080 273010 13150 273020
rect 12910 272990 13080 272996
rect 13840 273018 13848 273086
rect 13882 273018 13890 273086
rect 13150 272990 13801 272996
rect 12801 272956 12813 272990
rect 13789 272956 13801 272990
rect 12801 272950 12840 272956
rect 12910 272950 13080 272956
rect 12840 272930 12910 272940
rect 13150 272950 13801 272956
rect 13080 272930 13150 272940
rect 12710 272860 12720 272928
rect 12754 272860 12760 272928
rect 13840 272928 13890 273018
rect 13840 272860 13848 272928
rect 13882 272860 13890 272928
rect 12710 272770 12760 272860
rect 13450 272850 13520 272860
rect 12801 272832 13450 272838
rect 13690 272850 13760 272860
rect 13520 272832 13690 272838
rect 13760 272832 13801 272838
rect 12801 272798 12813 272832
rect 13789 272798 13801 272832
rect 12801 272792 13450 272798
rect 13520 272792 13690 272798
rect 13450 272770 13520 272780
rect 13760 272792 13801 272798
rect 13690 272770 13760 272780
rect 13840 272770 13890 272860
rect 12710 272702 12720 272770
rect 12754 272702 12760 272770
rect 12710 272612 12760 272702
rect 13840 272702 13848 272770
rect 13882 272702 13890 272770
rect 12840 272690 12910 272700
rect 12801 272674 12840 272680
rect 13080 272690 13150 272700
rect 12910 272674 13080 272680
rect 13150 272674 13801 272680
rect 12801 272640 12813 272674
rect 13789 272640 13801 272674
rect 12801 272634 12840 272640
rect 12710 272544 12720 272612
rect 12754 272544 12760 272612
rect 12910 272634 13080 272640
rect 12840 272610 12910 272620
rect 13150 272634 13801 272640
rect 13080 272610 13150 272620
rect 13840 272612 13890 272702
rect 12710 272454 12760 272544
rect 13840 272544 13848 272612
rect 13882 272544 13890 272612
rect 13450 272530 13520 272540
rect 12801 272516 13450 272522
rect 13690 272530 13760 272540
rect 13520 272516 13690 272522
rect 13760 272516 13801 272522
rect 12801 272482 12813 272516
rect 13789 272482 13801 272516
rect 12801 272476 13450 272482
rect 12710 272386 12720 272454
rect 12754 272386 12760 272454
rect 13520 272476 13690 272482
rect 13450 272450 13520 272460
rect 13760 272476 13801 272482
rect 13690 272450 13760 272460
rect 13840 272454 13890 272544
rect 12710 272296 12760 272386
rect 12840 272380 12910 272390
rect 12801 272358 12840 272364
rect 13080 272380 13150 272390
rect 12910 272358 13080 272364
rect 13840 272386 13848 272454
rect 13882 272386 13890 272454
rect 13150 272358 13801 272364
rect 12801 272324 12813 272358
rect 13789 272324 13801 272358
rect 12801 272318 12840 272324
rect 12910 272318 13080 272324
rect 12840 272300 12910 272310
rect 13150 272318 13801 272324
rect 13080 272300 13150 272310
rect 12710 272228 12720 272296
rect 12754 272228 12760 272296
rect 13840 272296 13890 272386
rect 12710 272138 12760 272228
rect 13450 272220 13520 272230
rect 12801 272200 13450 272206
rect 13690 272220 13760 272230
rect 13520 272200 13690 272206
rect 13840 272228 13848 272296
rect 13882 272228 13890 272296
rect 13760 272200 13801 272206
rect 12801 272166 12813 272200
rect 13789 272166 13801 272200
rect 12801 272160 13450 272166
rect 13520 272160 13690 272166
rect 13450 272140 13520 272150
rect 13760 272160 13801 272166
rect 13690 272140 13760 272150
rect 12710 272070 12720 272138
rect 12754 272070 12760 272138
rect 13840 272138 13890 272228
rect 13840 272070 13848 272138
rect 13882 272070 13890 272138
rect 12710 271980 12760 272070
rect 12840 272060 12910 272070
rect 12801 272042 12840 272048
rect 13080 272060 13150 272070
rect 12910 272042 13080 272048
rect 13150 272042 13801 272048
rect 12801 272008 12813 272042
rect 13789 272008 13801 272042
rect 12801 272002 12840 272008
rect 12910 272002 13080 272008
rect 12840 271980 12910 271990
rect 13150 272002 13801 272008
rect 13080 271980 13150 271990
rect 13840 271980 13890 272070
rect 12710 271912 12720 271980
rect 12754 271912 12760 271980
rect 12710 271822 12760 271912
rect 13840 271912 13848 271980
rect 13882 271912 13890 271980
rect 13450 271900 13520 271910
rect 12801 271884 13450 271890
rect 13690 271900 13760 271910
rect 13520 271884 13690 271890
rect 13760 271884 13801 271890
rect 12801 271850 12813 271884
rect 13789 271850 13801 271884
rect 12801 271844 13450 271850
rect 12710 271754 12720 271822
rect 12754 271754 12760 271822
rect 13520 271844 13690 271850
rect 13450 271820 13520 271830
rect 13760 271844 13801 271850
rect 13690 271820 13760 271830
rect 13840 271822 13890 271912
rect 12710 271664 12760 271754
rect 13840 271754 13848 271822
rect 13882 271754 13890 271822
rect 13940 271760 13950 273550
rect 12840 271740 12910 271750
rect 12801 271726 12840 271732
rect 13080 271740 13150 271750
rect 12910 271726 13080 271732
rect 13150 271726 13801 271732
rect 12801 271692 12813 271726
rect 13789 271692 13801 271726
rect 12801 271686 12840 271692
rect 12710 271596 12720 271664
rect 12754 271596 12760 271664
rect 12910 271686 13080 271692
rect 12840 271660 12910 271670
rect 13150 271686 13801 271692
rect 13080 271660 13150 271670
rect 13840 271664 13890 271754
rect 12710 271506 12760 271596
rect 13840 271596 13848 271664
rect 13882 271596 13890 271664
rect 13450 271580 13520 271590
rect 12801 271568 13450 271574
rect 13690 271580 13760 271590
rect 13520 271568 13690 271574
rect 13760 271568 13801 271574
rect 12801 271534 12813 271568
rect 13789 271534 13801 271568
rect 12801 271528 13450 271534
rect 12710 271438 12720 271506
rect 12754 271438 12760 271506
rect 13520 271528 13690 271534
rect 13450 271500 13520 271510
rect 13760 271528 13801 271534
rect 13690 271500 13760 271510
rect 13840 271506 13890 271596
rect 12710 271348 12760 271438
rect 12840 271430 12910 271440
rect 12801 271410 12840 271416
rect 13080 271430 13150 271440
rect 12910 271410 13080 271416
rect 13840 271438 13848 271506
rect 13882 271438 13890 271506
rect 13150 271410 13801 271416
rect 12801 271376 12813 271410
rect 13789 271376 13801 271410
rect 12801 271370 12840 271376
rect 12910 271370 13080 271376
rect 12840 271350 12910 271360
rect 13150 271370 13801 271376
rect 13080 271350 13150 271360
rect 12710 271280 12720 271348
rect 12754 271280 12760 271348
rect 13840 271348 13890 271438
rect 13840 271280 13848 271348
rect 13882 271280 13890 271348
rect 12710 271190 12760 271280
rect 13450 271270 13520 271280
rect 12801 271252 13450 271258
rect 13690 271270 13760 271280
rect 13520 271252 13690 271258
rect 13760 271252 13801 271258
rect 12801 271218 12813 271252
rect 13789 271218 13801 271252
rect 12801 271212 13450 271218
rect 13520 271212 13690 271218
rect 13450 271190 13520 271200
rect 13760 271212 13801 271218
rect 13690 271190 13760 271200
rect 13840 271190 13890 271280
rect 12710 271122 12720 271190
rect 12754 271122 12760 271190
rect 12710 271032 12760 271122
rect 13840 271122 13848 271190
rect 13882 271122 13890 271190
rect 12840 271110 12910 271120
rect 12801 271094 12840 271100
rect 13080 271110 13150 271120
rect 12910 271094 13080 271100
rect 13150 271094 13801 271100
rect 12801 271060 12813 271094
rect 13789 271060 13801 271094
rect 12801 271054 12840 271060
rect 12710 270964 12720 271032
rect 12754 270964 12760 271032
rect 12910 271054 13080 271060
rect 12840 271030 12910 271040
rect 13150 271054 13801 271060
rect 13080 271030 13150 271040
rect 13840 271032 13890 271122
rect 12710 270874 12760 270964
rect 13840 270964 13848 271032
rect 13882 270964 13890 271032
rect 13944 271029 13950 271760
rect 13984 273550 13990 274285
rect 14380 274270 14430 274400
rect 15150 274350 15220 274360
rect 14471 274332 15150 274338
rect 15360 274350 15430 274360
rect 15220 274332 15360 274338
rect 15430 274332 15471 274338
rect 14471 274298 14483 274332
rect 15459 274298 15471 274332
rect 14471 274292 15150 274298
rect 15220 274292 15360 274298
rect 15150 274270 15220 274280
rect 15430 274292 15471 274298
rect 15360 274270 15430 274280
rect 15510 274290 15560 274400
rect 16690 274350 16760 274360
rect 16011 274332 16690 274338
rect 16900 274350 16970 274360
rect 16760 274332 16900 274338
rect 16970 274332 17011 274338
rect 16011 274298 16023 274332
rect 16999 274298 17011 274332
rect 16011 274292 16690 274298
rect 15510 274270 15970 274290
rect 16760 274292 16900 274298
rect 16690 274270 16760 274280
rect 16970 274292 17011 274298
rect 16900 274270 16970 274280
rect 17050 274270 17100 274290
rect 14380 274202 14390 274270
rect 14424 274202 14430 274270
rect 14380 274112 14430 274202
rect 15510 274202 15518 274270
rect 15552 274202 15930 274270
rect 15964 274202 15970 274270
rect 14510 274190 14580 274200
rect 14471 274174 14510 274180
rect 14720 274190 14790 274200
rect 14580 274174 14720 274180
rect 14790 274174 15471 274180
rect 14471 274140 14483 274174
rect 15459 274140 15471 274174
rect 14471 274134 14510 274140
rect 14380 274044 14390 274112
rect 14424 274044 14430 274112
rect 14580 274134 14720 274140
rect 14510 274110 14580 274120
rect 14790 274134 15471 274140
rect 14720 274110 14790 274120
rect 15510 274112 15970 274202
rect 17050 274202 17058 274270
rect 17092 274202 17100 274270
rect 16060 274190 16130 274200
rect 16011 274174 16060 274180
rect 16270 274190 16340 274200
rect 16130 274174 16270 274180
rect 16340 274174 17011 274180
rect 16011 274140 16023 274174
rect 16999 274140 17011 274174
rect 16011 274134 16060 274140
rect 14380 273954 14430 274044
rect 15150 274040 15220 274050
rect 14471 274016 15150 274022
rect 15360 274040 15430 274050
rect 15220 274016 15360 274022
rect 15510 274044 15518 274112
rect 15552 274044 15930 274112
rect 15964 274044 15970 274112
rect 16130 274134 16270 274140
rect 16060 274110 16130 274120
rect 16340 274134 17011 274140
rect 16270 274110 16340 274120
rect 17050 274112 17100 274202
rect 15510 274030 15970 274044
rect 17050 274044 17058 274112
rect 17092 274044 17100 274112
rect 16690 274030 16760 274040
rect 16900 274030 16970 274040
rect 17050 274030 17100 274044
rect 15430 274016 15471 274022
rect 14471 273982 14483 274016
rect 15459 273982 15471 274016
rect 14471 273976 15150 273982
rect 15220 273976 15360 273982
rect 15150 273960 15220 273970
rect 15430 273976 15471 273982
rect 15510 274020 16690 274030
rect 15360 273960 15430 273970
rect 14380 273886 14390 273954
rect 14424 273886 14430 273954
rect 15510 273954 15560 274020
rect 14380 273796 14430 273886
rect 14510 273880 14580 273890
rect 14471 273858 14510 273864
rect 14720 273880 14790 273890
rect 14580 273858 14720 273864
rect 15510 273886 15518 273954
rect 15552 273886 15560 273954
rect 14790 273858 15471 273864
rect 14471 273824 14483 273858
rect 15459 273824 15471 273858
rect 14471 273818 14510 273824
rect 14580 273818 14720 273824
rect 14510 273800 14580 273810
rect 14790 273818 15471 273824
rect 14720 273800 14790 273810
rect 14380 273728 14390 273796
rect 14424 273728 14430 273796
rect 15510 273796 15560 273886
rect 14380 273638 14430 273728
rect 15150 273720 15220 273730
rect 14471 273700 15150 273706
rect 15360 273720 15430 273730
rect 15220 273700 15360 273706
rect 15510 273728 15518 273796
rect 15552 273728 15560 273796
rect 15430 273700 15471 273706
rect 14471 273666 14483 273700
rect 15459 273666 15471 273700
rect 14471 273660 15150 273666
rect 15220 273660 15360 273666
rect 15150 273640 15220 273650
rect 15430 273660 15471 273666
rect 15360 273640 15430 273650
rect 14380 273570 14390 273638
rect 14424 273570 14430 273638
rect 15510 273638 15560 273728
rect 15920 274016 16690 274020
rect 16760 274016 16900 274030
rect 16970 274016 17100 274030
rect 15920 273982 16023 274016
rect 16999 273982 17100 274016
rect 15920 273970 16690 273982
rect 15920 273954 15970 273970
rect 15920 273886 15930 273954
rect 15964 273886 15970 273954
rect 16760 273970 16900 273982
rect 16690 273950 16760 273960
rect 16970 273970 17100 273982
rect 16900 273950 16970 273960
rect 17050 273954 17100 273970
rect 15920 273796 15970 273886
rect 16060 273880 16130 273890
rect 16011 273858 16060 273864
rect 16270 273880 16340 273890
rect 16130 273858 16270 273864
rect 17050 273886 17058 273954
rect 17092 273886 17100 273954
rect 16340 273858 17011 273864
rect 16011 273824 16023 273858
rect 16999 273824 17011 273858
rect 16011 273818 16060 273824
rect 16130 273818 16270 273824
rect 16060 273800 16130 273810
rect 16340 273818 17011 273824
rect 16270 273800 16340 273810
rect 15920 273728 15930 273796
rect 15964 273728 15970 273796
rect 17050 273796 17100 273886
rect 15920 273710 15970 273728
rect 16690 273720 16760 273730
rect 15920 273700 16690 273710
rect 16900 273720 16970 273730
rect 16760 273700 16900 273710
rect 17050 273728 17058 273796
rect 17092 273728 17100 273796
rect 17050 273710 17100 273728
rect 16970 273700 17100 273710
rect 15510 273570 15518 273638
rect 15552 273570 15560 273638
rect 13984 273534 14330 273550
rect 13984 273330 14288 273534
rect 13984 273060 14000 273330
rect 14270 273060 14288 273330
rect 13984 272280 14288 273060
rect 13984 272010 14000 272280
rect 14270 272010 14288 272280
rect 13984 271778 14288 272010
rect 14322 271778 14330 273534
rect 13984 271760 14330 271778
rect 14380 273480 14430 273570
rect 14510 273560 14580 273570
rect 14471 273542 14510 273548
rect 14720 273560 14790 273570
rect 14580 273542 14720 273548
rect 14790 273542 15471 273548
rect 14471 273508 14483 273542
rect 15459 273508 15471 273542
rect 14471 273502 14510 273508
rect 14580 273502 14720 273508
rect 14510 273480 14580 273490
rect 14790 273502 15471 273508
rect 14720 273480 14790 273490
rect 15510 273480 15560 273570
rect 15614 273680 15866 273692
rect 15614 273550 15620 273680
rect 14380 273412 14390 273480
rect 14424 273412 14430 273480
rect 14380 273322 14430 273412
rect 15510 273412 15518 273480
rect 15552 273412 15560 273480
rect 15150 273400 15220 273410
rect 14471 273384 15150 273390
rect 15360 273400 15430 273410
rect 15220 273384 15360 273390
rect 15430 273384 15471 273390
rect 14471 273350 14483 273384
rect 15459 273350 15471 273384
rect 14471 273344 15150 273350
rect 14380 273254 14390 273322
rect 14424 273254 14430 273322
rect 15220 273344 15360 273350
rect 15150 273320 15220 273330
rect 15430 273344 15471 273350
rect 15360 273320 15430 273330
rect 15510 273322 15560 273412
rect 14380 273164 14430 273254
rect 14510 273250 14580 273260
rect 14471 273226 14510 273232
rect 14720 273250 14790 273260
rect 14580 273226 14720 273232
rect 15510 273254 15518 273322
rect 15552 273254 15560 273322
rect 15610 273540 15620 273550
rect 15860 273550 15866 273680
rect 15920 273666 16023 273700
rect 16999 273666 17100 273700
rect 15920 273650 16690 273666
rect 16760 273650 16900 273666
rect 16970 273650 17100 273666
rect 15920 273638 15970 273650
rect 16690 273640 16760 273650
rect 16900 273640 16970 273650
rect 15920 273570 15930 273638
rect 15964 273570 15970 273638
rect 17050 273638 17100 273650
rect 17050 273570 17058 273638
rect 17092 273570 17100 273638
rect 15860 273540 15870 273550
rect 15610 273270 15620 273280
rect 14790 273226 15471 273232
rect 14471 273192 14483 273226
rect 15459 273192 15471 273226
rect 14471 273186 14510 273192
rect 14580 273186 14720 273192
rect 14510 273170 14580 273180
rect 14790 273186 15471 273192
rect 14720 273170 14790 273180
rect 14380 273096 14390 273164
rect 14424 273096 14430 273164
rect 15510 273164 15560 273254
rect 14380 273006 14430 273096
rect 15150 273090 15220 273100
rect 14471 273068 15150 273074
rect 15360 273090 15430 273100
rect 15220 273068 15360 273074
rect 15510 273096 15518 273164
rect 15552 273096 15560 273164
rect 15614 273110 15620 273270
rect 15860 273270 15870 273280
rect 15920 273480 15970 273570
rect 16060 273560 16130 273570
rect 16011 273542 16060 273548
rect 16270 273560 16340 273570
rect 16130 273542 16270 273548
rect 16340 273542 17011 273548
rect 16011 273508 16023 273542
rect 16999 273508 17011 273542
rect 16011 273502 16060 273508
rect 16130 273502 16270 273508
rect 16060 273480 16130 273490
rect 16340 273502 17011 273508
rect 16270 273480 16340 273490
rect 17050 273480 17100 273570
rect 15920 273412 15930 273480
rect 15964 273412 15970 273480
rect 15920 273322 15970 273412
rect 17050 273412 17058 273480
rect 17092 273412 17100 273480
rect 17990 273430 18170 275100
rect 20540 275030 20590 275040
rect 21650 275030 21700 275040
rect 22060 275030 22110 275040
rect 23170 275030 23220 275040
rect 20510 275020 20620 275030
rect 20510 274900 20620 274910
rect 21620 275020 21730 275030
rect 21620 274900 21730 274910
rect 22030 275020 22140 275030
rect 22030 274900 22140 274910
rect 23140 275020 23250 275030
rect 23140 274900 23250 274910
rect 20540 274780 20590 274900
rect 21650 274780 21700 274900
rect 22060 274780 22110 274900
rect 23170 274780 23220 274900
rect 20510 274770 20620 274780
rect 20510 274650 20620 274660
rect 21620 274770 21730 274780
rect 21620 274650 21730 274660
rect 22030 274770 22140 274780
rect 22030 274650 22140 274660
rect 23140 274770 23250 274780
rect 23140 274650 23250 274660
rect 20540 274158 20590 274650
rect 20660 274240 20730 274250
rect 20620 274220 20660 274226
rect 20840 274240 20910 274250
rect 20730 274220 20840 274226
rect 20910 274220 21620 274226
rect 20620 274186 20632 274220
rect 21608 274186 21620 274220
rect 20620 274180 20660 274186
rect 20730 274180 20840 274186
rect 20660 274160 20730 274170
rect 20910 274180 21620 274186
rect 20840 274160 20910 274170
rect 20540 273990 20548 274158
rect 20582 273990 20590 274158
rect 21650 274158 21700 274650
rect 21650 273990 21658 274158
rect 21692 273990 21700 274158
rect 20540 273900 20590 273990
rect 21330 273980 21400 273990
rect 20620 273962 21330 273968
rect 21510 273980 21580 273990
rect 21400 273962 21510 273968
rect 21580 273962 21620 273968
rect 20620 273928 20632 273962
rect 21608 273928 21620 273962
rect 20620 273922 21330 273928
rect 21400 273922 21510 273928
rect 21330 273900 21400 273910
rect 21580 273922 21620 273928
rect 21510 273900 21580 273910
rect 21650 273900 21700 273990
rect 20540 273732 20548 273900
rect 20582 273732 20590 273900
rect 20540 273642 20590 273732
rect 21650 273732 21658 273900
rect 21692 273732 21700 273900
rect 20660 273720 20730 273730
rect 20620 273704 20660 273710
rect 20840 273720 20910 273730
rect 20730 273704 20840 273710
rect 20910 273704 21620 273710
rect 20620 273670 20632 273704
rect 21608 273670 21620 273704
rect 20620 273664 20660 273670
rect 20440 273477 20486 273489
rect 16690 273400 16760 273410
rect 16011 273384 16690 273390
rect 16900 273400 16970 273410
rect 16760 273384 16900 273390
rect 16970 273384 17011 273390
rect 16011 273350 16023 273384
rect 16999 273350 17011 273384
rect 16011 273344 16690 273350
rect 15860 273110 15866 273270
rect 15614 273098 15866 273110
rect 15920 273254 15930 273322
rect 15964 273254 15970 273322
rect 16760 273344 16900 273350
rect 16690 273320 16760 273330
rect 16970 273344 17011 273350
rect 16900 273320 16970 273330
rect 17050 273322 17100 273412
rect 15920 273164 15970 273254
rect 17050 273254 17058 273322
rect 17092 273254 17100 273322
rect 16060 273240 16130 273250
rect 16011 273226 16060 273232
rect 16270 273240 16340 273250
rect 16130 273226 16270 273232
rect 16340 273226 17011 273232
rect 16011 273192 16023 273226
rect 16999 273192 17011 273226
rect 16011 273186 16060 273192
rect 15430 273068 15471 273074
rect 14471 273034 14483 273068
rect 15459 273034 15471 273068
rect 14471 273028 15150 273034
rect 15220 273028 15360 273034
rect 15150 273010 15220 273020
rect 15430 273028 15471 273034
rect 15360 273010 15430 273020
rect 14380 272938 14390 273006
rect 14424 272938 14430 273006
rect 15510 273006 15560 273096
rect 14380 272848 14430 272938
rect 14510 272930 14580 272940
rect 14471 272910 14510 272916
rect 14720 272930 14790 272940
rect 14580 272910 14720 272916
rect 15510 272938 15518 273006
rect 15552 272938 15560 273006
rect 14790 272910 15471 272916
rect 14471 272876 14483 272910
rect 15459 272876 15471 272910
rect 14471 272870 14510 272876
rect 14580 272870 14720 272876
rect 14510 272850 14580 272860
rect 14790 272870 15471 272876
rect 14720 272850 14790 272860
rect 14380 272780 14390 272848
rect 14424 272780 14430 272848
rect 15510 272848 15560 272938
rect 15510 272780 15518 272848
rect 15552 272790 15560 272848
rect 15920 273096 15930 273164
rect 15964 273096 15970 273164
rect 16130 273186 16270 273192
rect 16060 273160 16130 273170
rect 16340 273186 17011 273192
rect 16270 273160 16340 273170
rect 17050 273164 17100 273254
rect 15920 273006 15970 273096
rect 16690 273090 16760 273100
rect 16011 273068 16690 273074
rect 16900 273090 16970 273100
rect 16760 273068 16900 273074
rect 17050 273096 17058 273164
rect 17092 273096 17100 273164
rect 16970 273068 17011 273074
rect 16011 273034 16023 273068
rect 16999 273034 17011 273068
rect 16011 273028 16690 273034
rect 16760 273028 16900 273034
rect 16690 273010 16760 273020
rect 16970 273028 17011 273034
rect 16900 273010 16970 273020
rect 15920 272938 15930 273006
rect 15964 272938 15970 273006
rect 17050 273006 17100 273096
rect 15920 272848 15970 272938
rect 16060 272930 16130 272940
rect 16011 272910 16060 272916
rect 16270 272930 16340 272940
rect 16130 272910 16270 272916
rect 17050 272938 17058 273006
rect 17092 272938 17100 273006
rect 17500 273350 18660 273430
rect 17500 273159 17550 273350
rect 18180 273240 18250 273250
rect 17579 273221 18180 273227
rect 18470 273240 18540 273250
rect 18250 273221 18470 273227
rect 18540 273221 18579 273227
rect 17579 273187 17591 273221
rect 18567 273187 18579 273221
rect 17579 273181 18180 273187
rect 18250 273181 18470 273187
rect 18180 273160 18250 273170
rect 18540 273181 18579 273187
rect 18470 273160 18540 273170
rect 17500 273091 17507 273159
rect 17541 273091 17550 273159
rect 17500 273001 17550 273091
rect 18610 273159 18660 273350
rect 18610 273091 18617 273159
rect 18651 273091 18660 273159
rect 17620 273080 17690 273090
rect 17579 273063 17620 273069
rect 17910 273080 17980 273090
rect 17690 273063 17910 273069
rect 17980 273063 18579 273069
rect 17579 273029 17591 273063
rect 18567 273029 18579 273063
rect 17579 273023 17620 273029
rect 16340 272910 17011 272916
rect 16011 272876 16023 272910
rect 16999 272876 17011 272910
rect 16011 272870 16060 272876
rect 16130 272870 16270 272876
rect 16060 272850 16130 272860
rect 16340 272870 17011 272876
rect 16270 272850 16340 272860
rect 15920 272790 15930 272848
rect 15552 272780 15930 272790
rect 15964 272780 15970 272848
rect 17050 272848 17100 272938
rect 17050 272780 17058 272848
rect 17092 272780 17100 272848
rect 14380 272690 14430 272780
rect 15150 272770 15220 272780
rect 14471 272752 15150 272758
rect 15360 272770 15430 272780
rect 15220 272752 15360 272758
rect 15430 272752 15471 272758
rect 14471 272718 14483 272752
rect 15459 272718 15471 272752
rect 14471 272712 15150 272718
rect 15220 272712 15360 272718
rect 15150 272690 15220 272700
rect 15430 272712 15471 272718
rect 15360 272690 15430 272700
rect 15510 272690 15970 272780
rect 16690 272770 16760 272780
rect 16011 272752 16690 272758
rect 16900 272770 16970 272780
rect 16760 272752 16900 272758
rect 16970 272752 17011 272758
rect 16011 272718 16023 272752
rect 16999 272718 17011 272752
rect 16011 272712 16690 272718
rect 16760 272712 16900 272718
rect 16690 272690 16760 272700
rect 16970 272712 17011 272718
rect 16900 272690 16970 272700
rect 17050 272690 17100 272780
rect 14380 272622 14390 272690
rect 14424 272622 14430 272690
rect 14380 272532 14430 272622
rect 15510 272622 15518 272690
rect 15552 272622 15930 272690
rect 15964 272622 15970 272690
rect 14510 272610 14580 272620
rect 14471 272594 14510 272600
rect 14720 272610 14790 272620
rect 14580 272594 14720 272600
rect 14790 272594 15471 272600
rect 14471 272560 14483 272594
rect 15459 272560 15471 272594
rect 14471 272554 14510 272560
rect 14380 272464 14390 272532
rect 14424 272464 14430 272532
rect 14580 272554 14720 272560
rect 14510 272530 14580 272540
rect 14790 272554 15471 272560
rect 14720 272530 14790 272540
rect 15510 272532 15970 272622
rect 17050 272622 17058 272690
rect 17092 272622 17100 272690
rect 16060 272610 16130 272620
rect 16011 272594 16060 272600
rect 16270 272610 16340 272620
rect 16130 272594 16270 272600
rect 16340 272594 17011 272600
rect 16011 272560 16023 272594
rect 16999 272560 17011 272594
rect 16011 272554 16060 272560
rect 14380 272374 14430 272464
rect 15150 272460 15220 272470
rect 14471 272436 15150 272442
rect 15360 272460 15430 272470
rect 15220 272436 15360 272442
rect 15510 272464 15518 272532
rect 15552 272520 15930 272532
rect 15552 272464 15560 272520
rect 15430 272436 15471 272442
rect 14471 272402 14483 272436
rect 15459 272402 15471 272436
rect 14471 272396 15150 272402
rect 15220 272396 15360 272402
rect 15150 272380 15220 272390
rect 15430 272396 15471 272402
rect 15360 272380 15430 272390
rect 14380 272306 14390 272374
rect 14424 272306 14430 272374
rect 15510 272374 15560 272464
rect 14380 272216 14430 272306
rect 14510 272300 14580 272310
rect 14471 272278 14510 272284
rect 14720 272300 14790 272310
rect 14580 272278 14720 272284
rect 15510 272306 15518 272374
rect 15552 272306 15560 272374
rect 14790 272278 15471 272284
rect 14471 272244 14483 272278
rect 15459 272244 15471 272278
rect 14471 272238 14510 272244
rect 14580 272238 14720 272244
rect 14510 272220 14580 272230
rect 14790 272238 15471 272244
rect 14720 272220 14790 272230
rect 14380 272148 14390 272216
rect 14424 272148 14430 272216
rect 15510 272216 15560 272306
rect 15920 272464 15930 272520
rect 15964 272464 15970 272532
rect 16130 272554 16270 272560
rect 16060 272530 16130 272540
rect 16340 272554 17011 272560
rect 16270 272530 16340 272540
rect 17050 272532 17100 272622
rect 15920 272374 15970 272464
rect 17050 272464 17058 272532
rect 17092 272464 17100 272532
rect 16690 272450 16760 272460
rect 16011 272436 16690 272442
rect 16900 272450 16970 272460
rect 16760 272436 16900 272442
rect 16970 272436 17011 272442
rect 16011 272402 16023 272436
rect 16999 272402 17011 272436
rect 16011 272396 16690 272402
rect 15920 272306 15930 272374
rect 15964 272306 15970 272374
rect 16760 272396 16900 272402
rect 16690 272370 16760 272380
rect 16970 272396 17011 272402
rect 16900 272370 16970 272380
rect 17050 272374 17100 272464
rect 14380 272058 14430 272148
rect 15150 272140 15220 272150
rect 14471 272120 15150 272126
rect 15360 272140 15430 272150
rect 15220 272120 15360 272126
rect 15510 272148 15518 272216
rect 15552 272148 15560 272216
rect 15430 272120 15471 272126
rect 14471 272086 14483 272120
rect 15459 272086 15471 272120
rect 14471 272080 15150 272086
rect 15220 272080 15360 272086
rect 15150 272060 15220 272070
rect 15430 272080 15471 272086
rect 15360 272060 15430 272070
rect 14380 271990 14390 272058
rect 14424 271990 14430 272058
rect 15510 272058 15560 272148
rect 15510 271990 15518 272058
rect 15552 271990 15560 272058
rect 15614 272210 15866 272222
rect 15614 272050 15620 272210
rect 14380 271900 14430 271990
rect 14510 271980 14580 271990
rect 14471 271962 14510 271968
rect 14720 271980 14790 271990
rect 14580 271962 14720 271968
rect 14790 271962 15471 271968
rect 14471 271928 14483 271962
rect 15459 271928 15471 271962
rect 14471 271922 14510 271928
rect 14580 271922 14720 271928
rect 14510 271900 14580 271910
rect 14790 271922 15471 271928
rect 14720 271900 14790 271910
rect 15510 271900 15560 271990
rect 14380 271832 14390 271900
rect 14424 271832 14430 271900
rect 13984 271029 13990 271760
rect 13944 271017 13990 271029
rect 14380 271742 14430 271832
rect 15510 271832 15518 271900
rect 15552 271832 15560 271900
rect 15150 271820 15220 271830
rect 14471 271804 15150 271810
rect 15360 271820 15430 271830
rect 15220 271804 15360 271810
rect 15430 271804 15471 271810
rect 14471 271770 14483 271804
rect 15459 271770 15471 271804
rect 14471 271764 15150 271770
rect 14380 271674 14390 271742
rect 14424 271674 14430 271742
rect 15220 271764 15360 271770
rect 15150 271740 15220 271750
rect 15430 271764 15471 271770
rect 15360 271740 15430 271750
rect 15510 271742 15560 271832
rect 15610 272040 15620 272050
rect 15860 272050 15866 272210
rect 15920 272216 15970 272306
rect 16060 272300 16130 272310
rect 16011 272278 16060 272284
rect 16270 272300 16340 272310
rect 16130 272278 16270 272284
rect 17050 272306 17058 272374
rect 17092 272306 17100 272374
rect 17399 272976 17445 272988
rect 17399 272326 17405 272976
rect 17439 272326 17445 272976
rect 17399 272314 17445 272326
rect 17500 272933 17507 273001
rect 17541 272933 17550 273001
rect 17690 273023 17910 273029
rect 17620 273000 17690 273010
rect 17980 273023 18579 273029
rect 17910 273000 17980 273010
rect 18610 273001 18660 273091
rect 17500 272843 17550 272933
rect 18610 272933 18617 273001
rect 18651 272933 18660 273001
rect 19020 273350 20180 273430
rect 19020 273159 19070 273350
rect 19700 273240 19770 273250
rect 19099 273221 19700 273227
rect 19990 273240 20060 273250
rect 19770 273221 19990 273227
rect 20060 273221 20099 273227
rect 19099 273187 19111 273221
rect 20087 273187 20099 273221
rect 19099 273181 19700 273187
rect 19770 273181 19990 273187
rect 19700 273160 19770 273170
rect 20060 273181 20099 273187
rect 19990 273160 20060 273170
rect 19020 273091 19027 273159
rect 19061 273091 19070 273159
rect 19020 273001 19070 273091
rect 20130 273159 20180 273350
rect 20130 273091 20137 273159
rect 20171 273091 20180 273159
rect 19140 273080 19210 273090
rect 19099 273063 19140 273069
rect 19430 273080 19500 273090
rect 19210 273063 19430 273069
rect 19500 273063 20099 273069
rect 19099 273029 19111 273063
rect 20087 273029 20099 273063
rect 19099 273023 19140 273029
rect 18180 272920 18250 272930
rect 17579 272905 18180 272911
rect 18470 272920 18540 272930
rect 18250 272905 18470 272911
rect 18540 272905 18579 272911
rect 17579 272871 17591 272905
rect 18567 272871 18579 272905
rect 17579 272865 18180 272871
rect 17500 272775 17507 272843
rect 17541 272775 17550 272843
rect 18250 272865 18470 272871
rect 18180 272840 18250 272850
rect 18540 272865 18579 272871
rect 18470 272840 18540 272850
rect 18610 272843 18660 272933
rect 17500 272685 17550 272775
rect 18610 272775 18617 272843
rect 18651 272775 18660 272843
rect 18713 272976 18759 272988
rect 18713 272790 18719 272976
rect 17620 272760 17690 272770
rect 17579 272747 17620 272753
rect 17910 272760 17980 272770
rect 17690 272747 17910 272753
rect 17980 272747 18579 272753
rect 17579 272713 17591 272747
rect 18567 272713 18579 272747
rect 17579 272707 17620 272713
rect 17500 272617 17507 272685
rect 17541 272617 17550 272685
rect 17690 272707 17910 272713
rect 17620 272680 17690 272690
rect 17980 272707 18579 272713
rect 17910 272680 17980 272690
rect 18610 272685 18660 272775
rect 17500 272527 17550 272617
rect 18610 272617 18617 272685
rect 18651 272617 18660 272685
rect 18180 272600 18250 272610
rect 17579 272589 18180 272595
rect 18470 272600 18540 272610
rect 18250 272589 18470 272595
rect 18540 272589 18579 272595
rect 17579 272555 17591 272589
rect 18567 272555 18579 272589
rect 17579 272549 18180 272555
rect 17500 272459 17507 272527
rect 17541 272459 17550 272527
rect 18250 272549 18470 272555
rect 18180 272520 18250 272530
rect 18540 272549 18579 272555
rect 18470 272520 18540 272530
rect 18610 272527 18660 272617
rect 17500 272369 17550 272459
rect 17620 272450 17690 272460
rect 17579 272431 17620 272437
rect 17910 272450 17980 272460
rect 17690 272431 17910 272437
rect 18610 272459 18617 272527
rect 18651 272459 18660 272527
rect 18710 272780 18719 272790
rect 18753 272790 18759 272976
rect 18919 272976 18965 272988
rect 18919 272790 18925 272976
rect 18753 272780 18925 272790
rect 18959 272790 18965 272976
rect 19020 272933 19027 273001
rect 19061 272933 19070 273001
rect 19210 273023 19430 273029
rect 19140 273000 19210 273010
rect 19500 273023 20099 273029
rect 19430 273000 19500 273010
rect 20130 273001 20180 273091
rect 19020 272843 19070 272933
rect 20130 272933 20137 273001
rect 20171 272933 20180 273001
rect 19700 272920 19770 272930
rect 19099 272905 19700 272911
rect 19990 272920 20060 272930
rect 19770 272905 19990 272911
rect 20060 272905 20099 272911
rect 19099 272871 19111 272905
rect 20087 272871 20099 272905
rect 19099 272865 19700 272871
rect 18959 272780 18970 272790
rect 18710 272510 18719 272520
rect 17980 272431 18579 272437
rect 17579 272397 17591 272431
rect 18567 272397 18579 272431
rect 17579 272391 17620 272397
rect 17690 272391 17910 272397
rect 17620 272370 17690 272380
rect 17980 272391 18579 272397
rect 17910 272370 17980 272380
rect 16340 272278 17011 272284
rect 16011 272244 16023 272278
rect 16999 272244 17011 272278
rect 16011 272238 16060 272244
rect 16130 272238 16270 272244
rect 16060 272220 16130 272230
rect 16340 272238 17011 272244
rect 16270 272220 16340 272230
rect 15920 272148 15930 272216
rect 15964 272148 15970 272216
rect 17050 272216 17100 272306
rect 15920 272058 15970 272148
rect 16690 272140 16760 272150
rect 16011 272120 16690 272126
rect 16900 272140 16970 272150
rect 16760 272120 16900 272126
rect 17050 272148 17058 272216
rect 17092 272148 17100 272216
rect 16970 272120 17011 272126
rect 16011 272086 16023 272120
rect 16999 272086 17011 272120
rect 16011 272080 16690 272086
rect 16760 272080 16900 272086
rect 16690 272060 16760 272070
rect 16970 272080 17011 272086
rect 16900 272060 16970 272070
rect 15860 272040 15870 272050
rect 15610 271770 15620 271780
rect 14380 271584 14430 271674
rect 15510 271674 15518 271742
rect 15552 271674 15560 271742
rect 14510 271660 14580 271670
rect 14471 271646 14510 271652
rect 14720 271660 14790 271670
rect 14580 271646 14720 271652
rect 14790 271646 15471 271652
rect 14471 271612 14483 271646
rect 15459 271612 15471 271646
rect 14471 271606 14510 271612
rect 14380 271516 14390 271584
rect 14424 271516 14430 271584
rect 14580 271606 14720 271612
rect 14510 271580 14580 271590
rect 14790 271606 15471 271612
rect 14720 271580 14790 271590
rect 15510 271584 15560 271674
rect 15614 271640 15620 271770
rect 15860 271770 15870 271780
rect 15920 271990 15930 272058
rect 15964 271990 15970 272058
rect 17050 272058 17100 272148
rect 17050 271990 17058 272058
rect 17092 271990 17100 272058
rect 15920 271900 15970 271990
rect 16060 271980 16130 271990
rect 16011 271962 16060 271968
rect 16270 271980 16340 271990
rect 16130 271962 16270 271968
rect 16340 271962 17011 271968
rect 16011 271928 16023 271962
rect 16999 271928 17011 271962
rect 16011 271922 16060 271928
rect 16130 271922 16270 271928
rect 16060 271900 16130 271910
rect 16340 271922 17011 271928
rect 16270 271900 16340 271910
rect 17050 271900 17100 271990
rect 15920 271832 15930 271900
rect 15964 271832 15970 271900
rect 15920 271820 15970 271832
rect 17050 271832 17058 271900
rect 17092 271832 17100 271900
rect 17500 272301 17507 272369
rect 17541 272301 17550 272369
rect 17500 272211 17550 272301
rect 18610 272369 18660 272459
rect 18610 272301 18617 272369
rect 18651 272301 18660 272369
rect 18713 272326 18719 272510
rect 18753 272510 18925 272520
rect 18753 272326 18759 272510
rect 18713 272314 18759 272326
rect 18919 272326 18925 272510
rect 18959 272510 18970 272520
rect 19020 272775 19027 272843
rect 19061 272775 19070 272843
rect 19770 272865 19990 272871
rect 19700 272840 19770 272850
rect 20060 272865 20099 272871
rect 19990 272840 20060 272850
rect 20130 272843 20180 272933
rect 19020 272685 19070 272775
rect 20130 272775 20137 272843
rect 20171 272775 20180 272843
rect 20233 272976 20279 272988
rect 20233 272790 20239 272976
rect 19140 272760 19210 272770
rect 19099 272747 19140 272753
rect 19430 272760 19500 272770
rect 19210 272747 19430 272753
rect 19500 272747 20099 272753
rect 19099 272713 19111 272747
rect 20087 272713 20099 272747
rect 19099 272707 19140 272713
rect 19020 272617 19027 272685
rect 19061 272617 19070 272685
rect 19210 272707 19430 272713
rect 19140 272680 19210 272690
rect 19500 272707 20099 272713
rect 19430 272680 19500 272690
rect 20130 272685 20180 272775
rect 19020 272527 19070 272617
rect 20130 272617 20137 272685
rect 20171 272617 20180 272685
rect 19700 272600 19770 272610
rect 19099 272589 19700 272595
rect 19990 272600 20060 272610
rect 19770 272589 19990 272595
rect 20060 272589 20099 272595
rect 19099 272555 19111 272589
rect 20087 272555 20099 272589
rect 19099 272549 19700 272555
rect 18959 272326 18965 272510
rect 18919 272314 18965 272326
rect 19020 272459 19027 272527
rect 19061 272459 19070 272527
rect 19770 272549 19990 272555
rect 19700 272520 19770 272530
rect 20060 272549 20099 272555
rect 19990 272520 20060 272530
rect 20130 272527 20180 272617
rect 19020 272369 19070 272459
rect 19140 272450 19210 272460
rect 19099 272431 19140 272437
rect 19430 272450 19500 272460
rect 19210 272431 19430 272437
rect 20130 272459 20137 272527
rect 20171 272459 20180 272527
rect 20230 272780 20239 272790
rect 20273 272790 20279 272976
rect 20440 272790 20446 273477
rect 20273 272780 20446 272790
rect 20480 272790 20486 273477
rect 20540 273474 20548 273642
rect 20582 273474 20590 273642
rect 20730 273664 20840 273670
rect 20660 273640 20730 273650
rect 20910 273664 21620 273670
rect 20840 273640 20910 273650
rect 21650 273642 21700 273732
rect 20540 273384 20590 273474
rect 21650 273474 21658 273642
rect 21692 273474 21700 273642
rect 22060 274414 22110 274650
rect 22180 274490 22250 274500
rect 22140 274476 22180 274482
rect 22360 274490 22430 274500
rect 22250 274476 22360 274482
rect 22430 274476 23140 274482
rect 22140 274442 22152 274476
rect 23128 274442 23140 274476
rect 22140 274436 22180 274442
rect 22060 274246 22068 274414
rect 22102 274246 22110 274414
rect 22250 274436 22360 274442
rect 22180 274410 22250 274420
rect 22430 274436 23140 274442
rect 22360 274410 22430 274420
rect 23170 274414 23220 274650
rect 22060 274156 22110 274246
rect 23170 274246 23178 274414
rect 23212 274246 23220 274414
rect 22850 274230 22920 274240
rect 22140 274218 22850 274224
rect 23030 274230 23100 274240
rect 22920 274218 23030 274224
rect 23100 274218 23140 274224
rect 22140 274184 22152 274218
rect 23128 274184 23140 274218
rect 22140 274178 22850 274184
rect 22060 273988 22068 274156
rect 22102 273988 22110 274156
rect 22920 274178 23030 274184
rect 22850 274150 22920 274160
rect 23100 274178 23140 274184
rect 23030 274150 23100 274160
rect 23170 274156 23220 274246
rect 22060 273898 22110 273988
rect 22180 273980 22250 273990
rect 22140 273960 22180 273966
rect 22360 273980 22430 273990
rect 22250 273960 22360 273966
rect 23170 273988 23178 274156
rect 23212 273988 23220 274156
rect 22430 273960 23140 273966
rect 22140 273926 22152 273960
rect 23128 273926 23140 273960
rect 22140 273920 22180 273926
rect 22250 273920 22360 273926
rect 22180 273900 22250 273910
rect 22430 273920 23140 273926
rect 22360 273900 22430 273910
rect 22060 273730 22068 273898
rect 22102 273730 22110 273898
rect 23170 273898 23220 273988
rect 23170 273730 23178 273898
rect 23212 273730 23220 273898
rect 22060 273640 22110 273730
rect 22850 273720 22920 273730
rect 22140 273702 22850 273708
rect 23030 273720 23100 273730
rect 22920 273702 23030 273708
rect 23100 273702 23140 273708
rect 22140 273668 22152 273702
rect 23128 273668 23140 273702
rect 22140 273662 22850 273668
rect 22920 273662 23030 273668
rect 22850 273640 22920 273650
rect 23100 273662 23140 273668
rect 23030 273640 23100 273650
rect 23170 273640 23220 273730
rect 21960 273604 22006 273616
rect 21330 273460 21400 273470
rect 20620 273446 21330 273452
rect 21510 273460 21580 273470
rect 21400 273446 21510 273452
rect 21580 273446 21620 273452
rect 20620 273412 20632 273446
rect 21608 273412 21620 273446
rect 20620 273406 21330 273412
rect 20540 273216 20548 273384
rect 20582 273216 20590 273384
rect 21400 273406 21510 273412
rect 21330 273380 21400 273390
rect 21580 273406 21620 273412
rect 21510 273380 21580 273390
rect 21650 273384 21700 273474
rect 20540 273126 20590 273216
rect 21650 273216 21658 273384
rect 21692 273216 21700 273384
rect 20660 273200 20730 273210
rect 20620 273188 20660 273194
rect 20840 273200 20910 273210
rect 20730 273188 20840 273194
rect 20910 273188 21620 273194
rect 20620 273154 20632 273188
rect 21608 273154 21620 273188
rect 20620 273148 20660 273154
rect 20540 272958 20548 273126
rect 20582 272958 20590 273126
rect 20730 273148 20840 273154
rect 20660 273120 20730 273130
rect 20910 273148 21620 273154
rect 20840 273120 20910 273130
rect 21650 273126 21700 273216
rect 20540 272868 20590 272958
rect 21330 272950 21400 272960
rect 20620 272930 21330 272936
rect 21510 272950 21580 272960
rect 21400 272930 21510 272936
rect 21650 272958 21658 273126
rect 21692 272958 21700 273126
rect 21580 272930 21620 272936
rect 20620 272896 20632 272930
rect 21608 272896 21620 272930
rect 20620 272890 21330 272896
rect 21400 272890 21510 272896
rect 21330 272870 21400 272880
rect 21580 272890 21620 272896
rect 21510 272870 21580 272880
rect 20480 272780 20490 272790
rect 20230 272510 20239 272520
rect 19500 272431 20099 272437
rect 19099 272397 19111 272431
rect 20087 272397 20099 272431
rect 19099 272391 19140 272397
rect 19210 272391 19430 272397
rect 19140 272370 19210 272380
rect 19500 272391 20099 272397
rect 19430 272370 19500 272380
rect 18180 272290 18250 272300
rect 17579 272273 18180 272279
rect 18470 272290 18540 272300
rect 18250 272273 18470 272279
rect 18540 272273 18579 272279
rect 17579 272239 17591 272273
rect 18567 272239 18579 272273
rect 17579 272233 18180 272239
rect 17500 272143 17507 272211
rect 17541 272143 17550 272211
rect 18250 272233 18470 272239
rect 18180 272210 18250 272220
rect 18540 272233 18579 272239
rect 18470 272210 18540 272220
rect 18610 272211 18660 272301
rect 17500 271950 17550 272143
rect 18610 272143 18617 272211
rect 18651 272143 18660 272211
rect 17620 272130 17690 272140
rect 17579 272115 17620 272121
rect 17910 272130 17980 272140
rect 17690 272115 17910 272121
rect 17980 272115 18579 272121
rect 17579 272081 17591 272115
rect 18567 272081 18579 272115
rect 17579 272075 17620 272081
rect 17690 272075 17910 272081
rect 17620 272050 17690 272060
rect 17980 272075 18579 272081
rect 17910 272050 17980 272060
rect 18610 271950 18660 272143
rect 17500 271870 18660 271950
rect 19020 272301 19027 272369
rect 19061 272301 19070 272369
rect 19020 272211 19070 272301
rect 20130 272369 20180 272459
rect 20130 272301 20137 272369
rect 20171 272301 20180 272369
rect 20233 272326 20239 272510
rect 20273 272510 20446 272520
rect 20273 272326 20279 272510
rect 20233 272314 20279 272326
rect 19700 272290 19770 272300
rect 19099 272273 19700 272279
rect 19990 272290 20060 272300
rect 19770 272273 19990 272279
rect 20060 272273 20099 272279
rect 19099 272239 19111 272273
rect 20087 272239 20099 272273
rect 19099 272233 19700 272239
rect 19020 272143 19027 272211
rect 19061 272143 19070 272211
rect 19770 272233 19990 272239
rect 19700 272210 19770 272220
rect 20060 272233 20099 272239
rect 19990 272210 20060 272220
rect 20130 272211 20180 272301
rect 19020 271950 19070 272143
rect 20130 272143 20137 272211
rect 20171 272143 20180 272211
rect 19140 272130 19210 272140
rect 19099 272115 19140 272121
rect 19430 272130 19500 272140
rect 19210 272115 19430 272121
rect 19500 272115 20099 272121
rect 19099 272081 19111 272115
rect 20087 272081 20099 272115
rect 19099 272075 19140 272081
rect 19210 272075 19430 272081
rect 19140 272050 19210 272060
rect 19500 272075 20099 272081
rect 19430 272050 19500 272060
rect 20130 271950 20180 272143
rect 19020 271870 20180 271950
rect 16690 271820 16760 271830
rect 16900 271820 16970 271830
rect 17050 271820 17100 271832
rect 15920 271804 16690 271820
rect 16760 271804 16900 271820
rect 16970 271804 17100 271820
rect 15920 271770 16023 271804
rect 16999 271770 17100 271804
rect 15860 271640 15866 271770
rect 15614 271628 15866 271640
rect 15920 271760 16690 271770
rect 15920 271742 15970 271760
rect 15920 271674 15930 271742
rect 15964 271674 15970 271742
rect 16760 271760 16900 271770
rect 16690 271740 16760 271750
rect 16970 271760 17100 271770
rect 16900 271740 16970 271750
rect 17050 271742 17100 271760
rect 14380 271426 14430 271516
rect 15150 271510 15220 271520
rect 14471 271488 15150 271494
rect 15360 271510 15430 271520
rect 15220 271488 15360 271494
rect 15510 271516 15518 271584
rect 15552 271516 15560 271584
rect 15430 271488 15471 271494
rect 14471 271454 14483 271488
rect 15459 271454 15471 271488
rect 14471 271448 15150 271454
rect 15220 271448 15360 271454
rect 15150 271430 15220 271440
rect 15430 271448 15471 271454
rect 15360 271430 15430 271440
rect 14380 271358 14390 271426
rect 14424 271358 14430 271426
rect 15510 271426 15560 271516
rect 14380 271268 14430 271358
rect 14510 271350 14580 271360
rect 14471 271330 14510 271336
rect 14720 271350 14790 271360
rect 14580 271330 14720 271336
rect 15510 271358 15518 271426
rect 15552 271358 15560 271426
rect 14790 271330 15471 271336
rect 14471 271296 14483 271330
rect 15459 271296 15471 271330
rect 14471 271290 14510 271296
rect 14580 271290 14720 271296
rect 14510 271270 14580 271280
rect 14790 271290 15471 271296
rect 15510 271290 15560 271358
rect 15920 271584 15970 271674
rect 17050 271674 17058 271742
rect 17092 271674 17100 271742
rect 16060 271660 16130 271670
rect 16011 271646 16060 271652
rect 16270 271660 16340 271670
rect 16130 271646 16270 271652
rect 16340 271646 17011 271652
rect 16011 271612 16023 271646
rect 16999 271612 17011 271646
rect 16011 271606 16060 271612
rect 15920 271516 15930 271584
rect 15964 271516 15970 271584
rect 16130 271606 16270 271612
rect 16060 271580 16130 271590
rect 16340 271606 17011 271612
rect 16270 271580 16340 271590
rect 17050 271584 17100 271674
rect 15920 271500 15970 271516
rect 16690 271510 16760 271520
rect 15920 271488 16690 271500
rect 16900 271510 16970 271520
rect 16760 271488 16900 271500
rect 17050 271516 17058 271584
rect 17092 271516 17100 271584
rect 17050 271500 17100 271516
rect 16970 271488 17100 271500
rect 15920 271454 16023 271488
rect 16999 271454 17100 271488
rect 15920 271440 16690 271454
rect 16760 271440 16900 271454
rect 16970 271440 17100 271454
rect 15920 271426 15970 271440
rect 16690 271430 16760 271440
rect 16900 271430 16970 271440
rect 15920 271358 15930 271426
rect 15964 271358 15970 271426
rect 17050 271426 17100 271440
rect 15920 271290 15970 271358
rect 16060 271350 16130 271360
rect 16011 271330 16060 271336
rect 16270 271350 16340 271360
rect 16130 271330 16270 271336
rect 17050 271358 17058 271426
rect 17092 271358 17100 271426
rect 16340 271330 17011 271336
rect 16011 271296 16023 271330
rect 16999 271296 17011 271330
rect 16011 271290 16060 271296
rect 14720 271270 14790 271280
rect 14380 271200 14390 271268
rect 14424 271200 14430 271268
rect 15510 271268 15970 271290
rect 16130 271290 16270 271296
rect 16060 271270 16130 271280
rect 16340 271290 17011 271296
rect 16270 271270 16340 271280
rect 15510 271200 15518 271268
rect 15552 271200 15930 271268
rect 15964 271200 15970 271268
rect 17050 271268 17100 271358
rect 17050 271200 17058 271268
rect 17092 271200 17100 271268
rect 14380 271110 14430 271200
rect 15150 271190 15220 271200
rect 14471 271172 15150 271178
rect 15360 271190 15430 271200
rect 15220 271172 15360 271178
rect 15430 271172 15471 271178
rect 14471 271138 14483 271172
rect 15459 271138 15471 271172
rect 14471 271132 15150 271138
rect 15220 271132 15360 271138
rect 15150 271110 15220 271120
rect 15430 271132 15471 271138
rect 15360 271110 15430 271120
rect 15510 271110 15970 271200
rect 16690 271190 16760 271200
rect 16011 271172 16690 271178
rect 16900 271190 16970 271200
rect 16760 271172 16900 271178
rect 16970 271172 17011 271178
rect 16011 271138 16023 271172
rect 16999 271138 17011 271172
rect 16011 271132 16690 271138
rect 16760 271132 16900 271138
rect 16690 271110 16760 271120
rect 16970 271132 17011 271138
rect 16900 271110 16970 271120
rect 17050 271110 17100 271200
rect 14380 271042 14390 271110
rect 14424 271042 14430 271110
rect 13450 270950 13520 270960
rect 12801 270936 13450 270942
rect 13690 270950 13760 270960
rect 13520 270936 13690 270942
rect 13760 270936 13801 270942
rect 12801 270902 12813 270936
rect 13789 270902 13801 270936
rect 12801 270896 13450 270902
rect 12710 270806 12720 270874
rect 12754 270806 12760 270874
rect 13520 270896 13690 270902
rect 13450 270870 13520 270880
rect 13760 270896 13801 270902
rect 13690 270870 13760 270880
rect 13840 270874 13890 270964
rect 12710 270716 12760 270806
rect 13840 270806 13848 270874
rect 13882 270806 13890 270874
rect 14380 270910 14430 271042
rect 15510 271042 15518 271110
rect 15552 271042 15930 271110
rect 15964 271042 15970 271110
rect 14510 271030 14580 271040
rect 14471 271014 14510 271020
rect 14720 271030 14790 271040
rect 14580 271014 14720 271020
rect 15510 271020 15970 271042
rect 17050 271042 17058 271110
rect 17092 271042 17100 271110
rect 16060 271030 16130 271040
rect 14790 271014 15471 271020
rect 14471 270980 14483 271014
rect 15459 270980 15471 271014
rect 14471 270974 14510 270980
rect 14580 270974 14720 270980
rect 14510 270950 14580 270960
rect 14790 270974 15471 270980
rect 14720 270950 14790 270960
rect 15510 270910 15560 271020
rect 16011 271014 16060 271020
rect 16270 271030 16340 271040
rect 16130 271014 16270 271020
rect 17050 271020 17100 271042
rect 16340 271014 17011 271020
rect 16011 270980 16023 271014
rect 16999 270980 17011 271014
rect 16011 270974 16060 270980
rect 16130 270974 16270 270980
rect 16060 270950 16130 270960
rect 16340 270974 17011 270980
rect 16270 270950 16340 270960
rect 14380 270830 15560 270910
rect 12840 270790 12910 270800
rect 12801 270778 12840 270784
rect 13080 270790 13150 270800
rect 12910 270778 13080 270784
rect 13150 270778 13801 270784
rect 12801 270744 12813 270778
rect 13789 270744 13801 270778
rect 12801 270738 12840 270744
rect 12710 270648 12720 270716
rect 12754 270648 12760 270716
rect 12910 270738 13080 270744
rect 12840 270710 12910 270720
rect 13150 270738 13801 270744
rect 13080 270710 13150 270720
rect 13840 270716 13890 270806
rect 12710 270558 12760 270648
rect 13450 270640 13520 270650
rect 12801 270620 13450 270626
rect 13690 270640 13760 270650
rect 13520 270620 13690 270626
rect 13840 270648 13848 270716
rect 13882 270700 13890 270716
rect 13882 270660 13950 270700
rect 13760 270620 13801 270626
rect 12801 270586 12813 270620
rect 13789 270586 13801 270620
rect 12801 270580 13450 270586
rect 13520 270580 13690 270586
rect 13450 270560 13520 270570
rect 13760 270580 13801 270586
rect 13840 270580 13860 270648
rect 13940 270580 13950 270660
rect 13690 270560 13760 270570
rect 12710 270490 12720 270558
rect 12754 270490 12760 270558
rect 13840 270558 13950 270580
rect 13840 270490 13848 270558
rect 13882 270540 13950 270558
rect 13882 270490 13890 270540
rect 12710 270400 12760 270490
rect 12840 270480 12910 270490
rect 12801 270462 12840 270468
rect 13080 270480 13150 270490
rect 12910 270462 13080 270468
rect 13150 270462 13801 270468
rect 12801 270428 12813 270462
rect 13789 270428 13801 270462
rect 12801 270422 12840 270428
rect 12910 270422 13080 270428
rect 12840 270400 12910 270410
rect 13150 270422 13801 270428
rect 13080 270400 13150 270410
rect 13840 270400 13890 270490
rect 12710 270332 12720 270400
rect 12754 270332 12760 270400
rect 12710 270242 12760 270332
rect 13840 270332 13848 270400
rect 13882 270332 13890 270400
rect 13450 270320 13520 270330
rect 12801 270304 13450 270310
rect 13690 270320 13760 270330
rect 13520 270304 13690 270310
rect 13760 270304 13801 270310
rect 12801 270270 12813 270304
rect 13789 270270 13801 270304
rect 12801 270264 13450 270270
rect 12710 270174 12720 270242
rect 12754 270174 12760 270242
rect 13520 270264 13690 270270
rect 13450 270240 13520 270250
rect 13760 270264 13801 270270
rect 13690 270240 13760 270250
rect 13840 270242 13890 270332
rect 12710 270084 12760 270174
rect 13840 270174 13848 270242
rect 13882 270174 13890 270242
rect 19510 270200 19690 271870
rect 20440 271833 20446 272510
rect 20480 272510 20490 272520
rect 20540 272700 20548 272868
rect 20582 272700 20590 272868
rect 21650 272868 21700 272958
rect 21650 272700 21658 272868
rect 21692 272700 21700 272868
rect 21754 273477 21800 273489
rect 21754 272790 21760 273477
rect 20540 272610 20590 272700
rect 20660 272690 20730 272700
rect 20620 272672 20660 272678
rect 20840 272690 20910 272700
rect 20730 272672 20840 272678
rect 20910 272672 21620 272678
rect 20620 272638 20632 272672
rect 21608 272638 21620 272672
rect 20620 272632 20660 272638
rect 20730 272632 20840 272638
rect 20660 272610 20730 272620
rect 20910 272632 21620 272638
rect 20840 272610 20910 272620
rect 21650 272610 21700 272700
rect 20480 271833 20486 272510
rect 20440 271821 20486 271833
rect 20540 272442 20548 272610
rect 20582 272442 20590 272610
rect 20540 272352 20590 272442
rect 21650 272442 21658 272610
rect 21692 272442 21700 272610
rect 21750 272780 21760 272790
rect 21794 272790 21800 273477
rect 21960 272790 21966 273604
rect 21794 272780 21966 272790
rect 22000 272790 22006 273604
rect 22060 273472 22068 273640
rect 22102 273472 22110 273640
rect 22060 273382 22110 273472
rect 23170 273472 23178 273640
rect 23212 273472 23220 273640
rect 24090 273630 25270 273700
rect 22180 273460 22250 273470
rect 22140 273444 22180 273450
rect 22360 273460 22430 273470
rect 22250 273444 22360 273450
rect 22430 273444 23140 273450
rect 22140 273410 22152 273444
rect 23128 273410 23140 273444
rect 22140 273404 22180 273410
rect 22060 273214 22068 273382
rect 22102 273214 22110 273382
rect 22250 273404 22360 273410
rect 22180 273380 22250 273390
rect 22430 273404 23140 273410
rect 22360 273380 22430 273390
rect 23170 273382 23220 273472
rect 22060 273124 22110 273214
rect 23170 273214 23178 273382
rect 23212 273214 23220 273382
rect 22850 273200 22920 273210
rect 22140 273186 22850 273192
rect 23030 273200 23100 273210
rect 22920 273186 23030 273192
rect 23100 273186 23140 273192
rect 22140 273152 22152 273186
rect 23128 273152 23140 273186
rect 22140 273146 22850 273152
rect 22060 272956 22068 273124
rect 22102 272956 22110 273124
rect 22920 273146 23030 273152
rect 22850 273120 22920 273130
rect 23100 273146 23140 273152
rect 23030 273120 23100 273130
rect 23170 273124 23220 273214
rect 22060 272866 22110 272956
rect 23170 272956 23178 273124
rect 23212 272956 23220 273124
rect 22180 272940 22250 272950
rect 22140 272928 22180 272934
rect 22360 272940 22430 272950
rect 22250 272928 22360 272934
rect 22430 272928 23140 272934
rect 22140 272894 22152 272928
rect 23128 272894 23140 272928
rect 22140 272888 22180 272894
rect 21750 272520 21760 272530
rect 21330 272430 21400 272440
rect 20620 272414 21330 272420
rect 21510 272430 21580 272440
rect 21400 272414 21510 272420
rect 21580 272414 21620 272420
rect 20620 272380 20632 272414
rect 21608 272380 21620 272414
rect 20620 272374 21330 272380
rect 20540 272184 20548 272352
rect 20582 272184 20590 272352
rect 21400 272374 21510 272380
rect 21330 272350 21400 272360
rect 21580 272374 21620 272380
rect 21510 272350 21580 272360
rect 21650 272352 21700 272442
rect 20540 272094 20590 272184
rect 21650 272184 21658 272352
rect 21692 272184 21700 272352
rect 20660 272170 20730 272180
rect 20620 272156 20660 272162
rect 20840 272170 20910 272180
rect 20730 272156 20840 272162
rect 20910 272156 21620 272162
rect 20620 272122 20632 272156
rect 21608 272122 21620 272156
rect 20620 272116 20660 272122
rect 20540 271926 20548 272094
rect 20582 271926 20590 272094
rect 20730 272116 20840 272122
rect 20660 272090 20730 272100
rect 20910 272116 21620 272122
rect 20840 272090 20910 272100
rect 21650 272094 21700 272184
rect 20540 271836 20590 271926
rect 21650 271926 21658 272094
rect 21692 271926 21700 272094
rect 21330 271910 21400 271920
rect 20620 271898 21330 271904
rect 21510 271910 21580 271920
rect 21400 271898 21510 271904
rect 21580 271898 21620 271904
rect 20620 271864 20632 271898
rect 21608 271864 21620 271898
rect 20620 271858 21330 271864
rect 20540 271668 20548 271836
rect 20582 271668 20590 271836
rect 21400 271858 21510 271864
rect 21330 271830 21400 271840
rect 21580 271858 21620 271864
rect 21510 271830 21580 271840
rect 21650 271836 21700 271926
rect 20540 271578 20590 271668
rect 20660 271660 20730 271670
rect 20620 271640 20660 271646
rect 20840 271660 20910 271670
rect 20730 271640 20840 271646
rect 21650 271668 21658 271836
rect 21692 271668 21700 271836
rect 21754 271833 21760 272520
rect 21794 272520 21966 272530
rect 21794 271833 21800 272520
rect 21754 271821 21800 271833
rect 21960 271702 21966 272520
rect 22000 272520 22010 272790
rect 22060 272698 22068 272866
rect 22102 272698 22110 272866
rect 22250 272888 22360 272894
rect 22180 272860 22250 272870
rect 22430 272888 23140 272894
rect 22360 272860 22430 272870
rect 23170 272866 23220 272956
rect 22060 272608 22110 272698
rect 22850 272690 22920 272700
rect 22140 272670 22850 272676
rect 23030 272690 23100 272700
rect 22920 272670 23030 272676
rect 23170 272698 23178 272866
rect 23212 272698 23220 272866
rect 23100 272670 23140 272676
rect 22140 272636 22152 272670
rect 23128 272636 23140 272670
rect 22140 272630 22850 272636
rect 22920 272630 23030 272636
rect 22850 272610 22920 272620
rect 23100 272630 23140 272636
rect 23030 272610 23100 272620
rect 22000 271702 22006 272520
rect 21960 271690 22006 271702
rect 22060 272440 22068 272608
rect 22102 272440 22110 272608
rect 23170 272608 23220 272698
rect 23170 272440 23178 272608
rect 23212 272440 23220 272608
rect 22060 272350 22110 272440
rect 22180 272430 22250 272440
rect 22140 272412 22180 272418
rect 22360 272430 22430 272440
rect 22250 272412 22360 272418
rect 22430 272412 23140 272418
rect 22140 272378 22152 272412
rect 23128 272378 23140 272412
rect 22140 272372 22180 272378
rect 22250 272372 22360 272378
rect 22180 272350 22250 272360
rect 22430 272372 23140 272378
rect 22360 272350 22430 272360
rect 23170 272350 23220 272440
rect 22060 272182 22068 272350
rect 22102 272182 22110 272350
rect 22060 272092 22110 272182
rect 23170 272182 23178 272350
rect 23212 272182 23220 272350
rect 22850 272170 22920 272180
rect 22140 272154 22850 272160
rect 23030 272170 23100 272180
rect 22920 272154 23030 272160
rect 23100 272154 23140 272160
rect 22140 272120 22152 272154
rect 23128 272120 23140 272154
rect 22140 272114 22850 272120
rect 22060 271924 22068 272092
rect 22102 271924 22110 272092
rect 22920 272114 23030 272120
rect 22850 272090 22920 272100
rect 23100 272114 23140 272120
rect 23030 272090 23100 272100
rect 23170 272092 23220 272182
rect 22060 271834 22110 271924
rect 23170 271924 23178 272092
rect 23212 271924 23220 272092
rect 22180 271910 22250 271920
rect 22140 271896 22180 271902
rect 22360 271910 22430 271920
rect 22250 271896 22360 271902
rect 22430 271896 23140 271902
rect 22140 271862 22152 271896
rect 23128 271862 23140 271896
rect 22140 271856 22180 271862
rect 20910 271640 21620 271646
rect 20620 271606 20632 271640
rect 21608 271606 21620 271640
rect 20620 271600 20660 271606
rect 20730 271600 20840 271606
rect 20660 271580 20730 271590
rect 20910 271600 21620 271606
rect 20840 271580 20910 271590
rect 20540 271410 20548 271578
rect 20582 271410 20590 271578
rect 21650 271578 21700 271668
rect 21650 271410 21658 271578
rect 21692 271410 21700 271578
rect 20540 271320 20590 271410
rect 21330 271400 21400 271410
rect 20620 271382 21330 271388
rect 21510 271400 21580 271410
rect 21400 271382 21510 271388
rect 21580 271382 21620 271388
rect 20620 271348 20632 271382
rect 21608 271348 21620 271382
rect 20620 271342 21330 271348
rect 21400 271342 21510 271348
rect 21330 271320 21400 271330
rect 21580 271342 21620 271348
rect 21510 271320 21580 271330
rect 21650 271320 21700 271410
rect 20540 271152 20548 271320
rect 20582 271152 20590 271320
rect 20540 270630 20590 271152
rect 21650 271152 21658 271320
rect 21692 271152 21700 271320
rect 20660 271140 20730 271150
rect 20620 271124 20660 271130
rect 20840 271140 20910 271150
rect 20730 271124 20840 271130
rect 20910 271124 21620 271130
rect 20620 271090 20632 271124
rect 21608 271090 21620 271124
rect 20620 271084 20660 271090
rect 20730 271084 20840 271090
rect 20660 271060 20730 271070
rect 20910 271084 21620 271090
rect 20840 271060 20910 271070
rect 21650 270630 21700 271152
rect 22060 271666 22068 271834
rect 22102 271666 22110 271834
rect 22250 271856 22360 271862
rect 22180 271830 22250 271840
rect 22430 271856 23140 271862
rect 22360 271830 22430 271840
rect 23170 271834 23220 271924
rect 22060 271576 22110 271666
rect 23170 271666 23178 271834
rect 23212 271666 23220 271834
rect 23274 273604 23320 273616
rect 23274 271702 23280 273604
rect 23314 272790 23320 273604
rect 24090 273380 24140 273630
rect 24550 273560 24820 273570
rect 24550 273520 24570 273560
rect 24800 273520 24820 273560
rect 24400 273470 24480 273480
rect 24181 273442 24400 273448
rect 24550 273448 24820 273520
rect 24480 273442 25181 273448
rect 24181 273408 24193 273442
rect 25169 273408 25181 273442
rect 24181 273402 24400 273408
rect 24480 273402 25181 273408
rect 24550 273400 24820 273402
rect 24400 273380 24480 273390
rect 25220 273390 25270 273630
rect 26060 273670 26320 273730
rect 26060 273590 26080 273670
rect 26160 273590 26220 273670
rect 26300 273590 26320 273670
rect 26060 273566 26320 273590
rect 26060 273560 26322 273566
rect 26060 273520 26080 273560
rect 26310 273520 26322 273560
rect 26060 273514 26322 273520
rect 26060 273510 26320 273514
rect 28960 273490 30120 273550
rect 25860 273470 25940 273480
rect 25681 273442 25860 273448
rect 26720 273460 26840 273480
rect 25940 273442 26681 273448
rect 25681 273408 25693 273442
rect 26669 273408 26681 273442
rect 25681 273402 25860 273408
rect 25590 273390 25640 273400
rect 25220 273380 25300 273390
rect 24090 273212 24100 273380
rect 24134 273212 24140 273380
rect 24090 273122 24140 273212
rect 24880 273210 24960 273220
rect 24181 273184 24880 273190
rect 25220 273212 25228 273380
rect 25262 273300 25300 273310
rect 25560 273380 25640 273390
rect 25940 273402 26681 273408
rect 25860 273380 25940 273390
rect 26720 273380 26730 273460
rect 25560 273300 25600 273310
rect 25262 273212 25270 273300
rect 24960 273184 25181 273190
rect 24181 273150 24193 273184
rect 25169 273150 25181 273184
rect 24181 273144 24880 273150
rect 24090 272954 24100 273122
rect 24134 272954 24140 273122
rect 24960 273144 25181 273150
rect 24880 273120 24960 273130
rect 25220 273122 25270 273212
rect 24090 272864 24140 272954
rect 24400 272950 24480 272960
rect 24181 272926 24400 272932
rect 25220 272954 25228 273122
rect 25262 272954 25270 273122
rect 24480 272926 25181 272932
rect 24181 272892 24193 272926
rect 25169 272892 25181 272926
rect 24181 272886 24400 272892
rect 23314 272780 23530 272790
rect 23314 272520 23530 272530
rect 24090 272696 24100 272864
rect 24134 272696 24140 272864
rect 24480 272886 25181 272892
rect 24400 272860 24480 272870
rect 25220 272864 25270 272954
rect 24090 272606 24140 272696
rect 24880 272690 24960 272700
rect 24181 272668 24880 272674
rect 25220 272696 25228 272864
rect 25262 272700 25270 272864
rect 25590 273212 25600 273300
rect 25634 273212 25640 273380
rect 25590 273190 25640 273212
rect 26720 273212 26728 273380
rect 26830 273360 26840 273460
rect 26762 273340 26840 273360
rect 28960 273365 29010 273490
rect 29310 273440 29370 273450
rect 29040 273427 29310 273433
rect 29370 273427 30040 273433
rect 29040 273393 29052 273427
rect 30028 273393 30040 273427
rect 29040 273387 29310 273393
rect 29370 273387 30040 273393
rect 29310 273370 29370 273380
rect 26762 273212 26770 273340
rect 28360 273300 28460 273320
rect 28360 273220 28370 273300
rect 28450 273220 28460 273300
rect 26720 273190 26770 273212
rect 25590 273184 26770 273190
rect 25590 273150 25693 273184
rect 26669 273150 26770 273184
rect 25590 273144 26770 273150
rect 25590 273140 25800 273144
rect 26560 273140 26770 273144
rect 25590 273122 25640 273140
rect 25590 272954 25600 273122
rect 25634 272954 25640 273122
rect 26720 273122 26770 273140
rect 25590 272864 25640 272954
rect 25860 272950 25940 272960
rect 25681 272926 25860 272932
rect 26720 272954 26728 273122
rect 26762 272954 26770 273122
rect 28170 273210 28260 273220
rect 28250 273130 28260 273210
rect 28360 273190 28460 273220
rect 28360 273172 28370 273190
rect 28170 273120 28260 273130
rect 28290 273166 28370 273172
rect 28960 273197 28968 273365
rect 29002 273197 29010 273365
rect 28460 273166 28540 273172
rect 28290 273132 28302 273166
rect 28528 273132 28540 273166
rect 28290 273126 28370 273132
rect 28210 273104 28260 273120
rect 25940 272926 26681 272932
rect 25681 272892 25693 272926
rect 26669 272892 26681 272926
rect 25681 272886 25860 272892
rect 25590 272700 25600 272864
rect 25262 272696 25300 272700
rect 25220 272690 25300 272696
rect 24960 272668 25181 272674
rect 24181 272634 24193 272668
rect 25169 272634 25181 272668
rect 24181 272628 24880 272634
rect 23314 271702 23320 272520
rect 23274 271690 23320 271702
rect 24090 272438 24100 272606
rect 24134 272438 24140 272606
rect 24960 272628 25181 272634
rect 24880 272600 24960 272610
rect 25220 272620 25230 272690
rect 25220 272610 25300 272620
rect 25560 272696 25600 272700
rect 25634 272696 25640 272864
rect 25940 272886 26681 272892
rect 25860 272860 25940 272870
rect 26720 272864 26770 272954
rect 27470 273010 27590 273020
rect 27408 272930 27470 272936
rect 28210 272936 28218 273104
rect 28252 272936 28260 273104
rect 28460 273126 28540 273132
rect 28370 273090 28460 273100
rect 28570 273104 28620 273120
rect 27590 272930 27662 272936
rect 27408 272890 27420 272930
rect 27650 272890 27662 272930
rect 27408 272884 27662 272890
rect 28210 272920 28260 272936
rect 28570 272936 28578 273104
rect 28612 273060 28620 273104
rect 28960 273107 29010 273197
rect 30070 273365 30120 273490
rect 30070 273197 30078 273365
rect 30112 273197 30120 273365
rect 29720 273180 29780 273190
rect 29040 273169 29720 273175
rect 29780 273169 30040 273175
rect 29040 273135 29052 273169
rect 30028 273135 30040 273169
rect 29040 273129 29720 273135
rect 29780 273129 30040 273135
rect 29720 273110 29780 273120
rect 28960 273060 28968 273107
rect 28612 273050 28640 273060
rect 28612 272980 28640 272990
rect 28940 273050 28968 273060
rect 28940 272980 28968 272990
rect 28612 272936 28620 272980
rect 28570 272920 28620 272936
rect 28210 272914 28290 272920
rect 28530 272914 28620 272920
rect 28210 272908 28620 272914
rect 27470 272880 27590 272884
rect 25560 272690 25640 272696
rect 25630 272680 25640 272690
rect 26720 272696 26728 272864
rect 26762 272696 26770 272864
rect 28210 272874 28302 272908
rect 28528 272874 28620 272908
rect 28210 272870 28620 272874
rect 28210 272846 28260 272870
rect 28290 272868 28540 272870
rect 26720 272680 26770 272696
rect 27210 272816 27450 272820
rect 27780 272816 27870 272820
rect 27210 272810 27870 272816
rect 27210 272776 27302 272810
rect 27778 272776 27870 272810
rect 27210 272770 27870 272776
rect 27210 272748 27260 272770
rect 27210 272680 27218 272748
rect 27252 272680 27260 272748
rect 27820 272748 27870 272770
rect 27820 272680 27828 272748
rect 27862 272680 27870 272748
rect 28210 272680 28218 272846
rect 25630 272674 25800 272680
rect 26550 272674 26800 272680
rect 25630 272670 26800 272674
rect 25630 272668 26730 272670
rect 25630 272634 25693 272668
rect 26669 272634 26730 272668
rect 25630 272630 26730 272634
rect 25630 272620 25640 272630
rect 25681 272628 26681 272630
rect 25560 272610 25640 272620
rect 25220 272606 25270 272610
rect 24090 272348 24140 272438
rect 24400 272430 24480 272440
rect 24181 272410 24400 272416
rect 25220 272438 25228 272606
rect 25262 272438 25270 272606
rect 24480 272410 25181 272416
rect 24181 272376 24193 272410
rect 25169 272376 25181 272410
rect 24181 272370 24400 272376
rect 24090 272180 24100 272348
rect 24134 272180 24140 272348
rect 24480 272370 25181 272376
rect 24400 272340 24480 272350
rect 25220 272348 25270 272438
rect 25220 272180 25228 272348
rect 25262 272180 25270 272348
rect 24090 272090 24140 272180
rect 24880 272170 24960 272180
rect 24181 272152 24880 272158
rect 24960 272152 25181 272158
rect 24181 272118 24193 272152
rect 25169 272118 25181 272152
rect 24181 272112 24880 272118
rect 24090 271922 24100 272090
rect 24134 271922 24140 272090
rect 24960 272112 25181 272118
rect 24880 272080 24960 272090
rect 25220 272090 25270 272180
rect 22850 271650 22920 271660
rect 22140 271638 22850 271644
rect 23030 271650 23100 271660
rect 22920 271638 23030 271644
rect 23100 271638 23140 271644
rect 22140 271604 22152 271638
rect 23128 271604 23140 271638
rect 22140 271598 22850 271604
rect 22060 271408 22068 271576
rect 22102 271408 22110 271576
rect 22920 271598 23030 271604
rect 22850 271570 22920 271580
rect 23100 271598 23140 271604
rect 23030 271570 23100 271580
rect 23170 271576 23220 271666
rect 24090 271670 24140 271922
rect 24400 271920 24480 271930
rect 24181 271894 24400 271900
rect 25220 271922 25228 272090
rect 25262 272000 25270 272090
rect 25590 272606 25640 272610
rect 25590 272438 25600 272606
rect 25634 272438 25640 272606
rect 26720 272606 26730 272630
rect 25590 272348 25640 272438
rect 25860 272430 25940 272440
rect 25681 272410 25860 272416
rect 26720 272438 26728 272606
rect 26762 272590 26800 272600
rect 27170 272670 27260 272680
rect 27240 272600 27260 272670
rect 27640 272670 27710 272680
rect 27290 272652 27640 272658
rect 27710 272652 27790 272658
rect 27290 272618 27302 272652
rect 27778 272618 27790 272652
rect 27290 272612 27640 272618
rect 27170 272590 27260 272600
rect 27710 272612 27790 272618
rect 27640 272590 27710 272600
rect 27820 272590 27870 272680
rect 28170 272678 28218 272680
rect 28252 272678 28260 272846
rect 28570 272846 28620 272870
rect 28170 272670 28260 272678
rect 28240 272600 28260 272670
rect 28370 272680 28460 272690
rect 28290 272650 28370 272656
rect 28570 272678 28578 272846
rect 28612 272678 28620 272846
rect 28960 272939 28968 272980
rect 29002 272939 29010 273107
rect 28960 272849 29010 272939
rect 30070 273107 30120 273197
rect 30070 272939 30078 273107
rect 30112 272939 30120 273107
rect 29310 272920 29370 272930
rect 29040 272911 29310 272917
rect 29370 272911 30040 272917
rect 29040 272877 29052 272911
rect 30028 272877 30040 272911
rect 29040 272871 29310 272877
rect 29370 272871 30040 272877
rect 29310 272850 29370 272860
rect 28460 272650 28540 272656
rect 28290 272616 28302 272650
rect 28528 272616 28540 272650
rect 28290 272610 28370 272616
rect 28170 272590 28260 272600
rect 26762 272438 26770 272590
rect 27210 272522 27218 272590
rect 27252 272522 27260 272590
rect 27210 272500 27260 272522
rect 27820 272522 27828 272590
rect 27862 272522 27870 272590
rect 27820 272500 27870 272522
rect 27210 272494 27870 272500
rect 27210 272460 27302 272494
rect 27778 272460 27870 272494
rect 27210 272454 27870 272460
rect 27210 272450 27450 272454
rect 27780 272450 27870 272454
rect 28210 272588 28260 272590
rect 25940 272410 26681 272416
rect 25681 272376 25693 272410
rect 26669 272376 26681 272410
rect 25681 272370 25860 272376
rect 25590 272180 25600 272348
rect 25634 272180 25640 272348
rect 25940 272370 26681 272376
rect 25860 272340 25940 272350
rect 26720 272348 26770 272438
rect 28210 272420 28218 272588
rect 28252 272420 28260 272588
rect 28460 272610 28540 272616
rect 28370 272580 28460 272590
rect 28570 272588 28620 272678
rect 28210 272400 28260 272420
rect 28570 272420 28578 272588
rect 28612 272420 28620 272588
rect 28670 272740 28910 272760
rect 28670 272500 28680 272740
rect 28720 272670 28860 272740
rect 28720 272580 28750 272670
rect 28840 272580 28860 272670
rect 28720 272500 28860 272580
rect 28900 272500 28910 272740
rect 28670 272480 28910 272500
rect 28960 272681 28968 272849
rect 29002 272681 29010 272849
rect 28960 272591 29010 272681
rect 30070 272849 30120 272939
rect 30070 272681 30078 272849
rect 30112 272681 30120 272849
rect 30460 273180 30900 275540
rect 30460 273120 30490 273180
rect 30550 273120 30610 273180
rect 30670 273120 30730 273180
rect 30790 273120 30900 273180
rect 29720 272670 29780 272680
rect 29040 272653 29720 272659
rect 29780 272653 30040 272659
rect 29040 272619 29052 272653
rect 30028 272619 30040 272653
rect 29040 272613 29720 272619
rect 29780 272613 30040 272619
rect 29720 272600 29780 272610
rect 28570 272400 28620 272420
rect 27480 272390 27600 272400
rect 25590 272160 25640 272180
rect 26720 272180 26728 272348
rect 26762 272180 26770 272348
rect 27408 272380 27480 272386
rect 28210 272398 28300 272400
rect 28530 272398 28620 272400
rect 28210 272392 28620 272398
rect 27600 272380 27662 272386
rect 27408 272340 27420 272380
rect 27650 272340 27662 272380
rect 27408 272334 27480 272340
rect 27600 272334 27662 272340
rect 28210 272358 28302 272392
rect 28528 272358 28620 272392
rect 28210 272352 28620 272358
rect 28210 272350 28300 272352
rect 28530 272350 28620 272352
rect 27480 272260 27600 272270
rect 28210 272330 28260 272350
rect 28210 272180 28218 272330
rect 26720 272160 26770 272180
rect 25590 272158 25800 272160
rect 26560 272158 26770 272160
rect 25590 272152 26770 272158
rect 25590 272118 25693 272152
rect 26669 272118 26770 272152
rect 25590 272112 26770 272118
rect 25590 272110 25800 272112
rect 26560 272110 26770 272112
rect 25590 272090 25640 272110
rect 25590 272000 25600 272090
rect 25262 271990 25300 272000
rect 25220 271920 25230 271922
rect 25220 271910 25300 271920
rect 25560 271990 25600 272000
rect 25634 271922 25640 272090
rect 26720 272090 26770 272110
rect 25630 271920 25640 271922
rect 25560 271910 25640 271920
rect 24480 271894 25181 271900
rect 24181 271860 24193 271894
rect 25169 271860 25181 271894
rect 24181 271854 24400 271860
rect 24480 271854 25181 271860
rect 24400 271830 24480 271840
rect 24550 271780 24820 271854
rect 24550 271740 24570 271780
rect 24800 271740 24820 271780
rect 24550 271730 24820 271740
rect 25220 271670 25270 271910
rect 25590 271900 25640 271910
rect 25860 271920 25940 271930
rect 25681 271894 25860 271900
rect 26720 271922 26728 272090
rect 26762 271930 26770 272090
rect 28170 272170 28218 272180
rect 28252 272162 28260 272330
rect 28570 272330 28620 272350
rect 28250 272090 28260 272162
rect 28360 272160 28470 272170
rect 28360 272140 28370 272160
rect 28290 272134 28370 272140
rect 28460 272140 28470 272160
rect 28570 272162 28578 272330
rect 28612 272290 28620 272330
rect 28960 272423 28968 272591
rect 29002 272423 29010 272591
rect 28960 272333 29010 272423
rect 30070 272591 30120 272681
rect 30070 272423 30078 272591
rect 30112 272423 30120 272591
rect 30170 272740 30290 272760
rect 30170 272500 30180 272740
rect 30220 272670 30290 272740
rect 30280 272580 30290 272670
rect 30220 272500 30290 272580
rect 30170 272480 30290 272500
rect 29310 272410 29370 272420
rect 29040 272395 29310 272401
rect 29370 272395 30040 272401
rect 29040 272361 29052 272395
rect 30028 272361 30040 272395
rect 29040 272355 29310 272361
rect 29370 272355 30040 272361
rect 29310 272340 29370 272350
rect 28960 272290 28968 272333
rect 28612 272280 28640 272290
rect 28612 272210 28640 272220
rect 28940 272280 28968 272290
rect 28940 272210 28968 272220
rect 28612 272162 28620 272210
rect 28570 272140 28620 272162
rect 28960 272165 28968 272210
rect 29002 272165 29010 272333
rect 28460 272134 28540 272140
rect 28290 272100 28302 272134
rect 28528 272100 28540 272134
rect 28290 272094 28370 272100
rect 28170 272080 28260 272090
rect 28360 272070 28370 272094
rect 28460 272094 28540 272100
rect 28460 272070 28470 272094
rect 28360 272050 28470 272070
rect 28360 271960 28370 272050
rect 28460 271960 28470 272050
rect 28360 271940 28470 271960
rect 28960 272075 29010 272165
rect 30070 272333 30120 272423
rect 30070 272165 30078 272333
rect 30112 272165 30120 272333
rect 29720 272150 29780 272160
rect 29040 272137 29720 272143
rect 29780 272137 30040 272143
rect 29040 272103 29052 272137
rect 30028 272103 30040 272137
rect 29040 272097 29720 272103
rect 29780 272097 30040 272103
rect 29720 272080 29780 272090
rect 26762 271922 26840 271930
rect 26720 271910 26840 271922
rect 25940 271894 26681 271900
rect 25681 271860 25693 271894
rect 26669 271860 26681 271894
rect 25681 271854 25860 271860
rect 25940 271854 26681 271860
rect 25860 271830 25940 271840
rect 26720 271810 26730 271910
rect 26830 271810 26840 271910
rect 26720 271790 26840 271810
rect 28960 271907 28968 272075
rect 29002 271907 29010 272075
rect 24090 271600 25270 271670
rect 26060 271786 26320 271790
rect 26060 271780 26322 271786
rect 26060 271740 26080 271780
rect 26310 271740 26322 271780
rect 26060 271734 26322 271740
rect 28960 271780 29010 271907
rect 30070 272075 30120 272165
rect 30070 271907 30078 272075
rect 30112 271907 30120 272075
rect 29310 271890 29370 271900
rect 29040 271879 29310 271885
rect 29370 271879 30040 271885
rect 29040 271845 29052 271879
rect 30028 271845 30040 271879
rect 29040 271839 29310 271845
rect 29370 271839 30040 271845
rect 29310 271820 29370 271830
rect 30070 271780 30120 271907
rect 26060 271710 26320 271734
rect 28960 271720 30120 271780
rect 30460 272150 30900 273120
rect 30460 272090 30490 272150
rect 30550 272090 30610 272150
rect 30670 272090 30730 272150
rect 30790 272090 30900 272150
rect 26060 271630 26080 271710
rect 26160 271630 26220 271710
rect 26300 271630 26320 271710
rect 22060 271318 22110 271408
rect 22180 271400 22250 271410
rect 22140 271380 22180 271386
rect 22360 271400 22430 271410
rect 22250 271380 22360 271386
rect 23170 271408 23178 271576
rect 23212 271408 23220 271576
rect 26060 271570 26320 271630
rect 22430 271380 23140 271386
rect 22140 271346 22152 271380
rect 23128 271346 23140 271380
rect 22140 271340 22180 271346
rect 22250 271340 22360 271346
rect 22180 271320 22250 271330
rect 22430 271340 23140 271346
rect 22360 271320 22430 271330
rect 22060 271150 22068 271318
rect 22102 271150 22110 271318
rect 23170 271318 23220 271408
rect 23170 271150 23178 271318
rect 23212 271150 23220 271318
rect 22060 271060 22110 271150
rect 22850 271140 22920 271150
rect 22140 271122 22850 271128
rect 23030 271140 23100 271150
rect 22920 271122 23030 271128
rect 23100 271122 23140 271128
rect 22140 271088 22152 271122
rect 23128 271088 23140 271122
rect 22140 271082 22850 271088
rect 22920 271082 23030 271088
rect 22850 271060 22920 271070
rect 23100 271082 23140 271088
rect 23030 271060 23100 271070
rect 23170 271060 23220 271150
rect 22060 270892 22068 271060
rect 22102 270892 22110 271060
rect 22060 270630 22110 270892
rect 23170 270892 23178 271060
rect 23212 270892 23220 271060
rect 22180 270880 22250 270890
rect 22140 270864 22180 270870
rect 22360 270880 22430 270890
rect 22250 270864 22360 270870
rect 22430 270864 23140 270870
rect 22140 270830 22152 270864
rect 23128 270830 23140 270864
rect 22140 270824 22180 270830
rect 22250 270824 22360 270830
rect 22180 270800 22250 270810
rect 22430 270824 23140 270830
rect 22360 270800 22430 270810
rect 23170 270630 23220 270892
rect 20510 270620 20620 270630
rect 20510 270500 20620 270510
rect 21620 270620 21730 270630
rect 21620 270500 21730 270510
rect 22030 270620 22140 270630
rect 22030 270500 22140 270510
rect 23140 270620 23250 270630
rect 23140 270500 23250 270510
rect 20540 270380 20590 270500
rect 21650 270380 21700 270500
rect 22060 270380 22110 270500
rect 23170 270380 23220 270500
rect 20510 270370 20620 270380
rect 20510 270250 20620 270260
rect 21620 270370 21730 270380
rect 21620 270250 21730 270260
rect 22030 270370 22140 270380
rect 22030 270250 22140 270260
rect 23140 270370 23250 270380
rect 23140 270250 23250 270260
rect 20540 270240 20590 270250
rect 21650 270240 21700 270250
rect 22060 270240 22110 270250
rect 23170 270240 23220 270250
rect 12840 270160 12910 270170
rect 12801 270146 12840 270152
rect 13080 270160 13150 270170
rect 12910 270146 13080 270152
rect 13150 270146 13801 270152
rect 12801 270112 12813 270146
rect 13789 270112 13801 270146
rect 12801 270106 12840 270112
rect 12710 270016 12720 270084
rect 12754 270016 12760 270084
rect 12910 270106 13080 270112
rect 12840 270080 12910 270090
rect 13150 270106 13801 270112
rect 13080 270080 13150 270090
rect 13840 270084 13890 270174
rect 12710 269926 12760 270016
rect 13840 270016 13848 270084
rect 13882 270016 13890 270084
rect 13450 270000 13520 270010
rect 12801 269988 13450 269994
rect 13690 270000 13760 270010
rect 13520 269988 13690 269994
rect 13760 269988 13801 269994
rect 12801 269954 12813 269988
rect 13789 269954 13801 269988
rect 12801 269948 13450 269954
rect 12710 269858 12720 269926
rect 12754 269858 12760 269926
rect 13520 269948 13690 269954
rect 13450 269920 13520 269930
rect 13760 269948 13801 269954
rect 13690 269920 13760 269930
rect 13840 269926 13890 270016
rect 12710 269768 12760 269858
rect 12840 269850 12910 269860
rect 12801 269830 12840 269836
rect 13080 269850 13150 269860
rect 12910 269830 13080 269836
rect 13840 269858 13848 269926
rect 13882 269858 13890 269926
rect 19200 270100 20000 270200
rect 19200 270000 19300 270100
rect 19400 270000 19500 270100
rect 19700 270000 19800 270100
rect 19900 270000 20000 270100
rect 19200 269900 20000 270000
rect 13150 269830 13801 269836
rect 12801 269796 12813 269830
rect 13789 269796 13801 269830
rect 12801 269790 12840 269796
rect 12910 269790 13080 269796
rect 12840 269770 12910 269780
rect 13150 269790 13801 269796
rect 13080 269770 13150 269780
rect 12710 269700 12720 269768
rect 12754 269700 12760 269768
rect 13840 269768 13890 269858
rect 13840 269700 13848 269768
rect 13882 269700 13890 269768
rect 12710 269610 12760 269700
rect 13450 269690 13520 269700
rect 12801 269672 13450 269678
rect 13690 269690 13760 269700
rect 13520 269672 13690 269678
rect 13760 269672 13801 269678
rect 12801 269638 12813 269672
rect 13789 269638 13801 269672
rect 12801 269632 13450 269638
rect 13520 269632 13690 269638
rect 13450 269610 13520 269620
rect 13760 269632 13801 269638
rect 13690 269610 13760 269620
rect 13840 269610 13890 269700
rect 30460 269640 30900 272090
rect 12710 269542 12720 269610
rect 12754 269542 12760 269610
rect 12710 269410 12760 269542
rect 13840 269542 13848 269610
rect 13882 269542 13890 269610
rect 12840 269530 12910 269540
rect 12801 269514 12840 269520
rect 13080 269530 13150 269540
rect 12910 269514 13080 269520
rect 13150 269514 13801 269520
rect 12801 269480 12813 269514
rect 13789 269480 13801 269514
rect 12801 269474 12840 269480
rect 12910 269474 13080 269480
rect 12840 269450 12910 269460
rect 13150 269474 13801 269480
rect 13080 269450 13150 269460
rect 13840 269410 13890 269542
rect 12710 269330 13890 269410
rect 31014 269440 31266 269452
rect 13140 268560 13430 269330
rect 31014 269200 31020 269440
rect 31260 269200 31266 269440
rect 31014 269188 31266 269200
rect 32734 269440 32986 269452
rect 32734 269200 32740 269440
rect 32980 269200 32986 269440
rect 32734 269188 32986 269200
rect 34454 269440 34706 269452
rect 34454 269200 34460 269440
rect 34700 269200 34706 269440
rect 34454 269188 34706 269200
rect 35934 269440 36186 269452
rect 35934 269200 35940 269440
rect 36180 269200 36186 269440
rect 35934 269188 36186 269200
rect 37654 269440 37906 269452
rect 37654 269200 37660 269440
rect 37900 269200 37906 269440
rect 37654 269188 37906 269200
rect 39254 269440 39506 269452
rect 39254 269200 39260 269440
rect 39500 269200 39506 269440
rect 39254 269188 39506 269200
rect 40974 269440 41226 269452
rect 40974 269200 40980 269440
rect 41220 269200 41226 269440
rect 40974 269188 41226 269200
rect 42574 269440 42826 269452
rect 42574 269200 42580 269440
rect 42820 269200 42826 269440
rect 42574 269188 42826 269200
rect 44294 269440 44546 269452
rect 44294 269200 44300 269440
rect 44540 269200 44546 269440
rect 44294 269188 44546 269200
rect 44600 269440 45200 275900
rect 537352 275058 537496 275064
rect 537352 274938 537364 275058
rect 537484 274938 537496 275058
rect 537352 274932 537496 274938
rect 543722 275058 543866 275064
rect 543722 274938 543734 275058
rect 543854 274938 543866 275058
rect 543722 274932 543866 274938
rect 537352 272058 537496 272064
rect 537352 271938 537364 272058
rect 537484 271938 537496 272058
rect 537352 271932 537496 271938
rect 543722 272058 543866 272064
rect 543722 271938 543734 272058
rect 543854 271938 543866 272058
rect 543722 271932 543866 271938
rect 44600 269200 44780 269440
rect 45020 269200 45200 269440
rect 44600 268600 45200 269200
rect 537352 269058 537496 269064
rect 537352 268938 537364 269058
rect 537484 268938 537496 269058
rect 537352 268932 537496 268938
rect 543722 269058 543866 269064
rect 543722 268938 543734 269058
rect 543854 268938 543866 269058
rect 543722 268932 543866 268938
rect 11860 268539 14480 268560
rect 11860 268142 11887 268539
rect 13001 268142 13347 268539
rect 14461 268142 14480 268539
rect 11860 268120 14480 268142
rect 44600 268300 44700 268600
rect 45000 268300 45200 268600
rect 44600 268100 45200 268300
rect 44600 267800 44700 268100
rect 45000 267800 45200 268100
rect 44600 267600 45200 267800
rect 14534 267300 14646 267312
rect 14534 267120 14540 267300
rect 14640 267120 14646 267300
rect 14534 267108 14646 267120
rect 44600 267300 44700 267600
rect 45000 267300 45200 267600
rect 44600 267100 45200 267300
rect 537604 267759 543604 267798
rect 537604 267753 540807 267759
rect 537604 267728 537777 267753
rect 538891 267728 539297 267753
rect 540411 267728 540807 267753
rect 541921 267738 542317 267759
rect 543431 267738 543604 267759
rect 541921 267728 542294 267738
rect 537604 267318 537744 267728
rect 538914 267318 539254 267728
rect 540424 267318 540774 267728
rect 541944 267328 542294 267728
rect 543464 267328 543604 267738
rect 541944 267318 543604 267328
rect 537604 267298 543604 267318
rect 14534 266880 14646 266892
rect 14534 266700 14540 266880
rect 14640 266700 14646 266880
rect 14534 266688 14646 266700
rect 44600 266800 44700 267100
rect 45000 266800 45200 267100
rect 44600 266600 45200 266800
rect 44600 266300 44700 266600
rect 45000 266300 45200 266600
rect 11870 266108 14480 266130
rect 11870 265711 11887 266108
rect 13001 265711 13347 266108
rect 14461 265711 14480 266108
rect 11870 265690 14480 265711
rect 44600 266100 45200 266300
rect 44600 265800 44700 266100
rect 45000 265800 45200 266100
rect 13060 265000 13280 265690
rect 13060 264930 13080 265000
rect 13150 264930 13280 265000
rect 13060 264890 13280 264930
rect 13060 264820 13190 264890
rect 13260 264820 13280 264890
rect 13060 264800 13280 264820
rect 44600 265600 45200 265800
rect 44600 265300 44700 265600
rect 45000 265300 45200 265600
rect 44600 265100 45200 265300
rect 44600 264800 44700 265100
rect 45000 264800 45200 265100
rect 44600 264600 45200 264800
rect 44600 264300 44700 264600
rect 45000 264300 45200 264600
rect 44600 264100 45200 264300
rect 44600 263800 44700 264100
rect 45000 263800 45200 264100
rect 44600 263600 45200 263800
rect 44600 263300 44700 263600
rect 45000 263300 45200 263600
rect 44600 263100 45200 263300
rect 44600 262800 44700 263100
rect 45000 262800 45200 263100
rect 44600 262600 45200 262800
rect 44600 262300 44700 262600
rect 45000 262300 45200 262600
rect 44600 262100 45200 262300
rect 44600 261800 44700 262100
rect 45000 261800 45200 262100
rect 44600 261600 45200 261800
rect 44600 261300 44700 261600
rect 45000 261300 45200 261600
rect 44600 261100 45200 261300
rect 44600 260800 44700 261100
rect 45000 260800 45200 261100
rect 44600 260600 45200 260800
rect 14940 252580 15820 252600
rect 14940 252490 14980 252580
rect 5900 252478 14980 252490
rect 5900 252444 8420 252478
rect 13560 252460 14980 252478
rect 15100 252460 15160 252580
rect 15280 252460 15340 252580
rect 15460 252460 15520 252580
rect 15640 252460 15700 252580
rect 15820 252460 16170 252490
rect 13560 252444 16170 252460
rect 5900 252440 16170 252444
rect 8408 252438 13572 252440
rect 9680 252380 9740 252390
rect 5990 252364 9680 252370
rect 9845 252380 9905 252390
rect 9740 252364 9845 252370
rect 10045 252380 10105 252390
rect 9905 252364 10045 252370
rect 10235 252380 10295 252390
rect 10105 252364 10235 252370
rect 10415 252380 10475 252390
rect 10295 252364 10415 252370
rect 10615 252380 10675 252390
rect 10475 252364 10615 252370
rect 10805 252380 10865 252390
rect 10675 252364 10805 252370
rect 10965 252380 11025 252390
rect 10865 252364 10965 252370
rect 11155 252380 11215 252390
rect 11025 252364 11155 252370
rect 11330 252380 11390 252390
rect 11215 252364 11330 252370
rect 11470 252380 11530 252390
rect 11390 252364 11470 252370
rect 11530 252364 15990 252370
rect 5800 252320 5960 252340
rect 5990 252330 6002 252364
rect 15978 252330 15990 252364
rect 5990 252324 9680 252330
rect 5800 252200 5820 252320
rect 5940 252315 5960 252320
rect 5952 252281 5960 252315
rect 9740 252324 9845 252330
rect 9680 252310 9740 252320
rect 9905 252324 10045 252330
rect 9845 252310 9905 252320
rect 10105 252324 10235 252330
rect 10045 252310 10105 252320
rect 10295 252324 10415 252330
rect 10235 252310 10295 252320
rect 10475 252324 10615 252330
rect 10415 252310 10475 252320
rect 10675 252324 10805 252330
rect 10615 252310 10675 252320
rect 10865 252324 10965 252330
rect 10805 252310 10865 252320
rect 11025 252324 11155 252330
rect 10965 252310 11025 252320
rect 11215 252324 11330 252330
rect 11155 252310 11215 252320
rect 11390 252324 11470 252330
rect 11330 252310 11390 252320
rect 11530 252324 15990 252330
rect 11470 252310 11530 252320
rect 5940 252270 5960 252281
rect 15970 252272 16060 252280
rect 5990 252270 16060 252272
rect 5940 252266 16060 252270
rect 5940 252232 6002 252266
rect 15978 252232 16060 252266
rect 5940 252229 16060 252232
rect 5940 252226 16068 252229
rect 5940 252220 6000 252226
rect 15970 252220 16068 252226
rect 5940 252200 5960 252220
rect 5800 252120 5960 252200
rect 16020 252217 16068 252220
rect 9680 252180 9740 252190
rect 5990 252168 9680 252174
rect 9845 252180 9905 252190
rect 9740 252168 9845 252174
rect 10045 252180 10105 252190
rect 9905 252168 10045 252174
rect 10235 252180 10295 252190
rect 10105 252168 10235 252174
rect 10415 252180 10475 252190
rect 10295 252168 10415 252174
rect 10615 252180 10675 252190
rect 10475 252168 10615 252174
rect 10805 252180 10865 252190
rect 10675 252168 10805 252174
rect 10965 252180 11025 252190
rect 10865 252168 10965 252174
rect 11155 252180 11215 252190
rect 11025 252168 11155 252174
rect 11330 252180 11390 252190
rect 11215 252168 11330 252174
rect 11470 252180 11530 252190
rect 11390 252168 11470 252174
rect 16020 252183 16028 252217
rect 16062 252183 16068 252217
rect 11530 252168 15990 252174
rect 5990 252134 6002 252168
rect 15978 252134 15990 252168
rect 5990 252128 9680 252134
rect 5800 252000 5820 252120
rect 5940 252119 5960 252120
rect 5952 252085 5960 252119
rect 9740 252128 9845 252134
rect 9680 252110 9740 252120
rect 9905 252128 10045 252134
rect 9845 252110 9905 252120
rect 10105 252128 10235 252134
rect 10045 252110 10105 252120
rect 10295 252128 10415 252134
rect 10235 252110 10295 252120
rect 10475 252128 10615 252134
rect 10415 252110 10475 252120
rect 10675 252128 10805 252134
rect 10615 252110 10675 252120
rect 10865 252128 10965 252134
rect 10805 252110 10865 252120
rect 11025 252128 11155 252134
rect 10965 252110 11025 252120
rect 11215 252128 11330 252134
rect 11155 252110 11215 252120
rect 11390 252128 11470 252134
rect 11330 252110 11390 252120
rect 11530 252128 15990 252134
rect 16020 252171 16068 252183
rect 11470 252110 11530 252120
rect 5940 252080 5960 252085
rect 16020 252080 16060 252171
rect 5940 252076 6000 252080
rect 15970 252076 16060 252080
rect 5940 252070 16060 252076
rect 5940 252036 6002 252070
rect 15978 252036 16060 252070
rect 5940 252033 16060 252036
rect 16120 252150 16170 252440
rect 5940 252030 16068 252033
rect 5940 252000 5960 252030
rect 15970 252021 16068 252030
rect 15970 252020 16028 252021
rect 5800 251923 5960 252000
rect 9680 251980 9740 251990
rect 5990 251972 9680 251978
rect 9845 251980 9905 251990
rect 9740 251972 9845 251978
rect 10045 251980 10105 251990
rect 9905 251972 10045 251978
rect 10235 251980 10295 251990
rect 10105 251972 10235 251978
rect 10415 251980 10475 251990
rect 10295 251972 10415 251978
rect 10615 251980 10675 251990
rect 10475 251972 10615 251978
rect 10805 251980 10865 251990
rect 10675 251972 10805 251978
rect 10965 251980 11025 251990
rect 10865 251972 10965 251978
rect 11155 251980 11215 251990
rect 11025 251972 11155 251978
rect 11330 251980 11390 251990
rect 11215 251972 11330 251978
rect 11470 251980 11530 251990
rect 11390 251972 11470 251978
rect 16020 251987 16028 252020
rect 16062 251987 16068 252021
rect 11530 251972 15990 251978
rect 5990 251938 6002 251972
rect 15978 251938 15990 251972
rect 5990 251932 9680 251938
rect 5800 251920 5918 251923
rect 5800 251800 5820 251920
rect 5952 251889 5960 251923
rect 9740 251932 9845 251938
rect 9680 251910 9740 251920
rect 9905 251932 10045 251938
rect 9845 251910 9905 251920
rect 10105 251932 10235 251938
rect 10045 251910 10105 251920
rect 10295 251932 10415 251938
rect 10235 251910 10295 251920
rect 10475 251932 10615 251938
rect 10415 251910 10475 251920
rect 10675 251932 10805 251938
rect 10615 251910 10675 251920
rect 10865 251932 10965 251938
rect 10805 251910 10865 251920
rect 11025 251932 11155 251938
rect 10965 251910 11025 251920
rect 11215 251932 11330 251938
rect 11155 251910 11215 251920
rect 11390 251932 11470 251938
rect 11330 251910 11390 251920
rect 11530 251932 15990 251938
rect 16020 251975 16068 251987
rect 11470 251910 11530 251920
rect 16020 251890 16060 251975
rect 5940 251880 5960 251889
rect 15970 251880 16060 251890
rect 5940 251874 16060 251880
rect 5940 251840 6002 251874
rect 15978 251840 16060 251874
rect 5940 251837 16060 251840
rect 5940 251834 16068 251837
rect 5940 251830 6000 251834
rect 15970 251830 16068 251834
rect 5940 251800 5960 251830
rect 16020 251825 16068 251830
rect 5800 251727 5960 251800
rect 9680 251790 9740 251800
rect 5990 251776 9680 251782
rect 9845 251790 9905 251800
rect 9740 251776 9845 251782
rect 10045 251790 10105 251800
rect 9905 251776 10045 251782
rect 10235 251790 10295 251800
rect 10105 251776 10235 251782
rect 10415 251790 10475 251800
rect 10295 251776 10415 251782
rect 10615 251790 10675 251800
rect 10475 251776 10615 251782
rect 10805 251790 10865 251800
rect 10675 251776 10805 251782
rect 10965 251790 11025 251800
rect 10865 251776 10965 251782
rect 11155 251790 11215 251800
rect 11025 251776 11155 251782
rect 11330 251790 11390 251800
rect 11215 251776 11330 251782
rect 11470 251790 11530 251800
rect 11390 251776 11470 251782
rect 16020 251791 16028 251825
rect 16062 251791 16068 251825
rect 11530 251776 15990 251782
rect 5990 251742 6002 251776
rect 15978 251742 15990 251776
rect 5990 251736 9680 251742
rect 5800 251720 5918 251727
rect 5800 251600 5820 251720
rect 5952 251693 5960 251727
rect 9740 251736 9845 251742
rect 9680 251720 9740 251730
rect 9905 251736 10045 251742
rect 9845 251720 9905 251730
rect 10105 251736 10235 251742
rect 10045 251720 10105 251730
rect 10295 251736 10415 251742
rect 10235 251720 10295 251730
rect 10475 251736 10615 251742
rect 10415 251720 10475 251730
rect 10675 251736 10805 251742
rect 10615 251720 10675 251730
rect 10865 251736 10965 251742
rect 10805 251720 10865 251730
rect 11025 251736 11155 251742
rect 10965 251720 11025 251730
rect 11215 251736 11330 251742
rect 11155 251720 11215 251730
rect 11390 251736 11470 251742
rect 11330 251720 11390 251730
rect 11530 251736 15990 251742
rect 16020 251779 16068 251791
rect 11470 251720 11530 251730
rect 5940 251690 5960 251693
rect 16020 251690 16060 251779
rect 5940 251684 6000 251690
rect 15970 251684 16060 251690
rect 5940 251678 16060 251684
rect 5940 251644 6002 251678
rect 15978 251644 16060 251678
rect 5940 251641 16060 251644
rect 5940 251640 16068 251641
rect 5940 251600 5960 251640
rect 5990 251638 16068 251640
rect 15970 251630 16068 251638
rect 16020 251629 16068 251630
rect 5800 251531 5960 251600
rect 9680 251590 9740 251600
rect 5990 251580 9680 251586
rect 9845 251590 9905 251600
rect 9740 251580 9845 251586
rect 10045 251590 10105 251600
rect 9905 251580 10045 251586
rect 10235 251590 10295 251600
rect 10105 251580 10235 251586
rect 10415 251590 10475 251600
rect 10295 251580 10415 251586
rect 10615 251590 10675 251600
rect 10475 251580 10615 251586
rect 10805 251590 10865 251600
rect 10675 251580 10805 251586
rect 10965 251590 11025 251600
rect 10865 251580 10965 251586
rect 11155 251590 11215 251600
rect 11025 251580 11155 251586
rect 11330 251590 11390 251600
rect 11215 251580 11330 251586
rect 11470 251590 11530 251600
rect 11390 251580 11470 251586
rect 16020 251595 16028 251629
rect 16062 251595 16068 251629
rect 11530 251580 15990 251586
rect 5990 251546 6002 251580
rect 15978 251546 15990 251580
rect 5990 251540 9680 251546
rect 5800 251520 5918 251531
rect 5800 251400 5820 251520
rect 5952 251497 5960 251531
rect 9740 251540 9845 251546
rect 9680 251520 9740 251530
rect 9905 251540 10045 251546
rect 9845 251520 9905 251530
rect 10105 251540 10235 251546
rect 10045 251520 10105 251530
rect 10295 251540 10415 251546
rect 10235 251520 10295 251530
rect 10475 251540 10615 251546
rect 10415 251520 10475 251530
rect 10675 251540 10805 251546
rect 10615 251520 10675 251530
rect 10865 251540 10965 251546
rect 10805 251520 10865 251530
rect 11025 251540 11155 251546
rect 10965 251520 11025 251530
rect 11215 251540 11330 251546
rect 11155 251520 11215 251530
rect 11390 251540 11470 251546
rect 11330 251520 11390 251530
rect 11530 251540 15990 251546
rect 16020 251583 16068 251595
rect 11470 251520 11530 251530
rect 5940 251490 5960 251497
rect 16020 251490 16060 251583
rect 5940 251488 6000 251490
rect 15970 251488 16060 251490
rect 5940 251482 16060 251488
rect 5940 251448 6002 251482
rect 15978 251448 16060 251482
rect 5940 251445 16060 251448
rect 16120 251564 16130 252150
rect 16164 251564 16170 252150
rect 5940 251442 16068 251445
rect 5940 251440 6000 251442
rect 15970 251440 16068 251442
rect 5940 251400 5960 251440
rect 16020 251433 16068 251440
rect 5800 251380 5960 251400
rect 9680 251400 9740 251410
rect 5990 251384 9680 251390
rect 9845 251390 9905 251400
rect 10045 251390 10105 251400
rect 10235 251390 10295 251400
rect 10415 251390 10475 251400
rect 10615 251390 10675 251400
rect 10805 251390 10865 251400
rect 10965 251390 11025 251400
rect 11155 251390 11215 251400
rect 11330 251390 11390 251400
rect 11470 251390 11530 251400
rect 16020 251399 16028 251433
rect 16062 251399 16068 251433
rect 9740 251384 9845 251390
rect 9905 251384 10045 251390
rect 10105 251384 10235 251390
rect 10295 251384 10415 251390
rect 10475 251384 10615 251390
rect 10675 251384 10805 251390
rect 10865 251384 10965 251390
rect 11025 251384 11155 251390
rect 11215 251384 11330 251390
rect 11390 251384 11470 251390
rect 11530 251384 15990 251390
rect 5990 251350 6002 251384
rect 15978 251350 15990 251384
rect 16020 251387 16068 251399
rect 16020 251380 16060 251387
rect 5990 251344 9680 251350
rect 9740 251344 9845 251350
rect 9680 251330 9740 251340
rect 9905 251344 10045 251350
rect 9845 251320 9905 251330
rect 10105 251344 10235 251350
rect 10045 251320 10105 251330
rect 10295 251344 10415 251350
rect 10235 251320 10295 251330
rect 10475 251344 10615 251350
rect 10415 251320 10475 251330
rect 10675 251344 10805 251350
rect 10615 251320 10675 251330
rect 10865 251344 10965 251350
rect 10805 251320 10865 251330
rect 11025 251344 11155 251350
rect 10965 251320 11025 251330
rect 11215 251344 11330 251350
rect 11155 251320 11215 251330
rect 11390 251344 11470 251350
rect 11330 251320 11390 251330
rect 11530 251344 15990 251350
rect 11470 251320 11530 251330
rect 16120 251280 16170 251564
rect 5900 251270 16170 251280
rect 5900 251236 8420 251270
rect 13560 251236 16170 251270
rect 5900 251230 16170 251236
rect 16020 242090 16400 242120
rect 5900 242078 16400 242090
rect 5900 242044 8420 242078
rect 13560 242044 16400 242078
rect 5900 242040 16400 242044
rect 8408 242038 13572 242040
rect 16020 242000 16400 242040
rect 9680 241980 9740 241990
rect 5990 241964 9680 241970
rect 9845 241980 9905 241990
rect 9740 241964 9845 241970
rect 10045 241980 10105 241990
rect 9905 241964 10045 241970
rect 10235 241980 10295 241990
rect 10105 241964 10235 241970
rect 10415 241980 10475 241990
rect 10295 241964 10415 241970
rect 10615 241980 10675 241990
rect 10475 241964 10615 241970
rect 10805 241980 10865 241990
rect 10675 241964 10805 241970
rect 10965 241980 11025 241990
rect 10865 241964 10965 241970
rect 11155 241980 11215 241990
rect 11025 241964 11155 241970
rect 11330 241980 11390 241990
rect 11215 241964 11330 241970
rect 11470 241980 11530 241990
rect 11390 241964 11470 241970
rect 11530 241964 15990 241970
rect 5990 241930 6002 241964
rect 15978 241930 15990 241964
rect 5910 241927 5950 241930
rect 5910 241915 5958 241927
rect 5990 241924 9680 241930
rect 5910 241881 5918 241915
rect 5952 241881 5958 241915
rect 9740 241924 9845 241930
rect 9680 241910 9740 241920
rect 9905 241924 10045 241930
rect 9845 241910 9905 241920
rect 10105 241924 10235 241930
rect 10045 241910 10105 241920
rect 10295 241924 10415 241930
rect 10235 241910 10295 241920
rect 10475 241924 10615 241930
rect 10415 241910 10475 241920
rect 10675 241924 10805 241930
rect 10615 241910 10675 241920
rect 10865 241924 10965 241930
rect 10805 241910 10865 241920
rect 11025 241924 11155 241930
rect 10965 241910 11025 241920
rect 11215 241924 11330 241930
rect 11155 241910 11215 241920
rect 11390 241924 11470 241930
rect 11330 241910 11390 241920
rect 11530 241924 15990 241930
rect 11470 241910 11530 241920
rect 5910 241870 5958 241881
rect 16020 241880 16100 242000
rect 15970 241872 16100 241880
rect 5990 241870 16100 241872
rect 5910 241866 16100 241870
rect 5910 241832 6002 241866
rect 15978 241832 16100 241866
rect 5910 241826 16100 241832
rect 5910 241820 6000 241826
rect 15970 241820 16100 241826
rect 5910 241731 5950 241820
rect 16020 241817 16100 241820
rect 9680 241780 9740 241790
rect 5990 241768 9680 241774
rect 9845 241780 9905 241790
rect 9740 241768 9845 241774
rect 10045 241780 10105 241790
rect 9905 241768 10045 241774
rect 10235 241780 10295 241790
rect 10105 241768 10235 241774
rect 10415 241780 10475 241790
rect 10295 241768 10415 241774
rect 10615 241780 10675 241790
rect 10475 241768 10615 241774
rect 10805 241780 10865 241790
rect 10675 241768 10805 241774
rect 10965 241780 11025 241790
rect 10865 241768 10965 241774
rect 11155 241780 11215 241790
rect 11025 241768 11155 241774
rect 11330 241780 11390 241790
rect 11215 241768 11330 241774
rect 11470 241780 11530 241790
rect 11390 241768 11470 241774
rect 16020 241783 16028 241817
rect 16062 241800 16100 241817
rect 16300 241800 16400 242000
rect 16062 241783 16400 241800
rect 11530 241768 15990 241774
rect 5990 241734 6002 241768
rect 15978 241734 15990 241768
rect 5910 241719 5958 241731
rect 5990 241728 9680 241734
rect 5910 241685 5918 241719
rect 5952 241685 5958 241719
rect 9740 241728 9845 241734
rect 9680 241710 9740 241720
rect 9905 241728 10045 241734
rect 9845 241710 9905 241720
rect 10105 241728 10235 241734
rect 10045 241710 10105 241720
rect 10295 241728 10415 241734
rect 10235 241710 10295 241720
rect 10475 241728 10615 241734
rect 10415 241710 10475 241720
rect 10675 241728 10805 241734
rect 10615 241710 10675 241720
rect 10865 241728 10965 241734
rect 10805 241710 10865 241720
rect 11025 241728 11155 241734
rect 10965 241710 11025 241720
rect 11215 241728 11330 241734
rect 11155 241710 11215 241720
rect 11390 241728 11470 241734
rect 11330 241710 11390 241720
rect 11530 241728 15990 241734
rect 16020 241750 16400 241783
rect 11470 241710 11530 241720
rect 5910 241680 5958 241685
rect 16020 241700 16130 241750
rect 16164 241700 16400 241750
rect 16020 241680 16100 241700
rect 5910 241676 6000 241680
rect 15970 241676 16100 241680
rect 5910 241670 16100 241676
rect 5910 241636 6002 241670
rect 15978 241636 16100 241670
rect 5910 241630 16100 241636
rect 5910 241535 5950 241630
rect 15970 241621 16100 241630
rect 15970 241620 16028 241621
rect 9680 241580 9740 241590
rect 5990 241572 9680 241578
rect 9845 241580 9905 241590
rect 9740 241572 9845 241578
rect 10045 241580 10105 241590
rect 9905 241572 10045 241578
rect 10235 241580 10295 241590
rect 10105 241572 10235 241578
rect 10415 241580 10475 241590
rect 10295 241572 10415 241578
rect 10615 241580 10675 241590
rect 10475 241572 10615 241578
rect 10805 241580 10865 241590
rect 10675 241572 10805 241578
rect 10965 241580 11025 241590
rect 10865 241572 10965 241578
rect 11155 241580 11215 241590
rect 11025 241572 11155 241578
rect 11330 241580 11390 241590
rect 11215 241572 11330 241578
rect 11470 241580 11530 241590
rect 11390 241572 11470 241578
rect 16020 241587 16028 241620
rect 16062 241587 16100 241621
rect 11530 241572 15990 241578
rect 5990 241538 6002 241572
rect 15978 241538 15990 241572
rect 5910 241523 5958 241535
rect 5990 241532 9680 241538
rect 5910 241489 5918 241523
rect 5952 241489 5958 241523
rect 9740 241532 9845 241538
rect 9680 241510 9740 241520
rect 9905 241532 10045 241538
rect 9845 241510 9905 241520
rect 10105 241532 10235 241538
rect 10045 241510 10105 241520
rect 10295 241532 10415 241538
rect 10235 241510 10295 241520
rect 10475 241532 10615 241538
rect 10415 241510 10475 241520
rect 10675 241532 10805 241538
rect 10615 241510 10675 241520
rect 10865 241532 10965 241538
rect 10805 241510 10865 241520
rect 11025 241532 11155 241538
rect 10965 241510 11025 241520
rect 11215 241532 11330 241538
rect 11155 241510 11215 241520
rect 11390 241532 11470 241538
rect 11330 241510 11390 241520
rect 11530 241532 15990 241538
rect 11470 241510 11530 241520
rect 16020 241500 16100 241587
rect 16300 241500 16400 241700
rect 16020 241490 16130 241500
rect 5910 241480 5958 241489
rect 15970 241480 16130 241490
rect 5910 241474 16130 241480
rect 5910 241440 6002 241474
rect 15978 241440 16130 241474
rect 5910 241434 16130 241440
rect 5910 241430 6000 241434
rect 15970 241430 16130 241434
rect 5910 241339 5950 241430
rect 16020 241425 16130 241430
rect 9680 241390 9740 241400
rect 5990 241376 9680 241382
rect 9845 241390 9905 241400
rect 9740 241376 9845 241382
rect 10045 241390 10105 241400
rect 9905 241376 10045 241382
rect 10235 241390 10295 241400
rect 10105 241376 10235 241382
rect 10415 241390 10475 241400
rect 10295 241376 10415 241382
rect 10615 241390 10675 241400
rect 10475 241376 10615 241382
rect 10805 241390 10865 241400
rect 10675 241376 10805 241382
rect 10965 241390 11025 241400
rect 10865 241376 10965 241382
rect 11155 241390 11215 241400
rect 11025 241376 11155 241382
rect 11330 241390 11390 241400
rect 11215 241376 11330 241382
rect 11470 241390 11530 241400
rect 11390 241376 11470 241382
rect 16020 241391 16028 241425
rect 16062 241400 16130 241425
rect 16164 241400 16400 241500
rect 16062 241391 16100 241400
rect 11530 241376 15990 241382
rect 5990 241342 6002 241376
rect 15978 241342 15990 241376
rect 5910 241327 5958 241339
rect 5990 241336 9680 241342
rect 5910 241293 5918 241327
rect 5952 241293 5958 241327
rect 9740 241336 9845 241342
rect 9680 241320 9740 241330
rect 9905 241336 10045 241342
rect 9845 241320 9905 241330
rect 10105 241336 10235 241342
rect 10045 241320 10105 241330
rect 10295 241336 10415 241342
rect 10235 241320 10295 241330
rect 10475 241336 10615 241342
rect 10415 241320 10475 241330
rect 10675 241336 10805 241342
rect 10615 241320 10675 241330
rect 10865 241336 10965 241342
rect 10805 241320 10865 241330
rect 11025 241336 11155 241342
rect 10965 241320 11025 241330
rect 11215 241336 11330 241342
rect 11155 241320 11215 241330
rect 11390 241336 11470 241342
rect 11330 241320 11390 241330
rect 11530 241336 15990 241342
rect 11470 241320 11530 241330
rect 5910 241290 5958 241293
rect 16020 241290 16100 241391
rect 5910 241284 6000 241290
rect 15970 241284 16100 241290
rect 5910 241278 16100 241284
rect 5910 241244 6002 241278
rect 15978 241244 16100 241278
rect 5910 241240 16100 241244
rect 5910 241143 5950 241240
rect 5990 241238 16100 241240
rect 15970 241230 16100 241238
rect 16020 241229 16100 241230
rect 9680 241190 9740 241200
rect 5990 241180 9680 241186
rect 9845 241190 9905 241200
rect 9740 241180 9845 241186
rect 10045 241190 10105 241200
rect 9905 241180 10045 241186
rect 10235 241190 10295 241200
rect 10105 241180 10235 241186
rect 10415 241190 10475 241200
rect 10295 241180 10415 241186
rect 10615 241190 10675 241200
rect 10475 241180 10615 241186
rect 10805 241190 10865 241200
rect 10675 241180 10805 241186
rect 10965 241190 11025 241200
rect 10865 241180 10965 241186
rect 11155 241190 11215 241200
rect 11025 241180 11155 241186
rect 11330 241190 11390 241200
rect 11215 241180 11330 241186
rect 11470 241190 11530 241200
rect 11390 241180 11470 241186
rect 16020 241195 16028 241229
rect 16062 241200 16100 241229
rect 16300 241200 16400 241400
rect 16062 241195 16130 241200
rect 11530 241180 15990 241186
rect 5990 241146 6002 241180
rect 15978 241146 15990 241180
rect 5910 241131 5958 241143
rect 5990 241140 9680 241146
rect 5910 241097 5918 241131
rect 5952 241097 5958 241131
rect 9740 241140 9845 241146
rect 9680 241120 9740 241130
rect 9905 241140 10045 241146
rect 9845 241120 9905 241130
rect 10105 241140 10235 241146
rect 10045 241120 10105 241130
rect 10295 241140 10415 241146
rect 10235 241120 10295 241130
rect 10475 241140 10615 241146
rect 10415 241120 10475 241130
rect 10675 241140 10805 241146
rect 10615 241120 10675 241130
rect 10865 241140 10965 241146
rect 10805 241120 10865 241130
rect 11025 241140 11155 241146
rect 10965 241120 11025 241130
rect 11215 241140 11330 241146
rect 11155 241120 11215 241130
rect 11390 241140 11470 241146
rect 11330 241120 11390 241130
rect 11530 241140 15990 241146
rect 16020 241164 16130 241195
rect 16164 241164 16400 241200
rect 11470 241120 11530 241130
rect 5910 241090 5958 241097
rect 16020 241100 16400 241164
rect 16020 241090 16100 241100
rect 5910 241088 6000 241090
rect 15970 241088 16100 241090
rect 5910 241082 16100 241088
rect 5910 241048 6002 241082
rect 15978 241048 16100 241082
rect 5910 241042 16100 241048
rect 5910 241040 6000 241042
rect 15970 241040 16100 241042
rect 16020 241033 16100 241040
rect 9680 241000 9740 241010
rect 5990 240984 9680 240990
rect 9845 240990 9905 241000
rect 10045 240990 10105 241000
rect 10235 240990 10295 241000
rect 10415 240990 10475 241000
rect 10615 240990 10675 241000
rect 10805 240990 10865 241000
rect 10965 240990 11025 241000
rect 11155 240990 11215 241000
rect 11330 240990 11390 241000
rect 11470 240990 11530 241000
rect 16020 240999 16028 241033
rect 16062 240999 16100 241033
rect 9740 240984 9845 240990
rect 9905 240984 10045 240990
rect 10105 240984 10235 240990
rect 10295 240984 10415 240990
rect 10475 240984 10615 240990
rect 10675 240984 10805 240990
rect 10865 240984 10965 240990
rect 11025 240984 11155 240990
rect 11215 240984 11330 240990
rect 11390 240984 11470 240990
rect 11530 240984 15990 240990
rect 5990 240950 6002 240984
rect 15978 240950 15990 240984
rect 5990 240944 9680 240950
rect 9740 240944 9845 240950
rect 9680 240930 9740 240940
rect 9905 240944 10045 240950
rect 9845 240920 9905 240930
rect 10105 240944 10235 240950
rect 10045 240920 10105 240930
rect 10295 240944 10415 240950
rect 10235 240920 10295 240930
rect 10475 240944 10615 240950
rect 10415 240920 10475 240930
rect 10675 240944 10805 240950
rect 10615 240920 10675 240930
rect 10865 240944 10965 240950
rect 10805 240920 10865 240930
rect 11025 240944 11155 240950
rect 10965 240920 11025 240930
rect 11215 240944 11330 240950
rect 11155 240920 11215 240930
rect 11390 240944 11470 240950
rect 11330 240920 11390 240930
rect 11530 240944 15990 240950
rect 11470 240920 11530 240930
rect 16020 240900 16100 240999
rect 16300 240900 16400 241100
rect 16020 240880 16400 240900
rect 5900 240870 16400 240880
rect 5900 240836 8420 240870
rect 13560 240836 16400 240870
rect 5900 240830 16400 240836
rect 16020 240800 16400 240830
<< via1 >>
rect 23400 702060 23520 702180
rect 23600 702060 23720 702180
rect 23800 702060 23920 702180
rect 24000 702060 24120 702180
rect 24200 702060 24320 702180
rect 65060 702080 65240 702260
rect 65400 702080 65580 702260
rect 65740 702080 65920 702260
rect 563840 702020 563940 702120
rect 563980 702020 564080 702120
rect 564120 702020 564220 702120
rect 564260 702020 564360 702120
rect 564400 702020 564500 702120
rect 564540 702020 564640 702120
rect 564680 702020 564780 702120
rect 564820 702020 564920 702120
rect 564960 702020 565060 702120
rect 563840 701880 563940 701980
rect 563980 701880 564080 701980
rect 564120 701880 564220 701980
rect 564260 701880 564360 701980
rect 564400 701880 564500 701980
rect 564540 701880 564640 701980
rect 564680 701880 564780 701980
rect 564820 701880 564920 701980
rect 564960 701880 565060 701980
rect 573280 702140 573380 702240
rect 573420 702140 573520 702240
rect 573560 702140 573660 702240
rect 573700 702140 573800 702240
rect 573840 702140 573940 702240
rect 573980 702140 574080 702240
rect 573280 701880 573380 701980
rect 573420 701880 573520 701980
rect 573560 701880 573660 701980
rect 573700 701880 573800 701980
rect 573840 701880 573940 701980
rect 573980 701880 574080 701980
rect 24460 692900 24580 693020
rect 24460 692720 24580 692840
rect 24460 692540 24580 692660
rect 64720 692860 64860 693000
rect 64720 692660 64860 692800
rect 66060 692860 66200 693000
rect 66060 692660 66200 692800
rect 75120 692860 75260 693000
rect 75120 692660 75260 692800
rect 24460 692360 24580 692480
rect 24460 692180 24580 692300
rect 12900 691700 13100 691900
rect 13200 691700 13400 691900
rect 13500 691700 13700 691900
rect 13800 691700 14000 691900
rect 566300 690900 566500 691100
rect 566700 690900 566900 691100
rect 567100 690900 567300 691100
rect 567500 690900 567700 691100
rect 567900 690900 568100 691100
rect 568300 690900 568500 691100
rect 568700 690900 568900 691100
rect 569100 690900 569300 691100
rect 569500 690900 569700 691100
rect 569900 690900 570100 691100
rect 570300 690900 570500 691100
rect 570700 690900 570900 691100
rect 571100 690900 571300 691100
rect 571500 690900 571700 691100
rect 566300 690500 566500 690700
rect 566700 690500 566900 690700
rect 567100 690500 567300 690700
rect 567500 690500 567700 690700
rect 567900 690500 568100 690700
rect 568300 690500 568500 690700
rect 568700 690500 568900 690700
rect 569100 690500 569300 690700
rect 569500 690500 569700 690700
rect 569900 690500 570100 690700
rect 570300 690500 570500 690700
rect 570700 690500 570900 690700
rect 571100 690500 571300 690700
rect 571500 690500 571700 690700
rect 47200 690200 47300 690300
rect 47200 689800 47300 690000
rect 47200 689500 47300 689600
rect 566300 690100 566500 690300
rect 566700 690100 566900 690300
rect 567100 690100 567300 690300
rect 567500 690100 567700 690300
rect 567900 690100 568100 690300
rect 568300 690100 568500 690300
rect 568700 690100 568900 690300
rect 569100 690100 569300 690300
rect 569500 690100 569700 690300
rect 569900 690100 570100 690300
rect 570300 690100 570500 690300
rect 570700 690100 570900 690300
rect 571100 690100 571300 690300
rect 571500 690100 571700 690300
rect 566300 689700 566500 689900
rect 566700 689700 566900 689900
rect 567100 689700 567300 689900
rect 567500 689700 567700 689900
rect 567900 689700 568100 689900
rect 568300 689700 568500 689900
rect 568700 689700 568900 689900
rect 569100 689700 569300 689900
rect 569500 689700 569700 689900
rect 569900 689700 570100 689900
rect 570300 689700 570500 689900
rect 570700 689700 570900 689900
rect 571100 689700 571300 689900
rect 571500 689700 571700 689900
rect 566300 689300 566500 689500
rect 566700 689300 566900 689500
rect 567100 689300 567300 689500
rect 567500 689300 567700 689500
rect 567900 689300 568100 689500
rect 568300 689300 568500 689500
rect 568700 689300 568900 689500
rect 569100 689300 569300 689500
rect 569500 689300 569700 689500
rect 569900 689300 570100 689500
rect 570300 689300 570500 689500
rect 570700 689300 570900 689500
rect 571100 689300 571300 689500
rect 571500 689300 571700 689500
rect 42000 688600 42100 688700
rect 42000 688300 42100 688500
rect 42000 688100 42100 688200
rect 582360 684520 582440 684600
rect 582540 684520 582620 684600
rect 582360 684360 582440 684440
rect 582540 684360 582620 684440
rect 582360 684200 582440 684280
rect 582540 684200 582620 684280
rect 582360 684020 582440 684100
rect 582540 684020 582620 684100
rect 582360 683860 582440 683940
rect 582540 683860 582620 683940
rect 561700 682000 561900 682200
rect 562100 682000 562300 682200
rect 562500 682000 562700 682200
rect 562900 682000 563100 682200
rect 563300 682000 563500 682200
rect 561700 681600 561900 681800
rect 562100 681600 562300 681800
rect 562500 681600 562700 681800
rect 562900 681600 563100 681800
rect 563300 681600 563500 681800
rect 561700 681200 561900 681400
rect 562100 681200 562300 681400
rect 562500 681200 562700 681400
rect 562900 681200 563100 681400
rect 563300 681200 563500 681400
rect 561700 680800 561900 681000
rect 562100 680800 562300 681000
rect 562500 680800 562700 681000
rect 562900 680800 563100 681000
rect 563300 680800 563500 681000
rect 561700 680400 561900 680600
rect 562100 680400 562300 680600
rect 562500 680400 562700 680600
rect 562900 680400 563100 680600
rect 563300 680400 563500 680600
rect 561700 680000 561900 680200
rect 562100 680000 562300 680200
rect 562500 680000 562700 680200
rect 562900 680000 563100 680200
rect 563300 680000 563500 680200
rect 561700 679600 561900 679800
rect 562100 679600 562300 679800
rect 562500 679600 562700 679800
rect 562900 679600 563100 679800
rect 563300 679600 563500 679800
rect 561700 679200 561900 679400
rect 562100 679200 562300 679400
rect 562500 679200 562700 679400
rect 562900 679200 563100 679400
rect 563300 679200 563500 679400
rect 561700 678800 561900 679000
rect 562100 678800 562300 679000
rect 562500 678800 562700 679000
rect 562900 678800 563100 679000
rect 563300 678800 563500 679000
rect 561700 678400 561900 678600
rect 562100 678400 562300 678600
rect 562500 678400 562700 678600
rect 562900 678400 563100 678600
rect 563300 678400 563500 678600
rect 571900 677100 572100 677300
rect 571900 676800 572100 677000
rect 571900 676500 572100 676700
rect 571900 676200 572100 676400
rect 32800 663000 33100 663300
rect 33300 663000 33600 663300
rect 33800 663000 34100 663300
rect 34300 663000 34600 663300
rect 34800 663000 35100 663300
rect 35300 663000 35600 663300
rect 35800 663000 36100 663300
rect 36300 663000 36600 663300
rect 36800 663000 37100 663300
rect 37300 663000 37600 663300
rect 37800 663000 38100 663300
rect 38300 663000 38600 663300
rect 38800 663000 39100 663300
rect 39300 663000 39600 663300
rect 39800 663000 40100 663300
rect 40300 663000 40600 663300
rect 559840 306020 559940 306120
rect 559980 306020 560080 306120
rect 560120 306020 560220 306120
rect 560260 306020 560360 306120
rect 560400 306020 560500 306120
rect 560540 306020 560640 306120
rect 560680 306020 560780 306120
rect 560820 306020 560920 306120
rect 560960 306020 561060 306120
rect 559840 305880 559940 305980
rect 559980 305880 560080 305980
rect 560120 305882 560220 305980
rect 560120 305880 560131 305882
rect 560131 305880 560220 305882
rect 560260 305882 560360 305980
rect 560260 305880 560293 305882
rect 560293 305880 560327 305882
rect 560327 305880 560360 305882
rect 560400 305882 560500 305980
rect 560400 305880 560489 305882
rect 560489 305880 560500 305882
rect 560540 305880 560640 305980
rect 560680 305882 560780 305980
rect 560680 305880 560685 305882
rect 560685 305880 560719 305882
rect 560719 305880 560780 305882
rect 560820 305882 560920 305980
rect 560820 305880 560881 305882
rect 560881 305880 560915 305882
rect 560915 305880 560920 305882
rect 560960 305880 561060 305980
rect 569280 306140 569380 306240
rect 569420 306140 569520 306240
rect 569560 306140 569660 306240
rect 569700 306140 569800 306240
rect 569840 306140 569940 306240
rect 569980 306140 570080 306240
rect 9680 304364 9740 304380
rect 9845 304364 9905 304380
rect 10045 304364 10105 304380
rect 10235 304364 10295 304380
rect 10415 304364 10475 304380
rect 10615 304364 10675 304380
rect 10805 304364 10865 304380
rect 10965 304364 11025 304380
rect 11155 304364 11215 304380
rect 11330 304364 11390 304380
rect 11470 304364 11530 304380
rect 9680 304330 9740 304364
rect 9845 304330 9905 304364
rect 10045 304330 10105 304364
rect 10235 304330 10295 304364
rect 10415 304330 10475 304364
rect 10615 304330 10675 304364
rect 10805 304330 10865 304364
rect 10965 304330 11025 304364
rect 11155 304330 11215 304364
rect 11330 304330 11390 304364
rect 11470 304330 11530 304364
rect 9680 304320 9740 304330
rect 9845 304320 9905 304330
rect 10045 304320 10105 304330
rect 10235 304320 10295 304330
rect 10415 304320 10475 304330
rect 10615 304320 10675 304330
rect 10805 304320 10865 304330
rect 10965 304320 11025 304330
rect 11155 304320 11215 304330
rect 11330 304320 11390 304330
rect 11470 304320 11530 304330
rect 9680 304168 9740 304180
rect 9845 304168 9905 304180
rect 10045 304168 10105 304180
rect 10235 304168 10295 304180
rect 10415 304168 10475 304180
rect 10615 304168 10675 304180
rect 10805 304168 10865 304180
rect 10965 304168 11025 304180
rect 11155 304168 11215 304180
rect 11330 304168 11390 304180
rect 11470 304168 11530 304180
rect 9680 304134 9740 304168
rect 9845 304134 9905 304168
rect 10045 304134 10105 304168
rect 10235 304134 10295 304168
rect 10415 304134 10475 304168
rect 10615 304134 10675 304168
rect 10805 304134 10865 304168
rect 10965 304134 11025 304168
rect 11155 304134 11215 304168
rect 11330 304134 11390 304168
rect 11470 304134 11530 304168
rect 9680 304120 9740 304134
rect 9845 304120 9905 304134
rect 10045 304120 10105 304134
rect 10235 304120 10295 304134
rect 10415 304120 10475 304134
rect 10615 304120 10675 304134
rect 10805 304120 10865 304134
rect 10965 304120 11025 304134
rect 11155 304120 11215 304134
rect 11330 304120 11390 304134
rect 11470 304120 11530 304134
rect 9680 303972 9740 303980
rect 9845 303972 9905 303980
rect 10045 303972 10105 303980
rect 10235 303972 10295 303980
rect 10415 303972 10475 303980
rect 10615 303972 10675 303980
rect 10805 303972 10865 303980
rect 10965 303972 11025 303980
rect 11155 303972 11215 303980
rect 11330 303972 11390 303980
rect 11470 303972 11530 303980
rect 9680 303938 9740 303972
rect 9845 303938 9905 303972
rect 10045 303938 10105 303972
rect 10235 303938 10295 303972
rect 10415 303938 10475 303972
rect 10615 303938 10675 303972
rect 10805 303938 10865 303972
rect 10965 303938 11025 303972
rect 11155 303938 11215 303972
rect 11330 303938 11390 303972
rect 11470 303938 11530 303972
rect 9680 303920 9740 303938
rect 9845 303920 9905 303938
rect 10045 303920 10105 303938
rect 10235 303920 10295 303938
rect 10415 303920 10475 303938
rect 10615 303920 10675 303938
rect 10805 303920 10865 303938
rect 10965 303920 11025 303938
rect 11155 303920 11215 303938
rect 11330 303920 11390 303938
rect 11470 303920 11530 303938
rect 9680 303776 9740 303790
rect 9845 303776 9905 303790
rect 10045 303776 10105 303790
rect 10235 303776 10295 303790
rect 10415 303776 10475 303790
rect 10615 303776 10675 303790
rect 10805 303776 10865 303790
rect 10965 303776 11025 303790
rect 11155 303776 11215 303790
rect 11330 303776 11390 303790
rect 11470 303776 11530 303790
rect 9680 303742 9740 303776
rect 9845 303742 9905 303776
rect 10045 303742 10105 303776
rect 10235 303742 10295 303776
rect 10415 303742 10475 303776
rect 10615 303742 10675 303776
rect 10805 303742 10865 303776
rect 10965 303742 11025 303776
rect 11155 303742 11215 303776
rect 11330 303742 11390 303776
rect 11470 303742 11530 303776
rect 9680 303730 9740 303742
rect 9845 303730 9905 303742
rect 10045 303730 10105 303742
rect 10235 303730 10295 303742
rect 10415 303730 10475 303742
rect 10615 303730 10675 303742
rect 10805 303730 10865 303742
rect 10965 303730 11025 303742
rect 11155 303730 11215 303742
rect 11330 303730 11390 303742
rect 11470 303730 11530 303742
rect 9680 303580 9740 303590
rect 9845 303580 9905 303590
rect 10045 303580 10105 303590
rect 10235 303580 10295 303590
rect 10415 303580 10475 303590
rect 10615 303580 10675 303590
rect 10805 303580 10865 303590
rect 10965 303580 11025 303590
rect 11155 303580 11215 303590
rect 11330 303580 11390 303590
rect 11470 303580 11530 303590
rect 9680 303546 9740 303580
rect 9845 303546 9905 303580
rect 10045 303546 10105 303580
rect 10235 303546 10295 303580
rect 10415 303546 10475 303580
rect 10615 303546 10675 303580
rect 10805 303546 10865 303580
rect 10965 303546 11025 303580
rect 11155 303546 11215 303580
rect 11330 303546 11390 303580
rect 11470 303546 11530 303580
rect 9680 303530 9740 303546
rect 9845 303530 9905 303546
rect 10045 303530 10105 303546
rect 10235 303530 10295 303546
rect 10415 303530 10475 303546
rect 10615 303530 10675 303546
rect 10805 303530 10865 303546
rect 10965 303530 11025 303546
rect 11155 303530 11215 303546
rect 11330 303530 11390 303546
rect 11470 303530 11530 303546
rect 9680 303384 9740 303400
rect 9845 303384 9905 303390
rect 10045 303384 10105 303390
rect 10235 303384 10295 303390
rect 10415 303384 10475 303390
rect 10615 303384 10675 303390
rect 10805 303384 10865 303390
rect 10965 303384 11025 303390
rect 11155 303384 11215 303390
rect 11330 303384 11390 303390
rect 11470 303384 11530 303390
rect 9680 303350 9740 303384
rect 9845 303350 9905 303384
rect 10045 303350 10105 303384
rect 10235 303350 10295 303384
rect 10415 303350 10475 303384
rect 10615 303350 10675 303384
rect 10805 303350 10865 303384
rect 10965 303350 11025 303384
rect 11155 303350 11215 303384
rect 11330 303350 11390 303384
rect 11470 303350 11530 303384
rect 9680 303340 9740 303350
rect 9845 303330 9905 303350
rect 10045 303330 10105 303350
rect 10235 303330 10295 303350
rect 10415 303330 10475 303350
rect 10615 303330 10675 303350
rect 10805 303330 10865 303350
rect 10965 303330 11025 303350
rect 11155 303330 11215 303350
rect 11330 303330 11390 303350
rect 11470 303330 11530 303350
rect 15000 303120 15140 303260
rect 15200 303120 15340 303260
rect 559940 302060 559950 302120
rect 559950 302060 559984 302120
rect 559984 302060 560000 302120
rect 559930 301895 559950 301955
rect 559950 301895 559984 301955
rect 559984 301895 559990 301955
rect 559930 301695 559950 301755
rect 559950 301695 559984 301755
rect 559984 301695 559990 301755
rect 559930 301505 559950 301565
rect 559950 301505 559984 301565
rect 559984 301505 559990 301565
rect 559930 301325 559950 301385
rect 559950 301325 559984 301385
rect 559984 301325 559990 301385
rect 559930 301125 559950 301185
rect 559950 301125 559984 301185
rect 559984 301125 559990 301185
rect 559930 300935 559950 300995
rect 559950 300935 559984 300995
rect 559984 300935 559990 300995
rect 559930 300775 559950 300835
rect 559950 300775 559984 300835
rect 559984 300775 559990 300835
rect 559930 300585 559950 300645
rect 559950 300585 559984 300645
rect 559984 300585 559990 300645
rect 559930 300410 559950 300470
rect 559950 300410 559984 300470
rect 559984 300410 559990 300470
rect 559930 300270 559950 300330
rect 559950 300270 559984 300330
rect 559984 300270 559990 300330
rect 560130 302060 560146 302120
rect 560146 302060 560180 302120
rect 560180 302060 560190 302120
rect 560130 301895 560146 301955
rect 560146 301895 560180 301955
rect 560180 301895 560190 301955
rect 560130 301695 560146 301755
rect 560146 301695 560180 301755
rect 560180 301695 560190 301755
rect 560130 301505 560146 301565
rect 560146 301505 560180 301565
rect 560180 301505 560190 301565
rect 560130 301325 560146 301385
rect 560146 301325 560180 301385
rect 560180 301325 560190 301385
rect 560130 301125 560146 301185
rect 560146 301125 560180 301185
rect 560180 301125 560190 301185
rect 560130 300935 560146 300995
rect 560146 300935 560180 300995
rect 560180 300935 560190 300995
rect 560130 300775 560146 300835
rect 560146 300775 560180 300835
rect 560180 300775 560190 300835
rect 560130 300585 560146 300645
rect 560146 300585 560180 300645
rect 560180 300585 560190 300645
rect 560130 300410 560146 300470
rect 560146 300410 560180 300470
rect 560180 300410 560190 300470
rect 560130 300270 560146 300330
rect 560146 300270 560180 300330
rect 560180 300270 560190 300330
rect 560330 302060 560342 302120
rect 560342 302060 560376 302120
rect 560376 302060 560390 302120
rect 560330 301895 560342 301955
rect 560342 301895 560376 301955
rect 560376 301895 560390 301955
rect 560330 301695 560342 301755
rect 560342 301695 560376 301755
rect 560376 301695 560390 301755
rect 560330 301505 560342 301565
rect 560342 301505 560376 301565
rect 560376 301505 560390 301565
rect 560330 301325 560342 301385
rect 560342 301325 560376 301385
rect 560376 301325 560390 301385
rect 560330 301125 560342 301185
rect 560342 301125 560376 301185
rect 560376 301125 560390 301185
rect 560330 300935 560342 300995
rect 560342 300935 560376 300995
rect 560376 300935 560390 300995
rect 560330 300775 560342 300835
rect 560342 300775 560376 300835
rect 560376 300775 560390 300835
rect 560330 300585 560342 300645
rect 560342 300585 560376 300645
rect 560376 300585 560390 300645
rect 560330 300410 560342 300470
rect 560342 300410 560376 300470
rect 560376 300410 560390 300470
rect 560330 300270 560342 300330
rect 560342 300270 560376 300330
rect 560376 300270 560390 300330
rect 560520 302060 560538 302120
rect 560538 302060 560572 302120
rect 560572 302060 560580 302120
rect 560520 301895 560538 301955
rect 560538 301895 560572 301955
rect 560572 301895 560580 301955
rect 560520 301695 560538 301755
rect 560538 301695 560572 301755
rect 560572 301695 560580 301755
rect 560520 301505 560538 301565
rect 560538 301505 560572 301565
rect 560572 301505 560580 301565
rect 560520 301325 560538 301385
rect 560538 301325 560572 301385
rect 560572 301325 560580 301385
rect 560520 301125 560538 301185
rect 560538 301125 560572 301185
rect 560572 301125 560580 301185
rect 560520 300935 560538 300995
rect 560538 300935 560572 300995
rect 560572 300935 560580 300995
rect 560520 300775 560538 300835
rect 560538 300775 560572 300835
rect 560572 300775 560580 300835
rect 560520 300585 560538 300645
rect 560538 300585 560572 300645
rect 560572 300585 560580 300645
rect 560520 300410 560538 300470
rect 560538 300410 560572 300470
rect 560572 300410 560580 300470
rect 560520 300270 560538 300330
rect 560538 300270 560572 300330
rect 560572 300270 560580 300330
rect 560720 302060 560734 302120
rect 560734 302060 560768 302120
rect 560768 302060 560780 302120
rect 560720 301895 560734 301955
rect 560734 301895 560768 301955
rect 560768 301895 560780 301955
rect 560720 301695 560734 301755
rect 560734 301695 560768 301755
rect 560768 301695 560780 301755
rect 560720 301505 560734 301565
rect 560734 301505 560768 301565
rect 560768 301505 560780 301565
rect 560720 301325 560734 301385
rect 560734 301325 560768 301385
rect 560768 301325 560780 301385
rect 560720 301125 560734 301185
rect 560734 301125 560768 301185
rect 560768 301125 560780 301185
rect 560720 300935 560734 300995
rect 560734 300935 560768 300995
rect 560768 300935 560780 300995
rect 560720 300775 560734 300835
rect 560734 300775 560768 300835
rect 560768 300775 560780 300835
rect 560720 300585 560734 300645
rect 560734 300585 560768 300645
rect 560768 300585 560780 300645
rect 560720 300410 560734 300470
rect 560734 300410 560768 300470
rect 560768 300410 560780 300470
rect 560720 300270 560734 300330
rect 560734 300270 560768 300330
rect 560768 300270 560780 300330
rect 569280 305882 569380 305980
rect 569280 305880 569297 305882
rect 569297 305880 569331 305882
rect 569331 305880 569380 305882
rect 569420 305882 569520 305980
rect 569420 305880 569493 305882
rect 569493 305880 569520 305882
rect 569560 305880 569660 305980
rect 569700 305882 569800 305980
rect 569700 305880 569723 305882
rect 569723 305880 569800 305882
rect 569840 305882 569940 305980
rect 569840 305880 569885 305882
rect 569885 305880 569919 305882
rect 569919 305880 569940 305882
rect 569980 305880 570080 305980
rect 560920 302060 560930 302120
rect 560930 302060 560964 302120
rect 560964 302060 560980 302120
rect 560920 301895 560930 301955
rect 560930 301895 560964 301955
rect 560964 301895 560980 301955
rect 560920 301695 560930 301755
rect 560930 301695 560964 301755
rect 560964 301695 560980 301755
rect 560920 301505 560930 301565
rect 560930 301505 560964 301565
rect 560964 301505 560980 301565
rect 560920 301325 560930 301385
rect 560930 301325 560964 301385
rect 560964 301325 560980 301385
rect 560920 301125 560930 301185
rect 560930 301125 560964 301185
rect 560964 301125 560980 301185
rect 560920 300935 560930 300995
rect 560930 300935 560964 300995
rect 560964 300935 560980 300995
rect 560920 300775 560930 300835
rect 560930 300775 560964 300835
rect 560964 300775 560980 300835
rect 560920 300585 560930 300645
rect 560930 300585 560964 300645
rect 560964 300585 560980 300645
rect 560920 300410 560930 300470
rect 560930 300410 560964 300470
rect 560964 300410 560980 300470
rect 560920 300270 560930 300330
rect 560930 300270 560964 300330
rect 560964 300270 560980 300330
rect 569140 302060 569150 302120
rect 569150 302060 569184 302120
rect 569184 302060 569200 302120
rect 569130 301895 569150 301955
rect 569150 301895 569184 301955
rect 569184 301895 569190 301955
rect 569130 301695 569150 301755
rect 569150 301695 569184 301755
rect 569184 301695 569190 301755
rect 569130 301505 569150 301565
rect 569150 301505 569184 301565
rect 569184 301505 569190 301565
rect 569130 301325 569150 301385
rect 569150 301325 569184 301385
rect 569184 301325 569190 301385
rect 569130 301125 569150 301185
rect 569150 301125 569184 301185
rect 569184 301125 569190 301185
rect 569130 300935 569150 300995
rect 569150 300935 569184 300995
rect 569184 300935 569190 300995
rect 569130 300775 569150 300835
rect 569150 300775 569184 300835
rect 569184 300775 569190 300835
rect 569130 300585 569150 300645
rect 569150 300585 569184 300645
rect 569184 300585 569190 300645
rect 569130 300410 569150 300470
rect 569150 300410 569184 300470
rect 569184 300410 569190 300470
rect 569130 300270 569150 300330
rect 569150 300270 569184 300330
rect 569184 300270 569190 300330
rect 569330 302060 569346 302120
rect 569346 302060 569380 302120
rect 569380 302060 569390 302120
rect 569330 301895 569346 301955
rect 569346 301895 569380 301955
rect 569380 301895 569390 301955
rect 569330 301695 569346 301755
rect 569346 301695 569380 301755
rect 569380 301695 569390 301755
rect 569330 301505 569346 301565
rect 569346 301505 569380 301565
rect 569380 301505 569390 301565
rect 569330 301325 569346 301385
rect 569346 301325 569380 301385
rect 569380 301325 569390 301385
rect 569330 301125 569346 301185
rect 569346 301125 569380 301185
rect 569380 301125 569390 301185
rect 569330 300935 569346 300995
rect 569346 300935 569380 300995
rect 569380 300935 569390 300995
rect 569330 300775 569346 300835
rect 569346 300775 569380 300835
rect 569380 300775 569390 300835
rect 569330 300585 569346 300645
rect 569346 300585 569380 300645
rect 569380 300585 569390 300645
rect 569330 300410 569346 300470
rect 569346 300410 569380 300470
rect 569380 300410 569390 300470
rect 569330 300270 569346 300330
rect 569346 300270 569380 300330
rect 569380 300270 569390 300330
rect 569530 302060 569542 302120
rect 569542 302060 569576 302120
rect 569576 302060 569590 302120
rect 569530 301895 569542 301955
rect 569542 301895 569576 301955
rect 569576 301895 569590 301955
rect 569530 301695 569542 301755
rect 569542 301695 569576 301755
rect 569576 301695 569590 301755
rect 569530 301505 569542 301565
rect 569542 301505 569576 301565
rect 569576 301505 569590 301565
rect 569530 301325 569542 301385
rect 569542 301325 569576 301385
rect 569576 301325 569590 301385
rect 569530 301125 569542 301185
rect 569542 301125 569576 301185
rect 569576 301125 569590 301185
rect 569530 300935 569542 300995
rect 569542 300935 569576 300995
rect 569576 300935 569590 300995
rect 569530 300775 569542 300835
rect 569542 300775 569576 300835
rect 569576 300775 569590 300835
rect 569530 300585 569542 300645
rect 569542 300585 569576 300645
rect 569576 300585 569590 300645
rect 569530 300410 569542 300470
rect 569542 300410 569576 300470
rect 569576 300410 569590 300470
rect 569530 300270 569542 300330
rect 569542 300270 569576 300330
rect 569576 300270 569590 300330
rect 569720 302060 569738 302120
rect 569738 302060 569772 302120
rect 569772 302060 569780 302120
rect 569720 301895 569738 301955
rect 569738 301895 569772 301955
rect 569772 301895 569780 301955
rect 569720 301695 569738 301755
rect 569738 301695 569772 301755
rect 569772 301695 569780 301755
rect 569720 301505 569738 301565
rect 569738 301505 569772 301565
rect 569772 301505 569780 301565
rect 569720 301325 569738 301385
rect 569738 301325 569772 301385
rect 569772 301325 569780 301385
rect 569720 301125 569738 301185
rect 569738 301125 569772 301185
rect 569772 301125 569780 301185
rect 569720 300935 569738 300995
rect 569738 300935 569772 300995
rect 569772 300935 569780 300995
rect 569720 300775 569738 300835
rect 569738 300775 569772 300835
rect 569772 300775 569780 300835
rect 569720 300585 569738 300645
rect 569738 300585 569772 300645
rect 569772 300585 569780 300645
rect 569720 300410 569738 300470
rect 569738 300410 569772 300470
rect 569772 300410 569780 300470
rect 569720 300270 569738 300330
rect 569738 300270 569772 300330
rect 569772 300270 569780 300330
rect 569920 302060 569934 302120
rect 569934 302060 569968 302120
rect 569968 302060 569980 302120
rect 569920 301895 569934 301955
rect 569934 301895 569968 301955
rect 569968 301895 569980 301955
rect 569920 301695 569934 301755
rect 569934 301695 569968 301755
rect 569968 301695 569980 301755
rect 569920 301505 569934 301565
rect 569934 301505 569968 301565
rect 569968 301505 569980 301565
rect 569920 301325 569934 301385
rect 569934 301325 569968 301385
rect 569968 301325 569980 301385
rect 569920 301125 569934 301185
rect 569934 301125 569968 301185
rect 569968 301125 569980 301185
rect 569920 300935 569934 300995
rect 569934 300935 569968 300995
rect 569968 300935 569980 300995
rect 569920 300775 569934 300835
rect 569934 300775 569968 300835
rect 569968 300775 569980 300835
rect 569920 300585 569934 300645
rect 569934 300585 569968 300645
rect 569968 300585 569980 300645
rect 569920 300410 569934 300470
rect 569934 300410 569968 300470
rect 569968 300410 569980 300470
rect 569920 300270 569934 300330
rect 569934 300270 569968 300330
rect 569968 300270 569980 300330
rect 570120 302060 570130 302120
rect 570130 302060 570164 302120
rect 570164 302060 570180 302120
rect 570120 301895 570130 301955
rect 570130 301895 570164 301955
rect 570164 301895 570180 301955
rect 570120 301695 570130 301755
rect 570130 301695 570164 301755
rect 570164 301695 570180 301755
rect 570120 301505 570130 301565
rect 570130 301505 570164 301565
rect 570164 301505 570180 301565
rect 570120 301325 570130 301385
rect 570130 301325 570164 301385
rect 570164 301325 570180 301385
rect 570120 301125 570130 301185
rect 570130 301125 570164 301185
rect 570164 301125 570180 301185
rect 570120 300935 570130 300995
rect 570130 300935 570164 300995
rect 570164 300935 570180 300995
rect 570120 300775 570130 300835
rect 570130 300775 570164 300835
rect 570164 300775 570180 300835
rect 570120 300585 570130 300645
rect 570130 300585 570164 300645
rect 570164 300585 570180 300645
rect 570120 300410 570130 300470
rect 570130 300410 570164 300470
rect 570164 300410 570180 300470
rect 570120 300270 570130 300330
rect 570130 300270 570164 300330
rect 570164 300270 570180 300330
rect 537969 294892 538059 294962
rect 538139 294892 538229 294962
rect 540459 294892 540549 294962
rect 540629 294892 540719 294962
rect 542919 294892 542999 294972
rect 543089 294892 543169 294972
rect 562300 294900 562500 295100
rect 562700 294900 562900 295100
rect 563100 294900 563300 295100
rect 563500 294900 563700 295100
rect 563900 294900 564100 295100
rect 564300 294900 564500 295100
rect 564700 294900 564900 295100
rect 565100 294900 565300 295100
rect 565500 294900 565700 295100
rect 565900 294900 566100 295100
rect 566300 294900 566500 295100
rect 566700 294900 566900 295100
rect 567100 294900 567300 295100
rect 567500 294900 567700 295100
rect 537969 294784 538049 294852
rect 538139 294784 538219 294852
rect 540459 294784 540539 294852
rect 540629 294784 540709 294852
rect 542919 294784 542999 294842
rect 543089 294784 543169 294842
rect 537969 294772 538049 294784
rect 538139 294772 538219 294784
rect 540459 294772 540539 294784
rect 540629 294772 540709 294784
rect 542919 294762 542999 294784
rect 543089 294762 543169 294784
rect 537089 294626 537169 294682
rect 537239 294626 537319 294682
rect 537419 294654 537449 294722
rect 537449 294654 537523 294722
rect 537523 294654 537549 294722
rect 538659 294654 538685 294722
rect 538685 294654 538759 294722
rect 538759 294654 538789 294722
rect 537419 294652 537549 294654
rect 538659 294652 538789 294654
rect 539579 294626 539659 294682
rect 539729 294626 539809 294682
rect 539889 294654 539921 294722
rect 539921 294654 539995 294722
rect 539995 294654 540019 294722
rect 541129 294654 541157 294722
rect 541157 294654 541231 294722
rect 541231 294654 541259 294722
rect 539889 294652 540019 294654
rect 541129 294652 541259 294654
rect 542059 294626 542139 294682
rect 542209 294626 542289 294682
rect 542369 294654 542393 294722
rect 542393 294654 542467 294722
rect 542467 294654 542499 294722
rect 543599 294654 543629 294722
rect 543629 294654 543703 294722
rect 543703 294654 543729 294722
rect 542369 294652 542499 294654
rect 543599 294652 543729 294654
rect 536699 294592 536779 294612
rect 536869 294592 536949 294612
rect 537089 294602 537169 294626
rect 537239 294602 537319 294626
rect 539219 294592 539299 294612
rect 539389 294592 539469 294612
rect 539579 294602 539659 294626
rect 539729 294602 539809 294626
rect 541709 294592 541789 294612
rect 541879 294592 541959 294612
rect 542059 294602 542139 294626
rect 542209 294602 542289 294626
rect 544159 294592 544239 294612
rect 544329 294592 544409 294612
rect 536699 294532 536779 294592
rect 536869 294532 536949 294592
rect 539219 294532 539299 294592
rect 539389 294532 539469 294592
rect 541709 294532 541789 294592
rect 541879 294532 541959 294592
rect 544159 294532 544239 294592
rect 544329 294532 544409 294592
rect 562300 294500 562500 294700
rect 562700 294500 562900 294700
rect 563100 294500 563300 294700
rect 563500 294500 563700 294700
rect 563900 294500 564100 294700
rect 564300 294500 564500 294700
rect 564700 294500 564900 294700
rect 565100 294500 565300 294700
rect 565500 294500 565700 294700
rect 565900 294500 566100 294700
rect 566300 294500 566500 294700
rect 566700 294500 566900 294700
rect 567100 294500 567300 294700
rect 567500 294500 567700 294700
rect 537969 294244 538049 294312
rect 538139 294244 538219 294312
rect 540459 294244 540539 294312
rect 540629 294244 540709 294312
rect 542919 294244 542999 294302
rect 543089 294244 543169 294302
rect 537969 294232 538049 294244
rect 538139 294232 538219 294244
rect 540459 294232 540539 294244
rect 540629 294232 540709 294244
rect 542919 294222 542999 294244
rect 543089 294222 543169 294244
rect 15000 294060 15140 294200
rect 15200 294060 15340 294200
rect 9680 293964 9740 293980
rect 9845 293964 9905 293980
rect 10045 293964 10105 293980
rect 10235 293964 10295 293980
rect 10415 293964 10475 293980
rect 10615 293964 10675 293980
rect 10805 293964 10865 293980
rect 10965 293964 11025 293980
rect 11155 293964 11215 293980
rect 11330 293964 11390 293980
rect 11470 293964 11530 293980
rect 9680 293930 9740 293964
rect 9845 293930 9905 293964
rect 10045 293930 10105 293964
rect 10235 293930 10295 293964
rect 10415 293930 10475 293964
rect 10615 293930 10675 293964
rect 10805 293930 10865 293964
rect 10965 293930 11025 293964
rect 11155 293930 11215 293964
rect 11330 293930 11390 293964
rect 11470 293930 11530 293964
rect 5740 293915 5920 293920
rect 5740 293881 5918 293915
rect 5918 293881 5920 293915
rect 9680 293920 9740 293930
rect 9845 293920 9905 293930
rect 10045 293920 10105 293930
rect 10235 293920 10295 293930
rect 10415 293920 10475 293930
rect 10615 293920 10675 293930
rect 10805 293920 10865 293930
rect 10965 293920 11025 293930
rect 11155 293920 11215 293930
rect 11330 293920 11390 293930
rect 11470 293920 11530 293930
rect 5740 293740 5920 293881
rect 9680 293768 9740 293780
rect 9845 293768 9905 293780
rect 10045 293768 10105 293780
rect 10235 293768 10295 293780
rect 10415 293768 10475 293780
rect 10615 293768 10675 293780
rect 10805 293768 10865 293780
rect 10965 293768 11025 293780
rect 11155 293768 11215 293780
rect 11330 293768 11390 293780
rect 11470 293768 11530 293780
rect 9680 293734 9740 293768
rect 9845 293734 9905 293768
rect 10045 293734 10105 293768
rect 10235 293734 10295 293768
rect 10415 293734 10475 293768
rect 10615 293734 10675 293768
rect 10805 293734 10865 293768
rect 10965 293734 11025 293768
rect 11155 293734 11215 293768
rect 11330 293734 11390 293768
rect 11470 293734 11530 293768
rect 9680 293720 9740 293734
rect 9845 293720 9905 293734
rect 10045 293720 10105 293734
rect 10235 293720 10295 293734
rect 10415 293720 10475 293734
rect 10615 293720 10675 293734
rect 10805 293720 10865 293734
rect 10965 293720 11025 293734
rect 11155 293720 11215 293734
rect 11330 293720 11390 293734
rect 11470 293720 11530 293734
rect 537089 294086 537169 294142
rect 537239 294086 537319 294142
rect 537419 294114 537449 294182
rect 537449 294114 537523 294182
rect 537523 294114 537549 294182
rect 538659 294114 538685 294182
rect 538685 294114 538759 294182
rect 538759 294114 538789 294182
rect 537419 294112 537549 294114
rect 538659 294112 538789 294114
rect 539579 294086 539659 294142
rect 539729 294086 539809 294142
rect 539889 294114 539921 294182
rect 539921 294114 539995 294182
rect 539995 294114 540019 294182
rect 541129 294114 541157 294182
rect 541157 294114 541231 294182
rect 541231 294114 541259 294182
rect 539889 294112 540019 294114
rect 541129 294112 541259 294114
rect 542059 294086 542139 294142
rect 542209 294086 542289 294142
rect 542369 294114 542393 294182
rect 542393 294114 542467 294182
rect 542467 294114 542499 294182
rect 543599 294114 543629 294182
rect 543629 294114 543703 294182
rect 543703 294114 543729 294182
rect 542369 294112 542499 294114
rect 543599 294112 543729 294114
rect 536699 294052 536779 294072
rect 536869 294052 536949 294072
rect 537089 294062 537169 294086
rect 537239 294062 537319 294086
rect 539219 294052 539299 294072
rect 539389 294052 539469 294072
rect 539579 294062 539659 294086
rect 539729 294062 539809 294086
rect 541709 294052 541789 294072
rect 541879 294052 541959 294072
rect 542059 294062 542139 294086
rect 542209 294062 542289 294086
rect 544159 294052 544239 294062
rect 544329 294052 544409 294062
rect 536699 293992 536779 294052
rect 536869 293992 536949 294052
rect 539219 293992 539299 294052
rect 539389 293992 539469 294052
rect 541709 293992 541789 294052
rect 541879 293992 541959 294052
rect 544159 293982 544239 294052
rect 544329 293982 544409 294052
rect 562300 294100 562500 294300
rect 562700 294100 562900 294300
rect 563100 294100 563300 294300
rect 563500 294100 563700 294300
rect 563900 294100 564100 294300
rect 564300 294100 564500 294300
rect 564700 294100 564900 294300
rect 565100 294100 565300 294300
rect 565500 294100 565700 294300
rect 565900 294100 566100 294300
rect 566300 294100 566500 294300
rect 566700 294100 566900 294300
rect 567100 294100 567300 294300
rect 567500 294100 567700 294300
rect 537979 293842 538069 293912
rect 538119 293842 538209 293912
rect 540459 293842 540549 293912
rect 540619 293852 540709 293922
rect 542919 293852 542999 293922
rect 543089 293852 543169 293922
rect 5740 293523 5920 293580
rect 9680 293572 9740 293580
rect 9845 293572 9905 293580
rect 10045 293572 10105 293580
rect 10235 293572 10295 293580
rect 10415 293572 10475 293580
rect 10615 293572 10675 293580
rect 10805 293572 10865 293580
rect 10965 293572 11025 293580
rect 11155 293572 11215 293580
rect 11330 293572 11390 293580
rect 11470 293572 11530 293580
rect 9680 293538 9740 293572
rect 9845 293538 9905 293572
rect 10045 293538 10105 293572
rect 10235 293538 10295 293572
rect 10415 293538 10475 293572
rect 10615 293538 10675 293572
rect 10805 293538 10865 293572
rect 10965 293538 11025 293572
rect 11155 293538 11215 293572
rect 11330 293538 11390 293572
rect 11470 293538 11530 293572
rect 5740 293489 5918 293523
rect 5918 293489 5920 293523
rect 9680 293520 9740 293538
rect 9845 293520 9905 293538
rect 10045 293520 10105 293538
rect 10235 293520 10295 293538
rect 10415 293520 10475 293538
rect 10615 293520 10675 293538
rect 10805 293520 10865 293538
rect 10965 293520 11025 293538
rect 11155 293520 11215 293538
rect 11330 293520 11390 293538
rect 11470 293520 11530 293538
rect 5740 293400 5920 293489
rect 9680 293376 9740 293390
rect 9845 293376 9905 293390
rect 10045 293376 10105 293390
rect 10235 293376 10295 293390
rect 10415 293376 10475 293390
rect 10615 293376 10675 293390
rect 10805 293376 10865 293390
rect 10965 293376 11025 293390
rect 11155 293376 11215 293390
rect 11330 293376 11390 293390
rect 11470 293376 11530 293390
rect 9680 293342 9740 293376
rect 9845 293342 9905 293376
rect 10045 293342 10105 293376
rect 10235 293342 10295 293376
rect 10415 293342 10475 293376
rect 10615 293342 10675 293376
rect 10805 293342 10865 293376
rect 10965 293342 11025 293376
rect 11155 293342 11215 293376
rect 11330 293342 11390 293376
rect 11470 293342 11530 293376
rect 9680 293330 9740 293342
rect 9845 293330 9905 293342
rect 10045 293330 10105 293342
rect 10235 293330 10295 293342
rect 10415 293330 10475 293342
rect 10615 293330 10675 293342
rect 10805 293330 10865 293342
rect 10965 293330 11025 293342
rect 11155 293330 11215 293342
rect 11330 293330 11390 293342
rect 11470 293330 11530 293342
rect 5740 293131 5920 293240
rect 9680 293180 9740 293190
rect 9845 293180 9905 293190
rect 10045 293180 10105 293190
rect 10235 293180 10295 293190
rect 10415 293180 10475 293190
rect 10615 293180 10675 293190
rect 10805 293180 10865 293190
rect 10965 293180 11025 293190
rect 11155 293180 11215 293190
rect 11330 293180 11390 293190
rect 11470 293180 11530 293190
rect 9680 293146 9740 293180
rect 9845 293146 9905 293180
rect 10045 293146 10105 293180
rect 10235 293146 10295 293180
rect 10415 293146 10475 293180
rect 10615 293146 10675 293180
rect 10805 293146 10865 293180
rect 10965 293146 11025 293180
rect 11155 293146 11215 293180
rect 11330 293146 11390 293180
rect 11470 293146 11530 293180
rect 5740 293097 5918 293131
rect 5918 293097 5920 293131
rect 9680 293130 9740 293146
rect 9845 293130 9905 293146
rect 10045 293130 10105 293146
rect 10235 293130 10295 293146
rect 10415 293130 10475 293146
rect 10615 293130 10675 293146
rect 10805 293130 10865 293146
rect 10965 293130 11025 293146
rect 11155 293130 11215 293146
rect 11330 293130 11390 293146
rect 11470 293130 11530 293146
rect 5740 293060 5920 293097
rect 537969 293704 538049 293772
rect 538139 293704 538219 293772
rect 540459 293704 540539 293782
rect 540629 293704 540709 293782
rect 542919 293704 542999 293762
rect 543089 293704 543169 293762
rect 537969 293692 538049 293704
rect 538139 293692 538219 293704
rect 540459 293702 540539 293704
rect 540629 293702 540709 293704
rect 542919 293682 542999 293704
rect 543089 293682 543169 293704
rect 562300 293700 562500 293900
rect 562700 293700 562900 293900
rect 563100 293700 563300 293900
rect 563500 293700 563700 293900
rect 563900 293700 564100 293900
rect 564300 293700 564500 293900
rect 564700 293700 564900 293900
rect 565100 293700 565300 293900
rect 565500 293700 565700 293900
rect 565900 293700 566100 293900
rect 566300 293700 566500 293900
rect 566700 293700 566900 293900
rect 567100 293700 567300 293900
rect 567500 293700 567700 293900
rect 537089 293546 537169 293602
rect 537239 293546 537319 293602
rect 537419 293574 537449 293642
rect 537449 293574 537523 293642
rect 537523 293574 537549 293642
rect 538659 293574 538685 293642
rect 538685 293574 538759 293642
rect 538759 293574 538789 293642
rect 537419 293572 537549 293574
rect 538659 293572 538789 293574
rect 539579 293546 539659 293602
rect 539729 293546 539809 293602
rect 539889 293574 539921 293642
rect 539921 293574 539995 293642
rect 539995 293574 540019 293642
rect 541129 293574 541157 293642
rect 541157 293574 541231 293642
rect 541231 293574 541259 293642
rect 539889 293572 540019 293574
rect 541129 293572 541259 293574
rect 542069 293546 542149 293602
rect 542209 293546 542289 293602
rect 542369 293574 542393 293642
rect 542393 293574 542467 293642
rect 542467 293574 542499 293642
rect 543599 293574 543629 293642
rect 543629 293574 543703 293642
rect 543703 293574 543729 293642
rect 542369 293572 542499 293574
rect 543599 293572 543729 293574
rect 536699 293512 536779 293532
rect 536869 293512 536949 293532
rect 537089 293522 537169 293546
rect 537239 293522 537319 293546
rect 539219 293512 539299 293532
rect 539389 293512 539469 293532
rect 539579 293522 539659 293546
rect 539729 293522 539809 293546
rect 542069 293522 542149 293546
rect 542209 293522 542289 293546
rect 541709 293512 541789 293522
rect 541879 293512 541959 293522
rect 544159 293512 544239 293532
rect 544329 293512 544409 293532
rect 536699 293452 536779 293512
rect 536869 293452 536949 293512
rect 539219 293452 539299 293512
rect 539389 293452 539469 293512
rect 541709 293442 541789 293512
rect 541879 293442 541959 293512
rect 544159 293452 544239 293512
rect 544329 293452 544409 293512
rect 537979 293302 538059 293382
rect 538149 293302 538229 293382
rect 540459 293302 540539 293382
rect 540629 293302 540709 293382
rect 542919 293302 542999 293382
rect 543089 293302 543169 293382
rect 562300 293300 562500 293500
rect 562700 293300 562900 293500
rect 563100 293300 563300 293500
rect 563500 293300 563700 293500
rect 563900 293300 564100 293500
rect 564300 293300 564500 293500
rect 564700 293300 564900 293500
rect 565100 293300 565300 293500
rect 565500 293300 565700 293500
rect 565900 293300 566100 293500
rect 566300 293300 566500 293500
rect 566700 293300 566900 293500
rect 567100 293300 567300 293500
rect 567500 293300 567700 293500
rect 537979 293172 538059 293252
rect 538149 293172 538229 293252
rect 540459 293182 540539 293262
rect 540629 293182 540709 293262
rect 542919 293172 542999 293252
rect 543089 293172 543169 293252
rect 9680 292984 9740 293000
rect 9845 292984 9905 292990
rect 10045 292984 10105 292990
rect 10235 292984 10295 292990
rect 10415 292984 10475 292990
rect 10615 292984 10675 292990
rect 10805 292984 10865 292990
rect 10965 292984 11025 292990
rect 11155 292984 11215 292990
rect 11330 292984 11390 292990
rect 11470 292984 11530 292990
rect 9680 292950 9740 292984
rect 9845 292950 9905 292984
rect 10045 292950 10105 292984
rect 10235 292950 10295 292984
rect 10415 292950 10475 292984
rect 10615 292950 10675 292984
rect 10805 292950 10865 292984
rect 10965 292950 11025 292984
rect 11155 292950 11215 292984
rect 11330 292950 11390 292984
rect 11470 292950 11530 292984
rect 9680 292940 9740 292950
rect 9845 292930 9905 292950
rect 10045 292930 10105 292950
rect 10235 292930 10295 292950
rect 10415 292930 10475 292950
rect 10615 292930 10675 292950
rect 10805 292930 10865 292950
rect 10965 292930 11025 292950
rect 11155 292930 11215 292950
rect 11330 292930 11390 292950
rect 11470 292930 11530 292950
rect 537419 293034 537449 293102
rect 537449 293034 537523 293102
rect 537523 293034 537549 293102
rect 537419 293032 537549 293034
rect 538659 293034 538685 293102
rect 538685 293034 538759 293102
rect 538759 293034 538789 293102
rect 538659 293032 538789 293034
rect 539889 293034 539921 293102
rect 539921 293034 539995 293102
rect 539995 293034 540019 293102
rect 539889 293032 540019 293034
rect 541129 293034 541157 293102
rect 541157 293034 541231 293102
rect 541231 293034 541259 293102
rect 541129 293032 541259 293034
rect 542359 293034 542393 293102
rect 542393 293034 542467 293102
rect 542467 293034 542489 293102
rect 542359 293032 542489 293034
rect 543599 293034 543629 293102
rect 543629 293034 543703 293102
rect 543703 293034 543729 293102
rect 543599 293032 543729 293034
rect 536699 292972 536779 292992
rect 536869 292972 536949 292992
rect 538379 292972 538459 293002
rect 538489 292972 538569 293002
rect 539209 292972 539289 292992
rect 539379 292972 539459 292992
rect 540789 292972 540869 293002
rect 540899 292972 540979 293002
rect 541699 292972 541779 292992
rect 541869 292972 541949 292992
rect 543249 292972 543329 292992
rect 543359 292972 543439 292992
rect 544189 292972 544269 292992
rect 544359 292972 544439 292992
rect 536699 292912 536779 292972
rect 536869 292912 536949 292972
rect 538379 292922 538459 292972
rect 538489 292922 538569 292972
rect 539209 292912 539289 292972
rect 539379 292912 539459 292972
rect 540789 292922 540869 292972
rect 540899 292922 540979 292972
rect 541699 292912 541779 292972
rect 541869 292912 541949 292972
rect 543249 292912 543329 292972
rect 543359 292912 543439 292972
rect 544189 292912 544269 292972
rect 544359 292912 544439 292972
rect 15000 292720 15140 292860
rect 15200 292720 15340 292860
rect 537979 292592 538059 292672
rect 538149 292592 538229 292672
rect 540459 292602 540539 292682
rect 540629 292602 540709 292682
rect 542919 292592 542999 292672
rect 543089 292592 543169 292672
rect 537419 292454 537449 292522
rect 537449 292454 537523 292522
rect 537523 292454 537549 292522
rect 537419 292452 537549 292454
rect 538659 292454 538685 292522
rect 538685 292454 538759 292522
rect 538759 292454 538789 292522
rect 538659 292452 538789 292454
rect 539899 292454 539921 292522
rect 539921 292454 539995 292522
rect 539995 292454 540029 292522
rect 539899 292452 540029 292454
rect 541129 292454 541157 292522
rect 541157 292454 541231 292522
rect 541231 292454 541259 292522
rect 541129 292452 541259 292454
rect 542359 292454 542393 292522
rect 542393 292454 542467 292522
rect 542467 292454 542489 292522
rect 542359 292452 542489 292454
rect 543599 292454 543629 292522
rect 543629 292454 543703 292522
rect 543703 292454 543729 292522
rect 543599 292452 543729 292454
rect 536699 292392 536779 292412
rect 536869 292392 536949 292412
rect 539209 292392 539289 292412
rect 539379 292392 539459 292412
rect 540789 292392 540869 292412
rect 540899 292392 540979 292412
rect 541699 292392 541779 292402
rect 541869 292392 541949 292402
rect 543249 292392 543329 292412
rect 543359 292392 543439 292412
rect 544189 292392 544269 292412
rect 544359 292392 544439 292412
rect 536699 292332 536779 292392
rect 536869 292332 536949 292392
rect 538379 292312 538459 292392
rect 538489 292312 538569 292392
rect 539209 292332 539289 292392
rect 539379 292332 539459 292392
rect 540789 292332 540869 292392
rect 540899 292332 540979 292392
rect 541699 292322 541779 292392
rect 541869 292322 541949 292392
rect 543249 292332 543329 292392
rect 543359 292332 543439 292392
rect 544189 292332 544269 292392
rect 544359 292332 544439 292392
rect 537979 292142 538069 292222
rect 538139 292142 538229 292222
rect 540459 292142 540539 292212
rect 540629 292142 540709 292212
rect 542919 292142 542999 292212
rect 543089 292142 543169 292212
rect 550129 292162 550259 292302
rect 550389 292162 550519 292302
rect 530629 291992 530759 292132
rect 530879 291992 531009 292132
rect 537979 292012 538059 292092
rect 538149 292012 538229 292092
rect 540459 292022 540539 292102
rect 540629 292022 540709 292102
rect 542919 292012 542999 292092
rect 543089 292012 543169 292092
rect 537419 291874 537449 291942
rect 537449 291874 537523 291942
rect 537523 291874 537549 291942
rect 537419 291872 537549 291874
rect 538659 291874 538685 291942
rect 538685 291874 538759 291942
rect 538759 291874 538789 291942
rect 538659 291872 538789 291874
rect 539889 291874 539921 291942
rect 539921 291874 539995 291942
rect 539995 291874 540019 291942
rect 539889 291872 540019 291874
rect 541129 291874 541157 291942
rect 541157 291874 541231 291942
rect 541231 291874 541259 291942
rect 541129 291872 541259 291874
rect 542359 291874 542393 291942
rect 542393 291874 542467 291942
rect 542467 291874 542489 291942
rect 542359 291872 542489 291874
rect 543599 291874 543629 291942
rect 543629 291874 543703 291942
rect 543703 291874 543729 291942
rect 543599 291872 543729 291874
rect 539209 291812 539289 291832
rect 539379 291812 539459 291832
rect 540789 291812 540869 291832
rect 540899 291812 540979 291832
rect 541699 291812 541779 291832
rect 541869 291812 541949 291832
rect 543249 291812 543329 291832
rect 543359 291812 543439 291832
rect 544189 291812 544269 291832
rect 544359 291812 544439 291832
rect 536679 291722 536759 291802
rect 536889 291722 536969 291802
rect 539209 291752 539289 291812
rect 539379 291752 539459 291812
rect 540789 291752 540869 291812
rect 540899 291752 540979 291812
rect 541699 291752 541779 291812
rect 541869 291752 541949 291812
rect 543249 291752 543329 291812
rect 543359 291752 543439 291812
rect 544189 291752 544269 291812
rect 544359 291752 544439 291812
rect 536099 291482 536179 291562
rect 536329 291482 536409 291562
rect 538649 291472 538729 291552
rect 538819 291472 538899 291552
rect 541109 291472 541189 291552
rect 541299 291472 541379 291552
rect 543559 291472 543639 291552
rect 543749 291472 543829 291552
rect 546069 291472 546149 291552
rect 546239 291472 546319 291552
rect 535579 291334 535609 291402
rect 535609 291334 535683 291402
rect 535683 291334 535709 291402
rect 535579 291332 535709 291334
rect 536819 291334 536845 291402
rect 536845 291334 536919 291402
rect 536919 291334 536949 291402
rect 536819 291332 536949 291334
rect 538049 291334 538081 291402
rect 538081 291334 538155 291402
rect 538155 291334 538179 291402
rect 538049 291332 538179 291334
rect 539289 291334 539317 291402
rect 539317 291334 539391 291402
rect 539391 291334 539419 291402
rect 539289 291332 539419 291334
rect 540529 291334 540553 291402
rect 540553 291334 540627 291402
rect 540627 291334 540659 291402
rect 540529 291332 540659 291334
rect 541759 291334 541789 291402
rect 541789 291334 541863 291402
rect 541863 291334 541889 291402
rect 541759 291332 541889 291334
rect 542999 291334 543025 291402
rect 543025 291334 543099 291402
rect 543099 291334 543129 291402
rect 542999 291332 543129 291334
rect 544229 291334 544261 291402
rect 544261 291334 544335 291402
rect 544335 291334 544359 291402
rect 544229 291332 544359 291334
rect 545469 291334 545497 291402
rect 545497 291334 545571 291402
rect 545571 291334 545599 291402
rect 545469 291332 545599 291334
rect 533080 290880 533140 290940
rect 533180 290880 533240 290940
rect 533280 290880 533340 290940
rect 534849 291272 534929 291282
rect 535059 291272 535139 291282
rect 537329 291272 537409 291282
rect 537549 291272 537629 291282
rect 539859 291272 539939 291282
rect 540039 291272 540119 291282
rect 534849 291202 534929 291272
rect 535059 291202 535139 291272
rect 537329 291202 537409 291272
rect 537549 291202 537629 291272
rect 539859 291202 539939 291272
rect 540039 291202 540119 291272
rect 542319 291192 542399 291272
rect 542499 291192 542579 291272
rect 544799 291192 544879 291272
rect 544969 291192 545049 291272
rect 536119 291062 536209 291142
rect 536299 291062 536389 291142
rect 538649 291062 538739 291142
rect 538809 291062 538899 291142
rect 541119 291062 541209 291142
rect 541279 291062 541369 291142
rect 543569 291062 543659 291142
rect 543729 291062 543819 291142
rect 546069 291062 546159 291142
rect 546229 291062 546319 291142
rect 536099 290942 536179 291022
rect 536329 290942 536409 291022
rect 538649 290932 538729 291012
rect 538819 290942 538899 291022
rect 541109 290942 541189 291022
rect 541299 290942 541379 291022
rect 543559 290932 543639 291012
rect 543749 290932 543829 291012
rect 546069 290932 546149 291012
rect 546239 290932 546319 291012
rect 533080 290760 533140 290820
rect 533180 290760 533240 290820
rect 533280 290760 533340 290820
rect 535579 290862 535709 290872
rect 535579 290802 535609 290862
rect 535609 290802 535683 290862
rect 535683 290802 535709 290862
rect 536819 290794 536845 290862
rect 536845 290794 536919 290862
rect 536919 290794 536949 290862
rect 536819 290792 536949 290794
rect 538049 290794 538081 290862
rect 538081 290794 538155 290862
rect 538155 290794 538179 290862
rect 538049 290792 538179 290794
rect 539289 290794 539317 290862
rect 539317 290794 539391 290862
rect 539391 290794 539419 290862
rect 539289 290792 539419 290794
rect 540529 290794 540553 290862
rect 540553 290794 540627 290862
rect 540627 290794 540659 290862
rect 540529 290792 540659 290794
rect 541759 290794 541789 290862
rect 541789 290794 541863 290862
rect 541863 290794 541889 290862
rect 541759 290792 541889 290794
rect 542999 290794 543025 290862
rect 543025 290794 543099 290862
rect 543099 290794 543129 290862
rect 542999 290792 543129 290794
rect 544229 290794 544261 290862
rect 544261 290794 544335 290862
rect 544335 290794 544359 290862
rect 544229 290792 544359 290794
rect 545469 290794 545497 290862
rect 545497 290794 545571 290862
rect 545571 290794 545599 290862
rect 545469 290792 545599 290794
rect 533080 290660 533140 290720
rect 533180 290660 533240 290720
rect 533280 290660 533340 290720
rect 534849 290732 534929 290742
rect 535059 290732 535139 290742
rect 537329 290732 537409 290742
rect 537549 290732 537629 290742
rect 539859 290732 539939 290742
rect 540049 290732 540129 290742
rect 534849 290662 534929 290732
rect 535059 290662 535139 290732
rect 537329 290662 537409 290732
rect 537549 290662 537629 290732
rect 539859 290662 539939 290732
rect 540049 290662 540129 290732
rect 542319 290652 542399 290732
rect 542499 290652 542579 290732
rect 544799 290652 544879 290732
rect 544969 290652 545049 290732
rect 533080 290520 533140 290580
rect 533180 290520 533240 290580
rect 533280 290520 533340 290580
rect 533080 290420 533140 290480
rect 533180 290420 533240 290480
rect 533280 290420 533340 290480
rect 533080 290320 533140 290380
rect 533180 290320 533240 290380
rect 533280 290320 533340 290380
rect 536099 290402 536179 290482
rect 536329 290402 536409 290482
rect 538639 290392 538719 290472
rect 538809 290392 538889 290472
rect 541109 290392 541189 290472
rect 541289 290392 541369 290472
rect 543559 290392 543639 290472
rect 543749 290392 543829 290472
rect 546069 290392 546149 290472
rect 546239 290392 546319 290472
rect 533080 290220 533140 290280
rect 533180 290220 533240 290280
rect 533280 290220 533340 290280
rect 535579 290254 535609 290322
rect 535609 290254 535683 290322
rect 535683 290254 535709 290322
rect 535579 290252 535709 290254
rect 536819 290254 536845 290322
rect 536845 290254 536919 290322
rect 536919 290254 536949 290322
rect 536819 290252 536949 290254
rect 538049 290254 538081 290322
rect 538081 290254 538155 290322
rect 538155 290254 538179 290322
rect 538049 290252 538179 290254
rect 539289 290254 539317 290322
rect 539317 290254 539391 290322
rect 539391 290254 539419 290322
rect 539289 290252 539419 290254
rect 540529 290254 540553 290322
rect 540553 290254 540627 290322
rect 540627 290254 540659 290322
rect 540529 290252 540659 290254
rect 541759 290254 541789 290322
rect 541789 290254 541863 290322
rect 541863 290254 541889 290322
rect 541759 290252 541889 290254
rect 542999 290254 543025 290322
rect 543025 290254 543099 290322
rect 543099 290254 543129 290322
rect 542999 290252 543129 290254
rect 544229 290254 544261 290322
rect 544261 290254 544335 290322
rect 544335 290254 544359 290322
rect 544229 290252 544359 290254
rect 545469 290254 545497 290322
rect 545497 290254 545571 290322
rect 545571 290254 545599 290322
rect 545469 290252 545599 290254
rect 534849 290192 534929 290202
rect 535059 290192 535139 290202
rect 537319 290192 537399 290202
rect 537559 290192 537639 290202
rect 539859 290192 539939 290202
rect 540039 290192 540119 290202
rect 534849 290122 534929 290192
rect 535059 290122 535139 290192
rect 537319 290122 537399 290192
rect 537559 290122 537639 290192
rect 539859 290122 539939 290192
rect 540039 290122 540119 290192
rect 542329 290112 542409 290192
rect 542499 290112 542579 290192
rect 544799 290112 544879 290192
rect 544969 290112 545049 290192
rect 536119 289982 536209 290062
rect 536299 289992 536389 290072
rect 538649 289982 538739 290062
rect 538809 289982 538899 290062
rect 541119 289982 541209 290062
rect 541279 289982 541369 290062
rect 543569 289982 543659 290062
rect 543729 289982 543819 290062
rect 546069 289982 546159 290062
rect 546229 289982 546319 290062
rect 536099 289852 536179 289932
rect 536329 289852 536409 289932
rect 538629 289862 538709 289942
rect 538819 289862 538899 289942
rect 541109 289852 541189 289932
rect 541299 289852 541379 289932
rect 543559 289852 543639 289932
rect 543749 289852 543829 289932
rect 546069 289844 546149 289922
rect 546239 289844 546319 289922
rect 546069 289842 546149 289844
rect 546239 289842 546319 289844
rect 535579 289714 535609 289782
rect 535609 289714 535683 289782
rect 535683 289714 535709 289782
rect 535579 289712 535709 289714
rect 536819 289714 536845 289782
rect 536845 289714 536919 289782
rect 536919 289714 536949 289782
rect 536819 289712 536949 289714
rect 538049 289714 538081 289782
rect 538081 289714 538155 289782
rect 538155 289714 538179 289782
rect 538049 289712 538179 289714
rect 539289 289714 539317 289782
rect 539317 289714 539391 289782
rect 539391 289714 539419 289782
rect 539289 289712 539419 289714
rect 540529 289714 540553 289782
rect 540553 289714 540627 289782
rect 540627 289714 540659 289782
rect 540529 289712 540659 289714
rect 541759 289714 541789 289782
rect 541789 289714 541863 289782
rect 541863 289714 541889 289782
rect 541759 289712 541889 289714
rect 542999 289714 543025 289782
rect 543025 289714 543099 289782
rect 543099 289714 543129 289782
rect 542999 289712 543129 289714
rect 544229 289714 544261 289782
rect 544261 289714 544335 289782
rect 544335 289714 544359 289782
rect 544229 289712 544359 289714
rect 545469 289714 545497 289782
rect 545497 289714 545571 289782
rect 545571 289714 545599 289782
rect 545469 289712 545599 289714
rect 534849 289652 534929 289662
rect 535059 289652 535139 289662
rect 539859 289652 539939 289662
rect 540049 289652 540129 289662
rect 534849 289582 534929 289652
rect 535059 289582 535139 289652
rect 537319 289572 537399 289652
rect 537559 289572 537639 289652
rect 539859 289582 539939 289652
rect 540049 289582 540129 289652
rect 542319 289572 542399 289652
rect 542509 289572 542589 289652
rect 544799 289562 544879 289642
rect 544969 289562 545049 289642
rect 531759 289122 531849 289252
rect 531969 289122 532059 289252
rect 549069 289152 549139 289242
rect 549229 289152 549299 289242
rect 536819 289064 536949 289132
rect 538049 289064 538179 289122
rect 538379 289064 538459 289132
rect 538489 289064 538569 289132
rect 539289 289064 539419 289122
rect 540529 289064 540659 289122
rect 540789 289064 540869 289132
rect 540899 289064 540979 289132
rect 541759 289064 541889 289122
rect 542999 289072 543129 289142
rect 543249 289064 543329 289142
rect 543359 289064 543439 289142
rect 544229 289064 544359 289122
rect 536819 289062 536949 289064
rect 538049 289052 538179 289064
rect 538379 289052 538459 289064
rect 538489 289052 538569 289064
rect 539289 289052 539419 289064
rect 540529 289052 540659 289064
rect 540789 289052 540869 289064
rect 540899 289052 540979 289064
rect 541759 289052 541889 289064
rect 543249 289062 543329 289064
rect 543359 289062 543439 289064
rect 544229 289052 544359 289064
rect 541769 288872 541859 288882
rect 541909 288872 541999 288882
rect 536759 288782 536849 288862
rect 536899 288782 536989 288862
rect 541769 288802 541859 288872
rect 541909 288802 541999 288872
rect 538279 288662 538389 288772
rect 539139 288662 539249 288772
rect 540349 288662 540459 288772
rect 541199 288662 541309 288772
rect 536759 288564 536849 288632
rect 536899 288564 536989 288632
rect 542769 288662 542879 288772
rect 543649 288662 543759 288772
rect 541769 288564 541859 288622
rect 541909 288564 541999 288622
rect 536759 288552 536849 288564
rect 536899 288552 536989 288564
rect 541769 288542 541859 288564
rect 541909 288542 541999 288564
rect 539579 288372 539659 288392
rect 539729 288372 539809 288392
rect 542059 288372 542139 288392
rect 542199 288372 542279 288392
rect 537089 288292 537169 288372
rect 537239 288292 537319 288372
rect 539579 288312 539659 288372
rect 539729 288312 539809 288372
rect 542059 288312 542139 288372
rect 542199 288312 542279 288372
rect 537539 288064 537619 288142
rect 537649 288064 537729 288142
rect 539949 288064 540029 288112
rect 542399 288064 542479 288132
rect 542519 288064 542599 288132
rect 543599 288064 543679 288122
rect 537539 288062 537619 288064
rect 537649 288062 537729 288064
rect 539949 288032 540029 288064
rect 542399 288052 542479 288064
rect 542519 288052 542599 288064
rect 543599 288042 543679 288064
rect 538719 287882 538799 287962
rect 541129 287882 541209 287962
rect 537459 287772 537539 287782
rect 542349 287772 542429 287782
rect 537459 287702 537539 287772
rect 542349 287702 542429 287772
rect 537569 287562 537679 287652
rect 542479 287562 542589 287652
rect 539949 287444 540029 287492
rect 543599 287444 543679 287502
rect 539949 287412 540029 287444
rect 543599 287422 543679 287444
rect 538109 287262 538165 287342
rect 538165 287262 538199 287342
rect 538229 287262 538319 287342
rect 538719 287262 538799 287342
rect 540559 287262 540601 287342
rect 540601 287262 540635 287342
rect 540635 287262 540649 287342
rect 540679 287262 540769 287342
rect 541129 287262 541209 287342
rect 542989 287262 543037 287342
rect 543037 287262 543071 287342
rect 543071 287262 543079 287342
rect 543109 287262 543199 287342
rect 537459 287152 537539 287162
rect 542349 287152 542429 287162
rect 537459 287082 537539 287152
rect 542349 287082 542429 287152
rect 539339 286844 539429 286912
rect 544219 286852 544309 286932
rect 539339 286832 539429 286844
rect 538109 286662 538199 286742
rect 538229 286662 538319 286742
rect 540559 286662 540649 286742
rect 540679 286662 540769 286742
rect 542989 286662 543079 286742
rect 543109 286662 543199 286742
rect 536759 286552 536849 286582
rect 536899 286552 536989 286582
rect 541769 286552 541859 286582
rect 541909 286552 541999 286582
rect 536759 286502 536849 286552
rect 536899 286502 536989 286552
rect 541769 286502 541859 286552
rect 541909 286502 541999 286552
rect 537509 286352 537629 286452
rect 538729 286352 538849 286452
rect 539939 286352 540059 286452
rect 539339 286244 539429 286312
rect 541159 286352 541279 286452
rect 542389 286342 542509 286442
rect 543599 286352 543719 286452
rect 544219 286252 544309 286332
rect 572750 288744 572810 288764
rect 572890 288744 572950 288764
rect 573065 288744 573125 288764
rect 573255 288744 573315 288764
rect 573415 288744 573475 288764
rect 573605 288744 573665 288764
rect 573805 288744 573865 288764
rect 573985 288744 574045 288764
rect 574175 288744 574235 288764
rect 574375 288744 574435 288764
rect 574540 288744 574600 288754
rect 572750 288710 572810 288744
rect 572890 288710 572950 288744
rect 573065 288710 573125 288744
rect 573255 288710 573315 288744
rect 573415 288710 573475 288744
rect 573605 288710 573665 288744
rect 573805 288710 573865 288744
rect 573985 288710 574045 288744
rect 574175 288710 574235 288744
rect 574375 288710 574435 288744
rect 574540 288710 574600 288744
rect 572750 288704 572810 288710
rect 572890 288704 572950 288710
rect 573065 288704 573125 288710
rect 573255 288704 573315 288710
rect 573415 288704 573475 288710
rect 573605 288704 573665 288710
rect 573805 288704 573865 288710
rect 573985 288704 574045 288710
rect 574175 288704 574235 288710
rect 574375 288704 574435 288710
rect 574540 288694 574600 288710
rect 578360 288597 578440 288600
rect 572750 288548 572810 288564
rect 572890 288548 572950 288564
rect 573065 288548 573125 288564
rect 573255 288548 573315 288564
rect 573415 288548 573475 288564
rect 573605 288548 573665 288564
rect 573805 288548 573865 288564
rect 573985 288548 574045 288564
rect 574175 288548 574235 288564
rect 574375 288548 574435 288564
rect 574540 288548 574600 288564
rect 578360 288563 578362 288597
rect 578362 288563 578440 288597
rect 572750 288514 572810 288548
rect 572890 288514 572950 288548
rect 573065 288514 573125 288548
rect 573255 288514 573315 288548
rect 573415 288514 573475 288548
rect 573605 288514 573665 288548
rect 573805 288514 573865 288548
rect 573985 288514 574045 288548
rect 574175 288514 574235 288548
rect 574375 288514 574435 288548
rect 574540 288514 574600 288548
rect 572750 288504 572810 288514
rect 572890 288504 572950 288514
rect 573065 288504 573125 288514
rect 573255 288504 573315 288514
rect 573415 288504 573475 288514
rect 573605 288504 573665 288514
rect 573805 288504 573865 288514
rect 573985 288504 574045 288514
rect 574175 288504 574235 288514
rect 574375 288504 574435 288514
rect 574540 288504 574600 288514
rect 578360 288520 578440 288563
rect 578540 288520 578620 288600
rect 578360 288401 578440 288440
rect 572750 288352 572810 288364
rect 572890 288352 572950 288364
rect 573065 288352 573125 288364
rect 573255 288352 573315 288364
rect 573415 288352 573475 288364
rect 573605 288352 573665 288364
rect 573805 288352 573865 288364
rect 573985 288352 574045 288364
rect 574175 288352 574235 288364
rect 574375 288352 574435 288364
rect 574540 288352 574600 288364
rect 578360 288367 578362 288401
rect 578362 288367 578440 288401
rect 578360 288360 578440 288367
rect 578540 288360 578620 288440
rect 572750 288318 572810 288352
rect 572890 288318 572950 288352
rect 573065 288318 573125 288352
rect 573255 288318 573315 288352
rect 573415 288318 573475 288352
rect 573605 288318 573665 288352
rect 573805 288318 573865 288352
rect 573985 288318 574045 288352
rect 574175 288318 574235 288352
rect 574375 288318 574435 288352
rect 574540 288318 574600 288352
rect 572750 288304 572810 288318
rect 572890 288304 572950 288318
rect 573065 288304 573125 288318
rect 573255 288304 573315 288318
rect 573415 288304 573475 288318
rect 573605 288304 573665 288318
rect 573805 288304 573865 288318
rect 573985 288304 574045 288318
rect 574175 288304 574235 288318
rect 574375 288304 574435 288318
rect 574540 288304 574600 288318
rect 578360 288205 578440 288280
rect 572750 288156 572810 288174
rect 572890 288156 572950 288174
rect 573065 288156 573125 288174
rect 573255 288156 573315 288174
rect 573415 288156 573475 288174
rect 573605 288156 573665 288174
rect 573805 288156 573865 288174
rect 573985 288156 574045 288174
rect 574175 288156 574235 288174
rect 574375 288156 574435 288174
rect 574540 288156 574600 288174
rect 578360 288200 578362 288205
rect 578362 288200 578440 288205
rect 578540 288200 578620 288280
rect 572750 288122 572810 288156
rect 572890 288122 572950 288156
rect 573065 288122 573125 288156
rect 573255 288122 573315 288156
rect 573415 288122 573475 288156
rect 573605 288122 573665 288156
rect 573805 288122 573865 288156
rect 573985 288122 574045 288156
rect 574175 288122 574235 288156
rect 574375 288122 574435 288156
rect 574540 288122 574600 288156
rect 572750 288114 572810 288122
rect 572890 288114 572950 288122
rect 573065 288114 573125 288122
rect 573255 288114 573315 288122
rect 573415 288114 573475 288122
rect 573605 288114 573665 288122
rect 573805 288114 573865 288122
rect 573985 288114 574045 288122
rect 574175 288114 574235 288122
rect 574375 288114 574435 288122
rect 574540 288114 574600 288122
rect 578360 288020 578440 288100
rect 578540 288020 578620 288100
rect 572750 287960 572810 287974
rect 572890 287960 572950 287974
rect 573065 287960 573125 287974
rect 573255 287960 573315 287974
rect 573415 287960 573475 287974
rect 573605 287960 573665 287974
rect 573805 287960 573865 287974
rect 573985 287960 574045 287974
rect 574175 287960 574235 287974
rect 574375 287960 574435 287974
rect 574540 287960 574600 287974
rect 572750 287926 572810 287960
rect 572890 287926 572950 287960
rect 573065 287926 573125 287960
rect 573255 287926 573315 287960
rect 573415 287926 573475 287960
rect 573605 287926 573665 287960
rect 573805 287926 573865 287960
rect 573985 287926 574045 287960
rect 574175 287926 574235 287960
rect 574375 287926 574435 287960
rect 574540 287926 574600 287960
rect 572750 287914 572810 287926
rect 572890 287914 572950 287926
rect 573065 287914 573125 287926
rect 573255 287914 573315 287926
rect 573415 287914 573475 287926
rect 573605 287914 573665 287926
rect 573805 287914 573865 287926
rect 573985 287914 574045 287926
rect 574175 287914 574235 287926
rect 574375 287914 574435 287926
rect 574540 287914 574600 287926
rect 578360 287860 578440 287940
rect 578540 287860 578620 287940
rect 572750 287764 572810 287774
rect 572890 287764 572950 287774
rect 573065 287764 573125 287774
rect 573255 287764 573315 287774
rect 573415 287764 573475 287774
rect 573605 287764 573665 287774
rect 573805 287764 573865 287774
rect 573985 287764 574045 287774
rect 574175 287764 574235 287774
rect 574375 287764 574435 287774
rect 574540 287764 574600 287774
rect 572750 287730 572810 287764
rect 572890 287730 572950 287764
rect 573065 287730 573125 287764
rect 573255 287730 573315 287764
rect 573415 287730 573475 287764
rect 573605 287730 573665 287764
rect 573805 287730 573865 287764
rect 573985 287730 574045 287764
rect 574175 287730 574235 287764
rect 574375 287730 574435 287764
rect 574540 287730 574600 287764
rect 572750 287714 572810 287730
rect 572890 287714 572950 287730
rect 573065 287714 573125 287730
rect 573255 287714 573315 287730
rect 573415 287714 573475 287730
rect 573605 287714 573665 287730
rect 573805 287714 573865 287730
rect 573985 287714 574045 287730
rect 574175 287714 574235 287730
rect 574375 287714 574435 287730
rect 574540 287714 574600 287730
rect 539339 286232 539429 286244
rect 538109 286062 538199 286142
rect 538229 286062 538319 286142
rect 540420 286056 540508 286146
rect 540559 286062 540649 286142
rect 540679 286062 540769 286142
rect 542989 286062 543079 286142
rect 543109 286062 543199 286142
rect 557700 286000 557900 286200
rect 558100 286000 558300 286200
rect 558500 286000 558700 286200
rect 558900 286000 559100 286200
rect 559300 286000 559500 286200
rect 536759 285952 536849 285962
rect 536899 285952 536989 285962
rect 541769 285952 541859 285982
rect 541909 285952 541999 285982
rect 536759 285882 536849 285952
rect 536899 285882 536989 285952
rect 541769 285902 541859 285952
rect 541909 285902 541999 285952
rect 557700 285600 557900 285800
rect 558100 285600 558300 285800
rect 558500 285600 558700 285800
rect 558900 285600 559100 285800
rect 559300 285600 559500 285800
rect 537384 285318 537544 285478
rect 538444 285318 538604 285478
rect 539904 285318 540064 285478
rect 541124 285318 541284 285478
rect 542604 285318 542764 285478
rect 543604 285318 543764 285478
rect 538884 285088 538954 285158
rect 539104 285088 539174 285158
rect 542064 285088 542134 285158
rect 542304 285088 542374 285158
rect 557700 285200 557900 285400
rect 558100 285200 558300 285400
rect 558500 285200 558700 285400
rect 558900 285200 559100 285400
rect 559300 285200 559500 285400
rect 537384 284738 537544 284898
rect 538444 284738 538604 284898
rect 539904 284738 540064 284898
rect 541124 284738 541284 284898
rect 542604 284738 542764 284898
rect 543604 284738 543764 284898
rect 557700 284800 557900 285000
rect 558100 284800 558300 285000
rect 558500 284800 558700 285000
rect 558900 284800 559100 285000
rect 559300 284800 559500 285000
rect 538884 284498 538954 284568
rect 539104 284498 539174 284568
rect 542064 284498 542134 284568
rect 542304 284498 542374 284568
rect 540044 284388 540114 284408
rect 540154 284388 540224 284408
rect 540984 284388 541054 284408
rect 541094 284388 541164 284408
rect 540044 284338 540114 284388
rect 540154 284338 540224 284388
rect 540984 284338 541054 284388
rect 541094 284338 541164 284388
rect 557700 284400 557900 284600
rect 558100 284400 558300 284600
rect 558500 284400 558700 284600
rect 558900 284400 559100 284600
rect 559300 284400 559500 284600
rect 557700 284000 557900 284200
rect 558100 284000 558300 284200
rect 558500 284000 558700 284200
rect 558900 284000 559100 284200
rect 559300 284000 559500 284200
rect 540410 283890 540470 283926
rect 540410 283866 540470 283890
rect 540510 283866 540570 283926
rect 540610 283866 540670 283926
rect 540710 283890 540770 283926
rect 540710 283866 540722 283890
rect 540722 283866 540770 283890
rect 540044 283828 540114 283838
rect 540044 283768 540062 283828
rect 540062 283768 540096 283828
rect 540096 283768 540114 283828
rect 540154 283828 540224 283838
rect 540984 283828 541054 283848
rect 540154 283768 540170 283828
rect 540170 283768 540204 283828
rect 540204 283768 540224 283828
rect 540984 283778 540998 283828
rect 540998 283778 541032 283828
rect 541032 283778 541054 283828
rect 541094 283828 541164 283848
rect 541094 283778 541106 283828
rect 541106 283778 541140 283828
rect 541140 283778 541164 283828
rect 557700 283600 557900 283800
rect 558100 283600 558300 283800
rect 558500 283600 558700 283800
rect 558900 283600 559100 283800
rect 559300 283600 559500 283800
rect 539764 283368 539984 283518
rect 540284 283368 540504 283518
rect 540704 283368 540924 283518
rect 541254 283368 541474 283518
rect 538884 283238 538954 283308
rect 539094 283238 539164 283308
rect 542064 283258 542134 283328
rect 542304 283258 542374 283328
rect 538884 283148 538954 283218
rect 539094 283148 539164 283218
rect 542064 283168 542134 283238
rect 542304 283168 542374 283238
rect 557700 283200 557900 283400
rect 558100 283200 558300 283400
rect 558500 283200 558700 283400
rect 558900 283200 559100 283400
rect 559300 283200 559500 283400
rect 540044 283073 540114 283088
rect 540154 283073 540224 283088
rect 540984 283073 541054 283088
rect 541094 283073 541164 283088
rect 540044 283018 540114 283073
rect 540154 283018 540224 283073
rect 540984 283018 541054 283073
rect 541094 283018 541164 283073
rect 537404 282828 537584 282958
rect 538544 282828 538724 282958
rect 539524 282838 539704 282968
rect 540294 282838 540474 282968
rect 540734 282838 540914 282968
rect 541454 282828 541634 282958
rect 542524 282838 542704 282968
rect 543524 282838 543704 282968
rect 557700 282800 557900 283000
rect 558100 282800 558300 283000
rect 558500 282800 558700 283000
rect 558900 282800 559100 283000
rect 559300 282800 559500 283000
rect 538884 282740 538954 282788
rect 539104 282740 539174 282788
rect 542064 282740 542134 282788
rect 542304 282740 542374 282788
rect 538884 282718 538954 282740
rect 539104 282718 539174 282740
rect 542064 282718 542134 282740
rect 542304 282718 542374 282740
rect 540044 282568 540114 282638
rect 540154 282568 540224 282638
rect 540984 282568 541054 282638
rect 541094 282568 541164 282638
rect 557700 282400 557900 282600
rect 558100 282400 558300 282600
rect 558500 282400 558700 282600
rect 558900 282400 559100 282600
rect 559300 282400 559500 282600
rect 567900 281100 568100 281300
rect 572770 281264 572830 281284
rect 572910 281264 572970 281284
rect 573085 281264 573145 281284
rect 573275 281264 573335 281284
rect 573435 281264 573495 281284
rect 573625 281264 573685 281284
rect 573825 281264 573885 281284
rect 574005 281264 574065 281284
rect 574195 281264 574255 281284
rect 574395 281264 574455 281284
rect 574560 281264 574620 281274
rect 572770 281230 572830 281264
rect 572910 281230 572970 281264
rect 573085 281230 573145 281264
rect 573275 281230 573335 281264
rect 573435 281230 573495 281264
rect 573625 281230 573685 281264
rect 573825 281230 573885 281264
rect 574005 281230 574065 281264
rect 574195 281230 574255 281264
rect 574395 281230 574455 281264
rect 574560 281230 574620 281264
rect 572770 281224 572830 281230
rect 572910 281224 572970 281230
rect 573085 281224 573145 281230
rect 573275 281224 573335 281230
rect 573435 281224 573495 281230
rect 573625 281224 573685 281230
rect 573825 281224 573885 281230
rect 574005 281224 574065 281230
rect 574195 281224 574255 281230
rect 574395 281224 574455 281230
rect 574560 281214 574620 281230
rect 537364 280938 537484 281058
rect 543734 280938 543854 281058
rect 567900 280800 568100 281000
rect 13190 280430 13260 280500
rect 13080 280320 13150 280390
rect 567900 280500 568100 280700
rect 572770 281068 572830 281084
rect 572910 281068 572970 281084
rect 573085 281068 573145 281084
rect 573275 281068 573335 281084
rect 573435 281068 573495 281084
rect 573625 281068 573685 281084
rect 573825 281068 573885 281084
rect 574005 281068 574065 281084
rect 574195 281068 574255 281084
rect 574395 281068 574455 281084
rect 574560 281068 574620 281084
rect 572770 281034 572830 281068
rect 572910 281034 572970 281068
rect 573085 281034 573145 281068
rect 573275 281034 573335 281068
rect 573435 281034 573495 281068
rect 573625 281034 573685 281068
rect 573825 281034 573885 281068
rect 574005 281034 574065 281068
rect 574195 281034 574255 281068
rect 574395 281034 574455 281068
rect 574560 281034 574620 281068
rect 572770 281024 572830 281034
rect 572910 281024 572970 281034
rect 573085 281024 573145 281034
rect 573275 281024 573335 281034
rect 573435 281024 573495 281034
rect 573625 281024 573685 281034
rect 573825 281024 573885 281034
rect 574005 281024 574065 281034
rect 574195 281024 574255 281034
rect 574395 281024 574455 281034
rect 574560 281024 574620 281034
rect 572770 280872 572830 280884
rect 572910 280872 572970 280884
rect 573085 280872 573145 280884
rect 573275 280872 573335 280884
rect 573435 280872 573495 280884
rect 573625 280872 573685 280884
rect 573825 280872 573885 280884
rect 574005 280872 574065 280884
rect 574195 280872 574255 280884
rect 574395 280872 574455 280884
rect 574560 280872 574620 280884
rect 572770 280838 572830 280872
rect 572910 280838 572970 280872
rect 573085 280838 573145 280872
rect 573275 280838 573335 280872
rect 573435 280838 573495 280872
rect 573625 280838 573685 280872
rect 573825 280838 573885 280872
rect 574005 280838 574065 280872
rect 574195 280838 574255 280872
rect 574395 280838 574455 280872
rect 574560 280838 574620 280872
rect 572770 280824 572830 280838
rect 572910 280824 572970 280838
rect 573085 280824 573145 280838
rect 573275 280824 573335 280838
rect 573435 280824 573495 280838
rect 573625 280824 573685 280838
rect 573825 280824 573885 280838
rect 574005 280824 574065 280838
rect 574195 280824 574255 280838
rect 574395 280824 574455 280838
rect 574560 280824 574620 280838
rect 572770 280676 572830 280694
rect 572910 280676 572970 280694
rect 573085 280676 573145 280694
rect 573275 280676 573335 280694
rect 573435 280676 573495 280694
rect 573625 280676 573685 280694
rect 573825 280676 573885 280694
rect 574005 280676 574065 280694
rect 574195 280676 574255 280694
rect 574395 280676 574455 280694
rect 574560 280676 574620 280694
rect 572770 280642 572830 280676
rect 572910 280642 572970 280676
rect 573085 280642 573145 280676
rect 573275 280642 573335 280676
rect 573435 280642 573495 280676
rect 573625 280642 573685 280676
rect 573825 280642 573885 280676
rect 574005 280642 574065 280676
rect 574195 280642 574255 280676
rect 574395 280642 574455 280676
rect 574560 280642 574620 280676
rect 572770 280634 572830 280642
rect 572910 280634 572970 280642
rect 573085 280634 573145 280642
rect 573275 280634 573335 280642
rect 573435 280634 573495 280642
rect 573625 280634 573685 280642
rect 573825 280634 573885 280642
rect 574005 280634 574065 280642
rect 574195 280634 574255 280642
rect 574395 280634 574455 280642
rect 574560 280634 574620 280642
rect 572770 280480 572830 280494
rect 572910 280480 572970 280494
rect 573085 280480 573145 280494
rect 573275 280480 573335 280494
rect 573435 280480 573495 280494
rect 573625 280480 573685 280494
rect 573825 280480 573885 280494
rect 574005 280480 574065 280494
rect 574195 280480 574255 280494
rect 574395 280480 574455 280494
rect 574560 280480 574620 280494
rect 572770 280446 572830 280480
rect 572910 280446 572970 280480
rect 573085 280446 573145 280480
rect 573275 280446 573335 280480
rect 573435 280446 573495 280480
rect 573625 280446 573685 280480
rect 573825 280446 573885 280480
rect 574005 280446 574065 280480
rect 574195 280446 574255 280480
rect 574395 280446 574455 280480
rect 574560 280446 574620 280480
rect 567900 280200 568100 280400
rect 572770 280434 572830 280446
rect 572910 280434 572970 280446
rect 573085 280434 573145 280446
rect 573275 280434 573335 280446
rect 573435 280434 573495 280446
rect 573625 280434 573685 280446
rect 573825 280434 573885 280446
rect 574005 280434 574065 280446
rect 574195 280434 574255 280446
rect 574395 280434 574455 280446
rect 574560 280434 574620 280446
rect 572770 280284 572830 280294
rect 572910 280284 572970 280294
rect 573085 280284 573145 280294
rect 573275 280284 573335 280294
rect 573435 280284 573495 280294
rect 573625 280284 573685 280294
rect 573825 280284 573885 280294
rect 574005 280284 574065 280294
rect 574195 280284 574255 280294
rect 574395 280284 574455 280294
rect 574560 280284 574620 280294
rect 572770 280250 572830 280284
rect 572910 280250 572970 280284
rect 573085 280250 573145 280284
rect 573275 280250 573335 280284
rect 573435 280250 573495 280284
rect 573625 280250 573685 280284
rect 573825 280250 573885 280284
rect 574005 280250 574065 280284
rect 574195 280250 574255 280284
rect 574395 280250 574455 280284
rect 574560 280250 574620 280284
rect 572770 280234 572830 280250
rect 572910 280234 572970 280250
rect 573085 280234 573145 280250
rect 573275 280234 573335 280250
rect 573435 280234 573495 280250
rect 573625 280234 573685 280250
rect 573825 280234 573885 280250
rect 574005 280234 574065 280250
rect 574195 280234 574255 280250
rect 574395 280234 574455 280250
rect 574560 280234 574620 280250
rect 14540 278370 14640 278550
rect 14540 277950 14640 278130
rect 537364 277938 537484 278058
rect 543734 277938 543854 278058
rect 12840 275834 12910 275850
rect 13080 275834 13150 275850
rect 12840 275800 12910 275834
rect 13080 275800 13150 275834
rect 12840 275780 12910 275800
rect 13080 275780 13150 275800
rect 31020 275900 31260 276140
rect 32740 275900 32980 276140
rect 34460 275900 34700 276140
rect 35940 275900 36180 276140
rect 37660 275900 37900 276140
rect 39260 275900 39500 276140
rect 40980 275900 41220 276140
rect 42580 275900 42820 276140
rect 44300 275900 44540 276140
rect 44780 275900 45020 276140
rect 13450 275676 13520 275700
rect 13690 275676 13760 275700
rect 13450 275642 13520 275676
rect 13690 275642 13760 275676
rect 13450 275630 13520 275642
rect 13690 275630 13760 275642
rect 12840 275518 12910 275540
rect 13080 275518 13150 275540
rect 12840 275484 12910 275518
rect 13080 275484 13150 275518
rect 12840 275470 12910 275484
rect 13080 275470 13150 275484
rect 13450 275360 13520 275380
rect 13690 275360 13760 275380
rect 13450 275326 13520 275360
rect 13690 275326 13760 275360
rect 13450 275310 13520 275326
rect 13690 275310 13760 275326
rect 12840 275202 12910 275220
rect 13080 275202 13150 275220
rect 12840 275168 12910 275202
rect 13080 275168 13150 275202
rect 12840 275150 12910 275168
rect 13080 275150 13150 275168
rect 17700 275200 17800 275300
rect 18000 275200 18200 275300
rect 18400 275200 18500 275300
rect 13450 275044 13520 275060
rect 13690 275044 13760 275060
rect 13450 275010 13520 275044
rect 13690 275010 13760 275044
rect 13450 274990 13520 275010
rect 13690 274990 13760 275010
rect 12840 274886 12910 274900
rect 13080 274886 13150 274900
rect 12840 274852 12910 274886
rect 13080 274852 13150 274886
rect 12840 274830 12910 274852
rect 13080 274830 13150 274852
rect 13450 274728 13520 274750
rect 13690 274728 13760 274750
rect 13450 274694 13520 274728
rect 13690 274694 13760 274728
rect 13450 274680 13520 274694
rect 13690 274680 13760 274694
rect 13860 274666 13940 274720
rect 12840 274570 12910 274590
rect 13080 274570 13150 274590
rect 13860 274640 13882 274666
rect 13882 274640 13940 274666
rect 12840 274536 12910 274570
rect 13080 274536 13150 274570
rect 12840 274520 12910 274536
rect 13080 274520 13150 274536
rect 13450 274412 13520 274430
rect 13690 274412 13760 274430
rect 13450 274378 13520 274412
rect 13690 274378 13760 274412
rect 13450 274360 13520 274378
rect 13690 274360 13760 274378
rect 12360 273060 12618 273330
rect 12618 273060 12630 273330
rect 12360 272010 12618 272280
rect 12618 272010 12630 272280
rect 12840 274254 12910 274270
rect 13080 274254 13150 274270
rect 12840 274220 12910 274254
rect 13080 274220 13150 274254
rect 12840 274200 12910 274220
rect 13080 274200 13150 274220
rect 13450 274096 13520 274110
rect 13690 274096 13760 274110
rect 13450 274062 13520 274096
rect 13690 274062 13760 274096
rect 13450 274040 13520 274062
rect 13690 274040 13760 274062
rect 12840 273938 12910 273960
rect 13080 273938 13150 273960
rect 12840 273904 12910 273938
rect 13080 273904 13150 273938
rect 12840 273890 12910 273904
rect 13080 273890 13150 273904
rect 13450 273780 13520 273800
rect 13690 273780 13760 273800
rect 13450 273746 13520 273780
rect 13690 273746 13760 273780
rect 13450 273730 13520 273746
rect 13690 273730 13760 273746
rect 12840 273622 12910 273640
rect 13080 273622 13150 273640
rect 12840 273588 12910 273622
rect 13080 273588 13150 273622
rect 12840 273570 12910 273588
rect 13080 273570 13150 273588
rect 13450 273464 13520 273480
rect 13690 273464 13760 273480
rect 13450 273430 13520 273464
rect 13690 273430 13760 273464
rect 13450 273410 13520 273430
rect 13690 273410 13760 273430
rect 12840 273306 12910 273320
rect 13080 273306 13150 273320
rect 12840 273272 12910 273306
rect 13080 273272 13150 273306
rect 12840 273250 12910 273272
rect 13080 273250 13150 273272
rect 13450 273148 13520 273170
rect 13690 273148 13760 273170
rect 13450 273114 13520 273148
rect 13690 273114 13760 273148
rect 13450 273100 13520 273114
rect 13690 273100 13760 273114
rect 12840 272990 12910 273010
rect 13080 272990 13150 273010
rect 12840 272956 12910 272990
rect 13080 272956 13150 272990
rect 12840 272940 12910 272956
rect 13080 272940 13150 272956
rect 13450 272832 13520 272850
rect 13690 272832 13760 272850
rect 13450 272798 13520 272832
rect 13690 272798 13760 272832
rect 13450 272780 13520 272798
rect 13690 272780 13760 272798
rect 12840 272674 12910 272690
rect 13080 272674 13150 272690
rect 12840 272640 12910 272674
rect 13080 272640 13150 272674
rect 12840 272620 12910 272640
rect 13080 272620 13150 272640
rect 13450 272516 13520 272530
rect 13690 272516 13760 272530
rect 13450 272482 13520 272516
rect 13690 272482 13760 272516
rect 13450 272460 13520 272482
rect 13690 272460 13760 272482
rect 12840 272358 12910 272380
rect 13080 272358 13150 272380
rect 12840 272324 12910 272358
rect 13080 272324 13150 272358
rect 12840 272310 12910 272324
rect 13080 272310 13150 272324
rect 13450 272200 13520 272220
rect 13690 272200 13760 272220
rect 13450 272166 13520 272200
rect 13690 272166 13760 272200
rect 13450 272150 13520 272166
rect 13690 272150 13760 272166
rect 12840 272042 12910 272060
rect 13080 272042 13150 272060
rect 12840 272008 12910 272042
rect 13080 272008 13150 272042
rect 12840 271990 12910 272008
rect 13080 271990 13150 272008
rect 13450 271884 13520 271900
rect 13690 271884 13760 271900
rect 13450 271850 13520 271884
rect 13690 271850 13760 271884
rect 13450 271830 13520 271850
rect 13690 271830 13760 271850
rect 12840 271726 12910 271740
rect 13080 271726 13150 271740
rect 12840 271692 12910 271726
rect 13080 271692 13150 271726
rect 12840 271670 12910 271692
rect 13080 271670 13150 271692
rect 13450 271568 13520 271580
rect 13690 271568 13760 271580
rect 13450 271534 13520 271568
rect 13690 271534 13760 271568
rect 13450 271510 13520 271534
rect 13690 271510 13760 271534
rect 12840 271410 12910 271430
rect 13080 271410 13150 271430
rect 12840 271376 12910 271410
rect 13080 271376 13150 271410
rect 12840 271360 12910 271376
rect 13080 271360 13150 271376
rect 13450 271252 13520 271270
rect 13690 271252 13760 271270
rect 13450 271218 13520 271252
rect 13690 271218 13760 271252
rect 13450 271200 13520 271218
rect 13690 271200 13760 271218
rect 12840 271094 12910 271110
rect 13080 271094 13150 271110
rect 12840 271060 12910 271094
rect 13080 271060 13150 271094
rect 12840 271040 12910 271060
rect 13080 271040 13150 271060
rect 15150 274332 15220 274350
rect 15360 274332 15430 274350
rect 15150 274298 15220 274332
rect 15360 274298 15430 274332
rect 15150 274280 15220 274298
rect 15360 274280 15430 274298
rect 16690 274332 16760 274350
rect 16900 274332 16970 274350
rect 16690 274298 16760 274332
rect 16900 274298 16970 274332
rect 16690 274280 16760 274298
rect 16900 274280 16970 274298
rect 14510 274174 14580 274190
rect 14720 274174 14790 274190
rect 14510 274140 14580 274174
rect 14720 274140 14790 274174
rect 14510 274120 14580 274140
rect 14720 274120 14790 274140
rect 16060 274174 16130 274190
rect 16270 274174 16340 274190
rect 16060 274140 16130 274174
rect 16270 274140 16340 274174
rect 15150 274016 15220 274040
rect 15360 274016 15430 274040
rect 16060 274120 16130 274140
rect 16270 274120 16340 274140
rect 15150 273982 15220 274016
rect 15360 273982 15430 274016
rect 15150 273970 15220 273982
rect 15360 273970 15430 273982
rect 14510 273858 14580 273880
rect 14720 273858 14790 273880
rect 14510 273824 14580 273858
rect 14720 273824 14790 273858
rect 14510 273810 14580 273824
rect 14720 273810 14790 273824
rect 15150 273700 15220 273720
rect 15360 273700 15430 273720
rect 15150 273666 15220 273700
rect 15360 273666 15430 273700
rect 15150 273650 15220 273666
rect 15360 273650 15430 273666
rect 16690 274016 16760 274030
rect 16900 274016 16970 274030
rect 16690 273982 16760 274016
rect 16900 273982 16970 274016
rect 16690 273960 16760 273982
rect 16900 273960 16970 273982
rect 16060 273858 16130 273880
rect 16270 273858 16340 273880
rect 16060 273824 16130 273858
rect 16270 273824 16340 273858
rect 16060 273810 16130 273824
rect 16270 273810 16340 273824
rect 16690 273700 16760 273720
rect 16900 273700 16970 273720
rect 14000 273060 14270 273330
rect 14000 272010 14270 272280
rect 14510 273542 14580 273560
rect 14720 273542 14790 273560
rect 14510 273508 14580 273542
rect 14720 273508 14790 273542
rect 14510 273490 14580 273508
rect 14720 273490 14790 273508
rect 15150 273384 15220 273400
rect 15360 273384 15430 273400
rect 15150 273350 15220 273384
rect 15360 273350 15430 273384
rect 15150 273330 15220 273350
rect 15360 273330 15430 273350
rect 14510 273226 14580 273250
rect 14720 273226 14790 273250
rect 16690 273666 16760 273700
rect 16900 273666 16970 273700
rect 16690 273650 16760 273666
rect 16900 273650 16970 273666
rect 15610 273280 15620 273540
rect 15620 273280 15860 273540
rect 15860 273280 15870 273540
rect 14510 273192 14580 273226
rect 14720 273192 14790 273226
rect 14510 273180 14580 273192
rect 14720 273180 14790 273192
rect 15150 273068 15220 273090
rect 15360 273068 15430 273090
rect 16060 273542 16130 273560
rect 16270 273542 16340 273560
rect 16060 273508 16130 273542
rect 16270 273508 16340 273542
rect 16060 273490 16130 273508
rect 16270 273490 16340 273508
rect 20510 274910 20620 275020
rect 21620 274910 21730 275020
rect 22030 274910 22140 275020
rect 23140 274910 23250 275020
rect 20510 274660 20620 274770
rect 21620 274660 21730 274770
rect 22030 274660 22140 274770
rect 23140 274660 23250 274770
rect 20660 274220 20730 274240
rect 20840 274220 20910 274240
rect 20660 274186 20730 274220
rect 20840 274186 20910 274220
rect 20660 274170 20730 274186
rect 20840 274170 20910 274186
rect 21330 273962 21400 273980
rect 21510 273962 21580 273980
rect 21330 273928 21400 273962
rect 21510 273928 21580 273962
rect 21330 273910 21400 273928
rect 21510 273910 21580 273928
rect 20660 273704 20730 273720
rect 20840 273704 20910 273720
rect 20660 273670 20730 273704
rect 20840 273670 20910 273704
rect 16690 273384 16760 273400
rect 16900 273384 16970 273400
rect 16690 273350 16760 273384
rect 16900 273350 16970 273384
rect 16690 273330 16760 273350
rect 16900 273330 16970 273350
rect 16060 273226 16130 273240
rect 16270 273226 16340 273240
rect 16060 273192 16130 273226
rect 16270 273192 16340 273226
rect 15150 273034 15220 273068
rect 15360 273034 15430 273068
rect 15150 273020 15220 273034
rect 15360 273020 15430 273034
rect 14510 272910 14580 272930
rect 14720 272910 14790 272930
rect 14510 272876 14580 272910
rect 14720 272876 14790 272910
rect 14510 272860 14580 272876
rect 14720 272860 14790 272876
rect 16060 273170 16130 273192
rect 16270 273170 16340 273192
rect 16690 273068 16760 273090
rect 16900 273068 16970 273090
rect 16690 273034 16760 273068
rect 16900 273034 16970 273068
rect 16690 273020 16760 273034
rect 16900 273020 16970 273034
rect 16060 272910 16130 272930
rect 16270 272910 16340 272930
rect 18180 273221 18250 273240
rect 18470 273221 18540 273240
rect 18180 273187 18250 273221
rect 18470 273187 18540 273221
rect 18180 273170 18250 273187
rect 18470 273170 18540 273187
rect 17620 273063 17690 273080
rect 17910 273063 17980 273080
rect 17620 273029 17690 273063
rect 17910 273029 17980 273063
rect 16060 272876 16130 272910
rect 16270 272876 16340 272910
rect 16060 272860 16130 272876
rect 16270 272860 16340 272876
rect 15150 272752 15220 272770
rect 15360 272752 15430 272770
rect 15150 272718 15220 272752
rect 15360 272718 15430 272752
rect 15150 272700 15220 272718
rect 15360 272700 15430 272718
rect 16690 272752 16760 272770
rect 16900 272752 16970 272770
rect 16690 272718 16760 272752
rect 16900 272718 16970 272752
rect 16690 272700 16760 272718
rect 16900 272700 16970 272718
rect 14510 272594 14580 272610
rect 14720 272594 14790 272610
rect 14510 272560 14580 272594
rect 14720 272560 14790 272594
rect 14510 272540 14580 272560
rect 14720 272540 14790 272560
rect 16060 272594 16130 272610
rect 16270 272594 16340 272610
rect 16060 272560 16130 272594
rect 16270 272560 16340 272594
rect 15150 272436 15220 272460
rect 15360 272436 15430 272460
rect 15150 272402 15220 272436
rect 15360 272402 15430 272436
rect 15150 272390 15220 272402
rect 15360 272390 15430 272402
rect 14510 272278 14580 272300
rect 14720 272278 14790 272300
rect 14510 272244 14580 272278
rect 14720 272244 14790 272278
rect 14510 272230 14580 272244
rect 14720 272230 14790 272244
rect 16060 272540 16130 272560
rect 16270 272540 16340 272560
rect 16690 272436 16760 272450
rect 16900 272436 16970 272450
rect 16690 272402 16760 272436
rect 16900 272402 16970 272436
rect 16690 272380 16760 272402
rect 16900 272380 16970 272402
rect 15150 272120 15220 272140
rect 15360 272120 15430 272140
rect 15150 272086 15220 272120
rect 15360 272086 15430 272120
rect 15150 272070 15220 272086
rect 15360 272070 15430 272086
rect 14510 271962 14580 271980
rect 14720 271962 14790 271980
rect 14510 271928 14580 271962
rect 14720 271928 14790 271962
rect 14510 271910 14580 271928
rect 14720 271910 14790 271928
rect 15150 271804 15220 271820
rect 15360 271804 15430 271820
rect 15150 271770 15220 271804
rect 15360 271770 15430 271804
rect 15150 271750 15220 271770
rect 15360 271750 15430 271770
rect 16060 272278 16130 272300
rect 16270 272278 16340 272300
rect 17620 273010 17690 273029
rect 17910 273010 17980 273029
rect 19700 273221 19770 273240
rect 19990 273221 20060 273240
rect 19700 273187 19770 273221
rect 19990 273187 20060 273221
rect 19700 273170 19770 273187
rect 19990 273170 20060 273187
rect 19140 273063 19210 273080
rect 19430 273063 19500 273080
rect 19140 273029 19210 273063
rect 19430 273029 19500 273063
rect 18180 272905 18250 272920
rect 18470 272905 18540 272920
rect 18180 272871 18250 272905
rect 18470 272871 18540 272905
rect 18180 272850 18250 272871
rect 18470 272850 18540 272871
rect 17620 272747 17690 272760
rect 17910 272747 17980 272760
rect 17620 272713 17690 272747
rect 17910 272713 17980 272747
rect 17620 272690 17690 272713
rect 17910 272690 17980 272713
rect 18180 272589 18250 272600
rect 18470 272589 18540 272600
rect 18180 272555 18250 272589
rect 18470 272555 18540 272589
rect 18180 272530 18250 272555
rect 18470 272530 18540 272555
rect 17620 272431 17690 272450
rect 17910 272431 17980 272450
rect 19140 273010 19210 273029
rect 19430 273010 19500 273029
rect 19700 272905 19770 272920
rect 19990 272905 20060 272920
rect 19700 272871 19770 272905
rect 19990 272871 20060 272905
rect 18710 272520 18719 272780
rect 18719 272520 18753 272780
rect 18753 272520 18925 272780
rect 18925 272520 18959 272780
rect 18959 272520 18970 272780
rect 17620 272397 17690 272431
rect 17910 272397 17980 272431
rect 17620 272380 17690 272397
rect 17910 272380 17980 272397
rect 16060 272244 16130 272278
rect 16270 272244 16340 272278
rect 16060 272230 16130 272244
rect 16270 272230 16340 272244
rect 16690 272120 16760 272140
rect 16900 272120 16970 272140
rect 16690 272086 16760 272120
rect 16900 272086 16970 272120
rect 16690 272070 16760 272086
rect 16900 272070 16970 272086
rect 15610 271780 15620 272040
rect 15620 271780 15860 272040
rect 15860 271780 15870 272040
rect 14510 271646 14580 271660
rect 14720 271646 14790 271660
rect 14510 271612 14580 271646
rect 14720 271612 14790 271646
rect 14510 271590 14580 271612
rect 14720 271590 14790 271612
rect 16060 271962 16130 271980
rect 16270 271962 16340 271980
rect 16060 271928 16130 271962
rect 16270 271928 16340 271962
rect 16060 271910 16130 271928
rect 16270 271910 16340 271928
rect 19700 272850 19770 272871
rect 19990 272850 20060 272871
rect 19140 272747 19210 272760
rect 19430 272747 19500 272760
rect 19140 272713 19210 272747
rect 19430 272713 19500 272747
rect 19140 272690 19210 272713
rect 19430 272690 19500 272713
rect 19700 272589 19770 272600
rect 19990 272589 20060 272600
rect 19700 272555 19770 272589
rect 19990 272555 20060 272589
rect 19700 272530 19770 272555
rect 19990 272530 20060 272555
rect 19140 272431 19210 272450
rect 19430 272431 19500 272450
rect 20660 273650 20730 273670
rect 20840 273650 20910 273670
rect 22180 274476 22250 274490
rect 22360 274476 22430 274490
rect 22180 274442 22250 274476
rect 22360 274442 22430 274476
rect 22180 274420 22250 274442
rect 22360 274420 22430 274442
rect 22850 274218 22920 274230
rect 23030 274218 23100 274230
rect 22850 274184 22920 274218
rect 23030 274184 23100 274218
rect 22850 274160 22920 274184
rect 23030 274160 23100 274184
rect 22180 273960 22250 273980
rect 22360 273960 22430 273980
rect 22180 273926 22250 273960
rect 22360 273926 22430 273960
rect 22180 273910 22250 273926
rect 22360 273910 22430 273926
rect 22850 273702 22920 273720
rect 23030 273702 23100 273720
rect 22850 273668 22920 273702
rect 23030 273668 23100 273702
rect 22850 273650 22920 273668
rect 23030 273650 23100 273668
rect 21330 273446 21400 273460
rect 21510 273446 21580 273460
rect 21330 273412 21400 273446
rect 21510 273412 21580 273446
rect 21330 273390 21400 273412
rect 21510 273390 21580 273412
rect 20660 273188 20730 273200
rect 20840 273188 20910 273200
rect 20660 273154 20730 273188
rect 20840 273154 20910 273188
rect 20660 273130 20730 273154
rect 20840 273130 20910 273154
rect 21330 272930 21400 272950
rect 21510 272930 21580 272950
rect 21330 272896 21400 272930
rect 21510 272896 21580 272930
rect 21330 272880 21400 272896
rect 21510 272880 21580 272896
rect 20230 272520 20239 272780
rect 20239 272520 20273 272780
rect 20273 272520 20446 272780
rect 20446 272520 20480 272780
rect 20480 272520 20490 272780
rect 19140 272397 19210 272431
rect 19430 272397 19500 272431
rect 19140 272380 19210 272397
rect 19430 272380 19500 272397
rect 18180 272273 18250 272290
rect 18470 272273 18540 272290
rect 18180 272239 18250 272273
rect 18470 272239 18540 272273
rect 18180 272220 18250 272239
rect 18470 272220 18540 272239
rect 17620 272115 17690 272130
rect 17910 272115 17980 272130
rect 17620 272081 17690 272115
rect 17910 272081 17980 272115
rect 17620 272060 17690 272081
rect 17910 272060 17980 272081
rect 19700 272273 19770 272290
rect 19990 272273 20060 272290
rect 19700 272239 19770 272273
rect 19990 272239 20060 272273
rect 19700 272220 19770 272239
rect 19990 272220 20060 272239
rect 19140 272115 19210 272130
rect 19430 272115 19500 272130
rect 19140 272081 19210 272115
rect 19430 272081 19500 272115
rect 19140 272060 19210 272081
rect 19430 272060 19500 272081
rect 16690 271804 16760 271820
rect 16900 271804 16970 271820
rect 16690 271770 16760 271804
rect 16900 271770 16970 271804
rect 16690 271750 16760 271770
rect 16900 271750 16970 271770
rect 15150 271488 15220 271510
rect 15360 271488 15430 271510
rect 15150 271454 15220 271488
rect 15360 271454 15430 271488
rect 15150 271440 15220 271454
rect 15360 271440 15430 271454
rect 14510 271330 14580 271350
rect 14720 271330 14790 271350
rect 14510 271296 14580 271330
rect 14720 271296 14790 271330
rect 14510 271280 14580 271296
rect 14720 271280 14790 271296
rect 16060 271646 16130 271660
rect 16270 271646 16340 271660
rect 16060 271612 16130 271646
rect 16270 271612 16340 271646
rect 16060 271590 16130 271612
rect 16270 271590 16340 271612
rect 16690 271488 16760 271510
rect 16900 271488 16970 271510
rect 16690 271454 16760 271488
rect 16900 271454 16970 271488
rect 16690 271440 16760 271454
rect 16900 271440 16970 271454
rect 16060 271330 16130 271350
rect 16270 271330 16340 271350
rect 16060 271296 16130 271330
rect 16270 271296 16340 271330
rect 16060 271280 16130 271296
rect 16270 271280 16340 271296
rect 15150 271172 15220 271190
rect 15360 271172 15430 271190
rect 15150 271138 15220 271172
rect 15360 271138 15430 271172
rect 15150 271120 15220 271138
rect 15360 271120 15430 271138
rect 16690 271172 16760 271190
rect 16900 271172 16970 271190
rect 16690 271138 16760 271172
rect 16900 271138 16970 271172
rect 16690 271120 16760 271138
rect 16900 271120 16970 271138
rect 13450 270936 13520 270950
rect 13690 270936 13760 270950
rect 13450 270902 13520 270936
rect 13690 270902 13760 270936
rect 13450 270880 13520 270902
rect 13690 270880 13760 270902
rect 14510 271014 14580 271030
rect 14720 271014 14790 271030
rect 14510 270980 14580 271014
rect 14720 270980 14790 271014
rect 14510 270960 14580 270980
rect 14720 270960 14790 270980
rect 16060 271014 16130 271030
rect 16270 271014 16340 271030
rect 16060 270980 16130 271014
rect 16270 270980 16340 271014
rect 16060 270960 16130 270980
rect 16270 270960 16340 270980
rect 12840 270778 12910 270790
rect 13080 270778 13150 270790
rect 12840 270744 12910 270778
rect 13080 270744 13150 270778
rect 12840 270720 12910 270744
rect 13080 270720 13150 270744
rect 13450 270620 13520 270640
rect 13690 270620 13760 270640
rect 13860 270648 13882 270660
rect 13882 270648 13940 270660
rect 13450 270586 13520 270620
rect 13690 270586 13760 270620
rect 13450 270570 13520 270586
rect 13690 270570 13760 270586
rect 13860 270580 13940 270648
rect 12840 270462 12910 270480
rect 13080 270462 13150 270480
rect 12840 270428 12910 270462
rect 13080 270428 13150 270462
rect 12840 270410 12910 270428
rect 13080 270410 13150 270428
rect 13450 270304 13520 270320
rect 13690 270304 13760 270320
rect 13450 270270 13520 270304
rect 13690 270270 13760 270304
rect 13450 270250 13520 270270
rect 13690 270250 13760 270270
rect 20660 272672 20730 272690
rect 20840 272672 20910 272690
rect 20660 272638 20730 272672
rect 20840 272638 20910 272672
rect 20660 272620 20730 272638
rect 20840 272620 20910 272638
rect 22180 273444 22250 273460
rect 22360 273444 22430 273460
rect 22180 273410 22250 273444
rect 22360 273410 22430 273444
rect 22180 273390 22250 273410
rect 22360 273390 22430 273410
rect 22850 273186 22920 273200
rect 23030 273186 23100 273200
rect 22850 273152 22920 273186
rect 23030 273152 23100 273186
rect 22850 273130 22920 273152
rect 23030 273130 23100 273152
rect 22180 272928 22250 272940
rect 22360 272928 22430 272940
rect 22180 272894 22250 272928
rect 22360 272894 22430 272928
rect 21750 272530 21760 272780
rect 21760 272530 21794 272780
rect 21794 272530 21966 272780
rect 21966 272530 22000 272780
rect 21330 272414 21400 272430
rect 21510 272414 21580 272430
rect 21330 272380 21400 272414
rect 21510 272380 21580 272414
rect 21330 272360 21400 272380
rect 21510 272360 21580 272380
rect 20660 272156 20730 272170
rect 20840 272156 20910 272170
rect 20660 272122 20730 272156
rect 20840 272122 20910 272156
rect 20660 272100 20730 272122
rect 20840 272100 20910 272122
rect 21330 271898 21400 271910
rect 21510 271898 21580 271910
rect 21330 271864 21400 271898
rect 21510 271864 21580 271898
rect 21330 271840 21400 271864
rect 21510 271840 21580 271864
rect 20660 271640 20730 271660
rect 20840 271640 20910 271660
rect 22180 272870 22250 272894
rect 22360 272870 22430 272894
rect 22850 272670 22920 272690
rect 23030 272670 23100 272690
rect 22850 272636 22920 272670
rect 23030 272636 23100 272670
rect 22850 272620 22920 272636
rect 23030 272620 23100 272636
rect 22180 272412 22250 272430
rect 22360 272412 22430 272430
rect 22180 272378 22250 272412
rect 22360 272378 22430 272412
rect 22180 272360 22250 272378
rect 22360 272360 22430 272378
rect 22850 272154 22920 272170
rect 23030 272154 23100 272170
rect 22850 272120 22920 272154
rect 23030 272120 23100 272154
rect 22850 272100 22920 272120
rect 23030 272100 23100 272120
rect 22180 271896 22250 271910
rect 22360 271896 22430 271910
rect 22180 271862 22250 271896
rect 22360 271862 22430 271896
rect 20660 271606 20730 271640
rect 20840 271606 20910 271640
rect 20660 271590 20730 271606
rect 20840 271590 20910 271606
rect 21330 271382 21400 271400
rect 21510 271382 21580 271400
rect 21330 271348 21400 271382
rect 21510 271348 21580 271382
rect 21330 271330 21400 271348
rect 21510 271330 21580 271348
rect 20660 271124 20730 271140
rect 20840 271124 20910 271140
rect 20660 271090 20730 271124
rect 20840 271090 20910 271124
rect 20660 271070 20730 271090
rect 20840 271070 20910 271090
rect 22180 271840 22250 271862
rect 22360 271840 22430 271862
rect 24400 273442 24480 273470
rect 24400 273408 24480 273442
rect 24400 273390 24480 273408
rect 26080 273590 26160 273670
rect 26220 273590 26300 273670
rect 25860 273442 25940 273470
rect 25860 273408 25940 273442
rect 24880 273184 24960 273210
rect 25230 273310 25262 273380
rect 25262 273310 25300 273380
rect 25860 273390 25940 273408
rect 26730 273380 26830 273460
rect 25560 273310 25600 273380
rect 25600 273310 25630 273380
rect 24880 273150 24960 273184
rect 24880 273130 24960 273150
rect 24400 272926 24480 272950
rect 24400 272892 24480 272926
rect 23280 272530 23314 272780
rect 23314 272530 23530 272780
rect 24400 272870 24480 272892
rect 24880 272668 24960 272690
rect 26730 273360 26762 273380
rect 26762 273360 26830 273380
rect 29310 273427 29370 273440
rect 29310 273393 29370 273427
rect 29310 273380 29370 273393
rect 25860 272926 25940 272950
rect 28170 273130 28250 273210
rect 28370 273166 28460 273190
rect 28370 273132 28460 273166
rect 25860 272892 25940 272926
rect 24880 272634 24960 272668
rect 24880 272610 24960 272634
rect 25230 272620 25300 272690
rect 25860 272870 25940 272892
rect 27470 272930 27590 273010
rect 28370 273100 28460 273132
rect 27470 272890 27590 272930
rect 29720 273169 29780 273180
rect 29720 273135 29780 273169
rect 29720 273120 29780 273135
rect 28580 272990 28612 273050
rect 28612 272990 28640 273050
rect 28940 272990 28968 273050
rect 28968 272990 29000 273050
rect 25560 272620 25630 272690
rect 24400 272410 24480 272430
rect 24400 272376 24480 272410
rect 24400 272350 24480 272376
rect 24880 272152 24960 272170
rect 24880 272118 24960 272152
rect 24880 272090 24960 272118
rect 22850 271638 22920 271650
rect 23030 271638 23100 271650
rect 22850 271604 22920 271638
rect 23030 271604 23100 271638
rect 22850 271580 22920 271604
rect 23030 271580 23100 271604
rect 24400 271894 24480 271920
rect 26730 272606 26800 272670
rect 25860 272410 25940 272430
rect 26730 272600 26762 272606
rect 26762 272600 26800 272606
rect 27170 272600 27240 272670
rect 27640 272652 27710 272670
rect 27640 272618 27710 272652
rect 27640 272600 27710 272618
rect 28170 272600 28240 272670
rect 28370 272650 28460 272680
rect 29310 272911 29370 272920
rect 29310 272877 29370 272911
rect 29310 272860 29370 272877
rect 28370 272616 28460 272650
rect 25860 272376 25940 272410
rect 25860 272350 25940 272376
rect 28370 272590 28460 272616
rect 28750 272580 28840 272670
rect 30490 273120 30550 273180
rect 30610 273120 30670 273180
rect 30730 273120 30790 273180
rect 29720 272653 29780 272670
rect 29720 272619 29780 272653
rect 29720 272610 29780 272619
rect 27480 272380 27600 272390
rect 27480 272340 27600 272380
rect 27480 272270 27600 272340
rect 25230 271922 25262 271990
rect 25262 271922 25300 271990
rect 25230 271920 25300 271922
rect 25560 271922 25600 271990
rect 25600 271922 25630 271990
rect 25560 271920 25630 271922
rect 24400 271860 24480 271894
rect 24400 271840 24480 271860
rect 25860 271894 25940 271920
rect 28170 272162 28218 272170
rect 28218 272162 28250 272170
rect 28170 272090 28250 272162
rect 28370 272134 28460 272160
rect 30190 272580 30220 272670
rect 30220 272580 30280 272670
rect 29310 272395 29370 272410
rect 29310 272361 29370 272395
rect 29310 272350 29370 272361
rect 28580 272220 28612 272280
rect 28612 272220 28640 272280
rect 28940 272220 28968 272280
rect 28968 272220 29000 272280
rect 28370 272100 28460 272134
rect 28370 272070 28460 272100
rect 29720 272137 29780 272150
rect 29720 272103 29780 272137
rect 29720 272090 29780 272103
rect 25860 271860 25940 271894
rect 25860 271840 25940 271860
rect 26730 271810 26830 271910
rect 29310 271879 29370 271890
rect 29310 271845 29370 271879
rect 29310 271830 29370 271845
rect 30490 272090 30550 272150
rect 30610 272090 30670 272150
rect 30730 272090 30790 272150
rect 26080 271630 26160 271710
rect 26220 271630 26300 271710
rect 22180 271380 22250 271400
rect 22360 271380 22430 271400
rect 22180 271346 22250 271380
rect 22360 271346 22430 271380
rect 22180 271330 22250 271346
rect 22360 271330 22430 271346
rect 22850 271122 22920 271140
rect 23030 271122 23100 271140
rect 22850 271088 22920 271122
rect 23030 271088 23100 271122
rect 22850 271070 22920 271088
rect 23030 271070 23100 271088
rect 22180 270864 22250 270880
rect 22360 270864 22430 270880
rect 22180 270830 22250 270864
rect 22360 270830 22430 270864
rect 22180 270810 22250 270830
rect 22360 270810 22430 270830
rect 20510 270510 20620 270620
rect 21620 270510 21730 270620
rect 22030 270510 22140 270620
rect 23140 270510 23250 270620
rect 20510 270260 20620 270370
rect 21620 270260 21730 270370
rect 22030 270260 22140 270370
rect 23140 270260 23250 270370
rect 12840 270146 12910 270160
rect 13080 270146 13150 270160
rect 12840 270112 12910 270146
rect 13080 270112 13150 270146
rect 12840 270090 12910 270112
rect 13080 270090 13150 270112
rect 13450 269988 13520 270000
rect 13690 269988 13760 270000
rect 13450 269954 13520 269988
rect 13690 269954 13760 269988
rect 13450 269930 13520 269954
rect 13690 269930 13760 269954
rect 12840 269830 12910 269850
rect 13080 269830 13150 269850
rect 19300 270000 19400 270100
rect 19500 270000 19700 270100
rect 19800 270000 19900 270100
rect 12840 269796 12910 269830
rect 13080 269796 13150 269830
rect 12840 269780 12910 269796
rect 13080 269780 13150 269796
rect 13450 269672 13520 269690
rect 13690 269672 13760 269690
rect 13450 269638 13520 269672
rect 13690 269638 13760 269672
rect 13450 269620 13520 269638
rect 13690 269620 13760 269638
rect 12840 269514 12910 269530
rect 13080 269514 13150 269530
rect 12840 269480 12910 269514
rect 13080 269480 13150 269514
rect 12840 269460 12910 269480
rect 13080 269460 13150 269480
rect 31020 269200 31260 269440
rect 32740 269200 32980 269440
rect 34460 269200 34700 269440
rect 35940 269200 36180 269440
rect 37660 269200 37900 269440
rect 39260 269200 39500 269440
rect 40980 269200 41220 269440
rect 42580 269200 42820 269440
rect 44300 269200 44540 269440
rect 537364 274938 537484 275058
rect 543734 274938 543854 275058
rect 537364 271938 537484 272058
rect 543734 271938 543854 272058
rect 44780 269200 45020 269440
rect 537364 268938 537484 269058
rect 543734 268938 543854 269058
rect 44700 268300 45000 268600
rect 44700 267800 45000 268100
rect 14540 267120 14640 267300
rect 44700 267300 45000 267600
rect 537744 267356 537777 267728
rect 537777 267356 538891 267728
rect 538891 267356 538914 267728
rect 537744 267318 538914 267356
rect 539254 267356 539297 267728
rect 539297 267356 540411 267728
rect 540411 267356 540424 267728
rect 539254 267318 540424 267356
rect 540774 267362 540807 267728
rect 540807 267362 541921 267728
rect 541921 267362 541944 267728
rect 540774 267318 541944 267362
rect 542294 267362 542317 267738
rect 542317 267362 543431 267738
rect 543431 267362 543464 267738
rect 542294 267328 543464 267362
rect 14540 266700 14640 266880
rect 44700 266800 45000 267100
rect 44700 266300 45000 266600
rect 44700 265800 45000 266100
rect 13080 264930 13150 265000
rect 13190 264820 13260 264890
rect 44700 265300 45000 265600
rect 44700 264800 45000 265100
rect 44700 264300 45000 264600
rect 44700 263800 45000 264100
rect 44700 263300 45000 263600
rect 44700 262800 45000 263100
rect 44700 262300 45000 262600
rect 44700 261800 45000 262100
rect 44700 261300 45000 261600
rect 44700 260800 45000 261100
rect 14980 252460 15100 252580
rect 15160 252460 15280 252580
rect 15340 252460 15460 252580
rect 15520 252460 15640 252580
rect 15700 252460 15820 252580
rect 9680 252364 9740 252380
rect 9845 252364 9905 252380
rect 10045 252364 10105 252380
rect 10235 252364 10295 252380
rect 10415 252364 10475 252380
rect 10615 252364 10675 252380
rect 10805 252364 10865 252380
rect 10965 252364 11025 252380
rect 11155 252364 11215 252380
rect 11330 252364 11390 252380
rect 11470 252364 11530 252380
rect 9680 252330 9740 252364
rect 9845 252330 9905 252364
rect 10045 252330 10105 252364
rect 10235 252330 10295 252364
rect 10415 252330 10475 252364
rect 10615 252330 10675 252364
rect 10805 252330 10865 252364
rect 10965 252330 11025 252364
rect 11155 252330 11215 252364
rect 11330 252330 11390 252364
rect 11470 252330 11530 252364
rect 5820 252315 5940 252320
rect 5820 252281 5918 252315
rect 5918 252281 5940 252315
rect 9680 252320 9740 252330
rect 9845 252320 9905 252330
rect 10045 252320 10105 252330
rect 10235 252320 10295 252330
rect 10415 252320 10475 252330
rect 10615 252320 10675 252330
rect 10805 252320 10865 252330
rect 10965 252320 11025 252330
rect 11155 252320 11215 252330
rect 11330 252320 11390 252330
rect 11470 252320 11530 252330
rect 5820 252200 5940 252281
rect 9680 252168 9740 252180
rect 9845 252168 9905 252180
rect 10045 252168 10105 252180
rect 10235 252168 10295 252180
rect 10415 252168 10475 252180
rect 10615 252168 10675 252180
rect 10805 252168 10865 252180
rect 10965 252168 11025 252180
rect 11155 252168 11215 252180
rect 11330 252168 11390 252180
rect 11470 252168 11530 252180
rect 9680 252134 9740 252168
rect 9845 252134 9905 252168
rect 10045 252134 10105 252168
rect 10235 252134 10295 252168
rect 10415 252134 10475 252168
rect 10615 252134 10675 252168
rect 10805 252134 10865 252168
rect 10965 252134 11025 252168
rect 11155 252134 11215 252168
rect 11330 252134 11390 252168
rect 11470 252134 11530 252168
rect 5820 252119 5940 252120
rect 5820 252085 5918 252119
rect 5918 252085 5940 252119
rect 9680 252120 9740 252134
rect 9845 252120 9905 252134
rect 10045 252120 10105 252134
rect 10235 252120 10295 252134
rect 10415 252120 10475 252134
rect 10615 252120 10675 252134
rect 10805 252120 10865 252134
rect 10965 252120 11025 252134
rect 11155 252120 11215 252134
rect 11330 252120 11390 252134
rect 11470 252120 11530 252134
rect 5820 252000 5940 252085
rect 9680 251972 9740 251980
rect 9845 251972 9905 251980
rect 10045 251972 10105 251980
rect 10235 251972 10295 251980
rect 10415 251972 10475 251980
rect 10615 251972 10675 251980
rect 10805 251972 10865 251980
rect 10965 251972 11025 251980
rect 11155 251972 11215 251980
rect 11330 251972 11390 251980
rect 11470 251972 11530 251980
rect 9680 251938 9740 251972
rect 9845 251938 9905 251972
rect 10045 251938 10105 251972
rect 10235 251938 10295 251972
rect 10415 251938 10475 251972
rect 10615 251938 10675 251972
rect 10805 251938 10865 251972
rect 10965 251938 11025 251972
rect 11155 251938 11215 251972
rect 11330 251938 11390 251972
rect 11470 251938 11530 251972
rect 5820 251889 5918 251920
rect 5918 251889 5940 251920
rect 9680 251920 9740 251938
rect 9845 251920 9905 251938
rect 10045 251920 10105 251938
rect 10235 251920 10295 251938
rect 10415 251920 10475 251938
rect 10615 251920 10675 251938
rect 10805 251920 10865 251938
rect 10965 251920 11025 251938
rect 11155 251920 11215 251938
rect 11330 251920 11390 251938
rect 11470 251920 11530 251938
rect 5820 251800 5940 251889
rect 9680 251776 9740 251790
rect 9845 251776 9905 251790
rect 10045 251776 10105 251790
rect 10235 251776 10295 251790
rect 10415 251776 10475 251790
rect 10615 251776 10675 251790
rect 10805 251776 10865 251790
rect 10965 251776 11025 251790
rect 11155 251776 11215 251790
rect 11330 251776 11390 251790
rect 11470 251776 11530 251790
rect 9680 251742 9740 251776
rect 9845 251742 9905 251776
rect 10045 251742 10105 251776
rect 10235 251742 10295 251776
rect 10415 251742 10475 251776
rect 10615 251742 10675 251776
rect 10805 251742 10865 251776
rect 10965 251742 11025 251776
rect 11155 251742 11215 251776
rect 11330 251742 11390 251776
rect 11470 251742 11530 251776
rect 5820 251693 5918 251720
rect 5918 251693 5940 251720
rect 9680 251730 9740 251742
rect 9845 251730 9905 251742
rect 10045 251730 10105 251742
rect 10235 251730 10295 251742
rect 10415 251730 10475 251742
rect 10615 251730 10675 251742
rect 10805 251730 10865 251742
rect 10965 251730 11025 251742
rect 11155 251730 11215 251742
rect 11330 251730 11390 251742
rect 11470 251730 11530 251742
rect 5820 251600 5940 251693
rect 9680 251580 9740 251590
rect 9845 251580 9905 251590
rect 10045 251580 10105 251590
rect 10235 251580 10295 251590
rect 10415 251580 10475 251590
rect 10615 251580 10675 251590
rect 10805 251580 10865 251590
rect 10965 251580 11025 251590
rect 11155 251580 11215 251590
rect 11330 251580 11390 251590
rect 11470 251580 11530 251590
rect 9680 251546 9740 251580
rect 9845 251546 9905 251580
rect 10045 251546 10105 251580
rect 10235 251546 10295 251580
rect 10415 251546 10475 251580
rect 10615 251546 10675 251580
rect 10805 251546 10865 251580
rect 10965 251546 11025 251580
rect 11155 251546 11215 251580
rect 11330 251546 11390 251580
rect 11470 251546 11530 251580
rect 5820 251497 5918 251520
rect 5918 251497 5940 251520
rect 9680 251530 9740 251546
rect 9845 251530 9905 251546
rect 10045 251530 10105 251546
rect 10235 251530 10295 251546
rect 10415 251530 10475 251546
rect 10615 251530 10675 251546
rect 10805 251530 10865 251546
rect 10965 251530 11025 251546
rect 11155 251530 11215 251546
rect 11330 251530 11390 251546
rect 11470 251530 11530 251546
rect 5820 251400 5940 251497
rect 9680 251384 9740 251400
rect 9845 251384 9905 251390
rect 10045 251384 10105 251390
rect 10235 251384 10295 251390
rect 10415 251384 10475 251390
rect 10615 251384 10675 251390
rect 10805 251384 10865 251390
rect 10965 251384 11025 251390
rect 11155 251384 11215 251390
rect 11330 251384 11390 251390
rect 11470 251384 11530 251390
rect 9680 251350 9740 251384
rect 9845 251350 9905 251384
rect 10045 251350 10105 251384
rect 10235 251350 10295 251384
rect 10415 251350 10475 251384
rect 10615 251350 10675 251384
rect 10805 251350 10865 251384
rect 10965 251350 11025 251384
rect 11155 251350 11215 251384
rect 11330 251350 11390 251384
rect 11470 251350 11530 251384
rect 9680 251340 9740 251350
rect 9845 251330 9905 251350
rect 10045 251330 10105 251350
rect 10235 251330 10295 251350
rect 10415 251330 10475 251350
rect 10615 251330 10675 251350
rect 10805 251330 10865 251350
rect 10965 251330 11025 251350
rect 11155 251330 11215 251350
rect 11330 251330 11390 251350
rect 11470 251330 11530 251350
rect 9680 241964 9740 241980
rect 9845 241964 9905 241980
rect 10045 241964 10105 241980
rect 10235 241964 10295 241980
rect 10415 241964 10475 241980
rect 10615 241964 10675 241980
rect 10805 241964 10865 241980
rect 10965 241964 11025 241980
rect 11155 241964 11215 241980
rect 11330 241964 11390 241980
rect 11470 241964 11530 241980
rect 9680 241930 9740 241964
rect 9845 241930 9905 241964
rect 10045 241930 10105 241964
rect 10235 241930 10295 241964
rect 10415 241930 10475 241964
rect 10615 241930 10675 241964
rect 10805 241930 10865 241964
rect 10965 241930 11025 241964
rect 11155 241930 11215 241964
rect 11330 241930 11390 241964
rect 11470 241930 11530 241964
rect 9680 241920 9740 241930
rect 9845 241920 9905 241930
rect 10045 241920 10105 241930
rect 10235 241920 10295 241930
rect 10415 241920 10475 241930
rect 10615 241920 10675 241930
rect 10805 241920 10865 241930
rect 10965 241920 11025 241930
rect 11155 241920 11215 241930
rect 11330 241920 11390 241930
rect 11470 241920 11530 241930
rect 9680 241768 9740 241780
rect 9845 241768 9905 241780
rect 10045 241768 10105 241780
rect 10235 241768 10295 241780
rect 10415 241768 10475 241780
rect 10615 241768 10675 241780
rect 10805 241768 10865 241780
rect 10965 241768 11025 241780
rect 11155 241768 11215 241780
rect 11330 241768 11390 241780
rect 11470 241768 11530 241780
rect 16100 241800 16300 242000
rect 9680 241734 9740 241768
rect 9845 241734 9905 241768
rect 10045 241734 10105 241768
rect 10235 241734 10295 241768
rect 10415 241734 10475 241768
rect 10615 241734 10675 241768
rect 10805 241734 10865 241768
rect 10965 241734 11025 241768
rect 11155 241734 11215 241768
rect 11330 241734 11390 241768
rect 11470 241734 11530 241768
rect 9680 241720 9740 241734
rect 9845 241720 9905 241734
rect 10045 241720 10105 241734
rect 10235 241720 10295 241734
rect 10415 241720 10475 241734
rect 10615 241720 10675 241734
rect 10805 241720 10865 241734
rect 10965 241720 11025 241734
rect 11155 241720 11215 241734
rect 11330 241720 11390 241734
rect 11470 241720 11530 241734
rect 9680 241572 9740 241580
rect 9845 241572 9905 241580
rect 10045 241572 10105 241580
rect 10235 241572 10295 241580
rect 10415 241572 10475 241580
rect 10615 241572 10675 241580
rect 10805 241572 10865 241580
rect 10965 241572 11025 241580
rect 11155 241572 11215 241580
rect 11330 241572 11390 241580
rect 11470 241572 11530 241580
rect 9680 241538 9740 241572
rect 9845 241538 9905 241572
rect 10045 241538 10105 241572
rect 10235 241538 10295 241572
rect 10415 241538 10475 241572
rect 10615 241538 10675 241572
rect 10805 241538 10865 241572
rect 10965 241538 11025 241572
rect 11155 241538 11215 241572
rect 11330 241538 11390 241572
rect 11470 241538 11530 241572
rect 9680 241520 9740 241538
rect 9845 241520 9905 241538
rect 10045 241520 10105 241538
rect 10235 241520 10295 241538
rect 10415 241520 10475 241538
rect 10615 241520 10675 241538
rect 10805 241520 10865 241538
rect 10965 241520 11025 241538
rect 11155 241520 11215 241538
rect 11330 241520 11390 241538
rect 11470 241520 11530 241538
rect 16100 241500 16130 241700
rect 16130 241500 16164 241700
rect 16164 241500 16300 241700
rect 9680 241376 9740 241390
rect 9845 241376 9905 241390
rect 10045 241376 10105 241390
rect 10235 241376 10295 241390
rect 10415 241376 10475 241390
rect 10615 241376 10675 241390
rect 10805 241376 10865 241390
rect 10965 241376 11025 241390
rect 11155 241376 11215 241390
rect 11330 241376 11390 241390
rect 11470 241376 11530 241390
rect 9680 241342 9740 241376
rect 9845 241342 9905 241376
rect 10045 241342 10105 241376
rect 10235 241342 10295 241376
rect 10415 241342 10475 241376
rect 10615 241342 10675 241376
rect 10805 241342 10865 241376
rect 10965 241342 11025 241376
rect 11155 241342 11215 241376
rect 11330 241342 11390 241376
rect 11470 241342 11530 241376
rect 9680 241330 9740 241342
rect 9845 241330 9905 241342
rect 10045 241330 10105 241342
rect 10235 241330 10295 241342
rect 10415 241330 10475 241342
rect 10615 241330 10675 241342
rect 10805 241330 10865 241342
rect 10965 241330 11025 241342
rect 11155 241330 11215 241342
rect 11330 241330 11390 241342
rect 11470 241330 11530 241342
rect 9680 241180 9740 241190
rect 9845 241180 9905 241190
rect 10045 241180 10105 241190
rect 10235 241180 10295 241190
rect 10415 241180 10475 241190
rect 10615 241180 10675 241190
rect 10805 241180 10865 241190
rect 10965 241180 11025 241190
rect 11155 241180 11215 241190
rect 11330 241180 11390 241190
rect 11470 241180 11530 241190
rect 16100 241200 16130 241400
rect 16130 241200 16164 241400
rect 16164 241200 16300 241400
rect 9680 241146 9740 241180
rect 9845 241146 9905 241180
rect 10045 241146 10105 241180
rect 10235 241146 10295 241180
rect 10415 241146 10475 241180
rect 10615 241146 10675 241180
rect 10805 241146 10865 241180
rect 10965 241146 11025 241180
rect 11155 241146 11215 241180
rect 11330 241146 11390 241180
rect 11470 241146 11530 241180
rect 9680 241130 9740 241146
rect 9845 241130 9905 241146
rect 10045 241130 10105 241146
rect 10235 241130 10295 241146
rect 10415 241130 10475 241146
rect 10615 241130 10675 241146
rect 10805 241130 10865 241146
rect 10965 241130 11025 241146
rect 11155 241130 11215 241146
rect 11330 241130 11390 241146
rect 11470 241130 11530 241146
rect 9680 240984 9740 241000
rect 9845 240984 9905 240990
rect 10045 240984 10105 240990
rect 10235 240984 10295 240990
rect 10415 240984 10475 240990
rect 10615 240984 10675 240990
rect 10805 240984 10865 240990
rect 10965 240984 11025 240990
rect 11155 240984 11215 240990
rect 11330 240984 11390 240990
rect 11470 240984 11530 240990
rect 9680 240950 9740 240984
rect 9845 240950 9905 240984
rect 10045 240950 10105 240984
rect 10235 240950 10295 240984
rect 10415 240950 10475 240984
rect 10615 240950 10675 240984
rect 10805 240950 10865 240984
rect 10965 240950 11025 240984
rect 11155 240950 11215 240984
rect 11330 240950 11390 240984
rect 11470 240950 11530 240984
rect 9680 240940 9740 240950
rect 9845 240930 9905 240950
rect 10045 240930 10105 240950
rect 10235 240930 10295 240950
rect 10415 240930 10475 240950
rect 10615 240930 10675 240950
rect 10805 240930 10865 240950
rect 10965 240930 11025 240950
rect 11155 240930 11215 240950
rect 11330 240930 11390 240950
rect 11470 240930 11530 240950
rect 16100 240900 16300 241100
<< metal2 >>
rect 65060 702260 65240 702270
rect 23400 702180 23520 702190
rect 23400 702050 23520 702060
rect 23600 702180 23720 702190
rect 23600 702050 23720 702060
rect 23800 702180 23920 702190
rect 23800 702050 23920 702060
rect 24000 702180 24120 702190
rect 24000 702050 24120 702060
rect 24200 702180 24320 702190
rect 65060 702070 65240 702080
rect 65400 702260 65580 702270
rect 65400 702070 65580 702080
rect 65740 702260 65920 702270
rect 573280 702240 573380 702250
rect 65740 702070 65920 702080
rect 563800 702120 565120 702160
rect 573280 702130 573380 702140
rect 573420 702240 573520 702250
rect 573420 702130 573520 702140
rect 573560 702240 573660 702250
rect 573560 702130 573660 702140
rect 573700 702240 573800 702250
rect 573700 702130 573800 702140
rect 573840 702240 573940 702250
rect 573840 702130 573940 702140
rect 573980 702240 574080 702250
rect 573980 702130 574080 702140
rect 24200 702050 24320 702060
rect 563800 702020 563840 702120
rect 563940 702020 563980 702120
rect 564080 702020 564120 702120
rect 564220 702020 564260 702120
rect 564360 702020 564400 702120
rect 564500 702020 564540 702120
rect 564640 702020 564680 702120
rect 564780 702020 564820 702120
rect 564920 702020 564960 702120
rect 565060 702020 565120 702120
rect 563800 701980 565120 702020
rect 563800 701880 563840 701980
rect 563940 701880 563980 701980
rect 564080 701880 564120 701980
rect 564220 701880 564260 701980
rect 564360 701880 564400 701980
rect 564500 701880 564540 701980
rect 564640 701880 564680 701980
rect 564780 701880 564820 701980
rect 564920 701880 564960 701980
rect 565060 701880 565120 701980
rect 563800 701840 565120 701880
rect 573280 701980 573380 701990
rect 573280 701870 573380 701880
rect 573420 701980 573520 701990
rect 573420 701870 573520 701880
rect 573560 701980 573660 701990
rect 573560 701870 573660 701880
rect 573700 701980 573800 701990
rect 573700 701870 573800 701880
rect 573840 701980 573940 701990
rect 573840 701870 573940 701880
rect 573980 701980 574080 701990
rect 573980 701870 574080 701880
rect 24460 693020 24580 693030
rect 24460 692890 24580 692900
rect 64720 693000 64860 693010
rect 64720 692850 64860 692860
rect 66060 693000 66200 693010
rect 66060 692850 66200 692860
rect 75120 693000 75260 693010
rect 75120 692850 75260 692860
rect 24460 692840 24580 692850
rect 24460 692710 24580 692720
rect 64720 692800 64860 692810
rect 24460 692660 24580 692670
rect 64720 692650 64860 692660
rect 66060 692800 66200 692810
rect 66060 692650 66200 692660
rect 75120 692800 75260 692810
rect 75120 692650 75260 692660
rect 24460 692530 24580 692540
rect 24460 692480 24580 692490
rect 24460 692350 24580 692360
rect 24460 692300 24580 692310
rect 24460 692170 24580 692180
rect 12900 691900 13100 691910
rect 12900 691690 13100 691700
rect 13200 691900 13400 691910
rect 13200 691690 13400 691700
rect 13500 691900 13700 691910
rect 13500 691690 13700 691700
rect 13800 691900 14000 691910
rect 13800 691690 14000 691700
rect 566290 690900 566300 691100
rect 566500 690900 566510 691100
rect 566690 690900 566700 691100
rect 566900 690900 566910 691100
rect 567090 690900 567100 691100
rect 567300 690900 567310 691100
rect 567490 690900 567500 691100
rect 567700 690900 567710 691100
rect 567890 690900 567900 691100
rect 568100 690900 568110 691100
rect 568290 690900 568300 691100
rect 568500 690900 568510 691100
rect 568690 690900 568700 691100
rect 568900 690900 568910 691100
rect 569090 690900 569100 691100
rect 569300 690900 569310 691100
rect 569490 690900 569500 691100
rect 569700 690900 569710 691100
rect 569890 690900 569900 691100
rect 570100 690900 570110 691100
rect 570290 690900 570300 691100
rect 570500 690900 570510 691100
rect 570690 690900 570700 691100
rect 570900 690900 570910 691100
rect 571090 690900 571100 691100
rect 571300 690900 571310 691100
rect 571490 690900 571500 691100
rect 571700 690900 571710 691100
rect 566290 690500 566300 690700
rect 566500 690500 566510 690700
rect 566690 690500 566700 690700
rect 566900 690500 566910 690700
rect 567090 690500 567100 690700
rect 567300 690500 567310 690700
rect 567490 690500 567500 690700
rect 567700 690500 567710 690700
rect 567890 690500 567900 690700
rect 568100 690500 568110 690700
rect 568290 690500 568300 690700
rect 568500 690500 568510 690700
rect 568690 690500 568700 690700
rect 568900 690500 568910 690700
rect 569090 690500 569100 690700
rect 569300 690500 569310 690700
rect 569490 690500 569500 690700
rect 569700 690500 569710 690700
rect 569890 690500 569900 690700
rect 570100 690500 570110 690700
rect 570290 690500 570300 690700
rect 570500 690500 570510 690700
rect 570690 690500 570700 690700
rect 570900 690500 570910 690700
rect 571090 690500 571100 690700
rect 571300 690500 571310 690700
rect 571490 690500 571500 690700
rect 571700 690500 571710 690700
rect 47200 690300 47300 690310
rect 47200 690190 47300 690200
rect 566290 690100 566300 690300
rect 566500 690100 566510 690300
rect 566690 690100 566700 690300
rect 566900 690100 566910 690300
rect 567090 690100 567100 690300
rect 567300 690100 567310 690300
rect 567490 690100 567500 690300
rect 567700 690100 567710 690300
rect 567890 690100 567900 690300
rect 568100 690100 568110 690300
rect 568290 690100 568300 690300
rect 568500 690100 568510 690300
rect 568690 690100 568700 690300
rect 568900 690100 568910 690300
rect 569090 690100 569100 690300
rect 569300 690100 569310 690300
rect 569490 690100 569500 690300
rect 569700 690100 569710 690300
rect 569890 690100 569900 690300
rect 570100 690100 570110 690300
rect 570290 690100 570300 690300
rect 570500 690100 570510 690300
rect 570690 690100 570700 690300
rect 570900 690100 570910 690300
rect 571090 690100 571100 690300
rect 571300 690100 571310 690300
rect 571490 690100 571500 690300
rect 571700 690100 571710 690300
rect 47200 690000 47300 690010
rect 47200 689790 47300 689800
rect 566290 689700 566300 689900
rect 566500 689700 566510 689900
rect 566690 689700 566700 689900
rect 566900 689700 566910 689900
rect 567090 689700 567100 689900
rect 567300 689700 567310 689900
rect 567490 689700 567500 689900
rect 567700 689700 567710 689900
rect 567890 689700 567900 689900
rect 568100 689700 568110 689900
rect 568290 689700 568300 689900
rect 568500 689700 568510 689900
rect 568690 689700 568700 689900
rect 568900 689700 568910 689900
rect 569090 689700 569100 689900
rect 569300 689700 569310 689900
rect 569490 689700 569500 689900
rect 569700 689700 569710 689900
rect 569890 689700 569900 689900
rect 570100 689700 570110 689900
rect 570290 689700 570300 689900
rect 570500 689700 570510 689900
rect 570690 689700 570700 689900
rect 570900 689700 570910 689900
rect 571090 689700 571100 689900
rect 571300 689700 571310 689900
rect 571490 689700 571500 689900
rect 571700 689700 571710 689900
rect 47200 689600 47300 689610
rect 47200 689490 47300 689500
rect 566290 689300 566300 689500
rect 566500 689300 566510 689500
rect 566690 689300 566700 689500
rect 566900 689300 566910 689500
rect 567090 689300 567100 689500
rect 567300 689300 567310 689500
rect 567490 689300 567500 689500
rect 567700 689300 567710 689500
rect 567890 689300 567900 689500
rect 568100 689300 568110 689500
rect 568290 689300 568300 689500
rect 568500 689300 568510 689500
rect 568690 689300 568700 689500
rect 568900 689300 568910 689500
rect 569090 689300 569100 689500
rect 569300 689300 569310 689500
rect 569490 689300 569500 689500
rect 569700 689300 569710 689500
rect 569890 689300 569900 689500
rect 570100 689300 570110 689500
rect 570290 689300 570300 689500
rect 570500 689300 570510 689500
rect 570690 689300 570700 689500
rect 570900 689300 570910 689500
rect 571090 689300 571100 689500
rect 571300 689300 571310 689500
rect 571490 689300 571500 689500
rect 571700 689300 571710 689500
rect 42000 688700 42100 688710
rect 42000 688590 42100 688600
rect 42000 688500 42100 688510
rect 42000 688290 42100 688300
rect 42000 688200 42100 688210
rect 42000 688090 42100 688100
rect 42240 683120 42640 684610
rect 42240 683040 42260 683120
rect 42340 683040 42400 683120
rect 42480 683040 42540 683120
rect 42620 683040 42640 683120
rect 42240 683020 42640 683040
rect 46640 683120 47040 684610
rect 582360 684600 582440 684610
rect 582360 684510 582440 684520
rect 582540 684600 582620 684610
rect 582540 684510 582620 684520
rect 582360 684440 582440 684450
rect 582360 684350 582440 684360
rect 582540 684440 582620 684450
rect 582540 684350 582620 684360
rect 582360 684280 582440 684290
rect 582360 684190 582440 684200
rect 582540 684280 582620 684290
rect 582540 684190 582620 684200
rect 582360 684100 582440 684110
rect 582360 684010 582440 684020
rect 582540 684100 582620 684110
rect 582540 684010 582620 684020
rect 582360 683940 582440 683950
rect 582360 683850 582440 683860
rect 582540 683940 582620 683950
rect 582540 683850 582620 683860
rect 46640 683040 46660 683120
rect 46740 683040 46800 683120
rect 46880 683040 46940 683120
rect 47020 683040 47040 683120
rect 46640 683020 47040 683040
rect 561700 682200 561900 682210
rect 561700 681990 561900 682000
rect 562100 682200 562300 682210
rect 562100 681990 562300 682000
rect 562500 682200 562700 682210
rect 562500 681990 562700 682000
rect 562900 682200 563100 682210
rect 562900 681990 563100 682000
rect 563300 682200 563500 682210
rect 563300 681990 563500 682000
rect 561700 681800 561900 681810
rect 561700 681590 561900 681600
rect 562100 681800 562300 681810
rect 562100 681590 562300 681600
rect 562500 681800 562700 681810
rect 562500 681590 562700 681600
rect 562900 681800 563100 681810
rect 562900 681590 563100 681600
rect 563300 681800 563500 681810
rect 563300 681590 563500 681600
rect 561700 681400 561900 681410
rect 561700 681190 561900 681200
rect 562100 681400 562300 681410
rect 562100 681190 562300 681200
rect 562500 681400 562700 681410
rect 562500 681190 562700 681200
rect 562900 681400 563100 681410
rect 562900 681190 563100 681200
rect 563300 681400 563500 681410
rect 563300 681190 563500 681200
rect 561700 681000 561900 681010
rect 561700 680790 561900 680800
rect 562100 681000 562300 681010
rect 562100 680790 562300 680800
rect 562500 681000 562700 681010
rect 562500 680790 562700 680800
rect 562900 681000 563100 681010
rect 562900 680790 563100 680800
rect 563300 681000 563500 681010
rect 563300 680790 563500 680800
rect 561700 680600 561900 680610
rect 561700 680390 561900 680400
rect 562100 680600 562300 680610
rect 562100 680390 562300 680400
rect 562500 680600 562700 680610
rect 562500 680390 562700 680400
rect 562900 680600 563100 680610
rect 562900 680390 563100 680400
rect 563300 680600 563500 680610
rect 563300 680390 563500 680400
rect 561700 680200 561900 680210
rect 561700 679990 561900 680000
rect 562100 680200 562300 680210
rect 562100 679990 562300 680000
rect 562500 680200 562700 680210
rect 562500 679990 562700 680000
rect 562900 680200 563100 680210
rect 562900 679990 563100 680000
rect 563300 680200 563500 680210
rect 563300 679990 563500 680000
rect 561700 679800 561900 679810
rect 561700 679590 561900 679600
rect 562100 679800 562300 679810
rect 562100 679590 562300 679600
rect 562500 679800 562700 679810
rect 562500 679590 562700 679600
rect 562900 679800 563100 679810
rect 562900 679590 563100 679600
rect 563300 679800 563500 679810
rect 563300 679590 563500 679600
rect 561700 679400 561900 679410
rect 561700 679190 561900 679200
rect 562100 679400 562300 679410
rect 562100 679190 562300 679200
rect 562500 679400 562700 679410
rect 562500 679190 562700 679200
rect 562900 679400 563100 679410
rect 562900 679190 563100 679200
rect 563300 679400 563500 679410
rect 563300 679190 563500 679200
rect 561700 679000 561900 679010
rect 561700 678790 561900 678800
rect 562100 679000 562300 679010
rect 562100 678790 562300 678800
rect 562500 679000 562700 679010
rect 562500 678790 562700 678800
rect 562900 679000 563100 679010
rect 562900 678790 563100 678800
rect 563300 679000 563500 679010
rect 563300 678790 563500 678800
rect 561700 678600 561900 678610
rect 561700 678390 561900 678400
rect 562100 678600 562300 678610
rect 562100 678390 562300 678400
rect 562500 678600 562700 678610
rect 562500 678390 562700 678400
rect 562900 678600 563100 678610
rect 562900 678390 563100 678400
rect 563300 678600 563500 678610
rect 563300 678390 563500 678400
rect 571900 677300 572100 677310
rect 571900 677090 572100 677100
rect 571900 677000 572100 677010
rect 571900 676790 572100 676800
rect 571900 676700 572100 676710
rect 571900 676490 572100 676500
rect 571900 676400 572100 676410
rect 571900 676190 572100 676200
rect 32800 663300 33100 663310
rect 32800 662990 33100 663000
rect 33300 663300 33600 663310
rect 33300 662990 33600 663000
rect 33800 663300 34100 663310
rect 33800 662990 34100 663000
rect 34300 663300 34600 663310
rect 34300 662990 34600 663000
rect 34800 663300 35100 663310
rect 34800 662990 35100 663000
rect 35300 663300 35600 663310
rect 35300 662990 35600 663000
rect 35800 663300 36100 663310
rect 35800 662990 36100 663000
rect 36300 663300 36600 663310
rect 36300 662990 36600 663000
rect 36800 663300 37100 663310
rect 36800 662990 37100 663000
rect 37300 663300 37600 663310
rect 37300 662990 37600 663000
rect 37800 663300 38100 663310
rect 37800 662990 38100 663000
rect 38300 663300 38600 663310
rect 38300 662990 38600 663000
rect 38800 663300 39100 663310
rect 38800 662990 39100 663000
rect 39300 663300 39600 663310
rect 39300 662990 39600 663000
rect 39800 663300 40100 663310
rect 39800 662990 40100 663000
rect 40300 663300 40600 663310
rect 40300 662990 40600 663000
rect 294760 352660 294820 352670
rect 281080 352640 281140 352650
rect 281080 352570 281140 352580
rect 281180 352640 281240 352650
rect 294760 352590 294820 352600
rect 294860 352660 294920 352670
rect 294860 352590 294920 352600
rect 281180 352570 281240 352580
rect 294760 352560 294820 352570
rect 281080 352540 281140 352550
rect 281080 352470 281140 352480
rect 281180 352540 281240 352550
rect 294760 352490 294820 352500
rect 294860 352560 294920 352570
rect 294860 352490 294920 352500
rect 281180 352470 281240 352480
rect 281060 351080 281120 351090
rect 281060 351010 281120 351020
rect 281160 351080 281220 351090
rect 281160 351010 281220 351020
rect 281060 350980 281120 350990
rect 281060 350910 281120 350920
rect 281160 350980 281220 350990
rect 281160 350910 281220 350920
rect 294760 350920 294820 350930
rect 294760 350850 294820 350860
rect 294860 350920 294920 350930
rect 294860 350850 294920 350860
rect 294760 350820 294820 350830
rect 294760 350750 294820 350760
rect 294860 350820 294920 350830
rect 294860 350750 294920 350760
rect 281060 349380 281120 349390
rect 281060 349310 281120 349320
rect 281160 349380 281220 349390
rect 281160 349310 281220 349320
rect 281060 349280 281120 349290
rect 281060 349210 281120 349220
rect 281160 349280 281220 349290
rect 281160 349210 281220 349220
rect 294760 349220 294820 349230
rect 294760 349150 294820 349160
rect 294860 349220 294920 349230
rect 294860 349150 294920 349160
rect 294760 349120 294820 349130
rect 294760 349050 294820 349060
rect 294860 349120 294920 349130
rect 294860 349050 294920 349060
rect 281040 347680 281100 347690
rect 281040 347610 281100 347620
rect 281140 347680 281200 347690
rect 281140 347610 281200 347620
rect 281040 347580 281100 347590
rect 281040 347510 281100 347520
rect 281140 347580 281200 347590
rect 281140 347510 281200 347520
rect 294760 347520 294820 347530
rect 294760 347450 294820 347460
rect 294860 347520 294920 347530
rect 294860 347450 294920 347460
rect 294760 347420 294820 347430
rect 294760 347350 294820 347360
rect 294860 347420 294920 347430
rect 294860 347350 294920 347360
rect 281060 345980 281120 345990
rect 281060 345910 281120 345920
rect 281160 345980 281220 345990
rect 281160 345910 281220 345920
rect 281060 345880 281120 345890
rect 281060 345810 281120 345820
rect 281160 345880 281220 345890
rect 281160 345810 281220 345820
rect 294760 345820 294820 345830
rect 294760 345750 294820 345760
rect 294860 345820 294920 345830
rect 294860 345750 294920 345760
rect 294760 345720 294820 345730
rect 294760 345650 294820 345660
rect 294860 345720 294920 345730
rect 294860 345650 294920 345660
rect 281060 344260 281120 344270
rect 281060 344190 281120 344200
rect 281160 344260 281220 344270
rect 281160 344190 281220 344200
rect 294800 344200 295100 344210
rect 281060 344160 281120 344170
rect 281060 344090 281120 344100
rect 281160 344160 281220 344170
rect 281160 344090 281220 344100
rect 294800 343890 295100 343900
rect 281040 342560 281100 342570
rect 281040 342490 281100 342500
rect 281140 342560 281200 342570
rect 281140 342490 281200 342500
rect 281040 342460 281100 342470
rect 281040 342390 281100 342400
rect 281140 342460 281200 342470
rect 281140 342390 281200 342400
rect 294760 342420 294820 342430
rect 294760 342350 294820 342360
rect 294860 342420 294920 342430
rect 294860 342350 294920 342360
rect 294760 342320 294820 342330
rect 294760 342250 294820 342260
rect 294860 342320 294920 342330
rect 294860 342250 294920 342260
rect 288300 340800 288600 340810
rect 281060 340720 281120 340730
rect 281060 340650 281120 340660
rect 281160 340720 281220 340730
rect 281160 340650 281220 340660
rect 281060 340620 281120 340630
rect 281060 340550 281120 340560
rect 281160 340620 281220 340630
rect 281160 340550 281220 340560
rect 288300 340490 288600 340500
rect 569280 306240 569380 306250
rect 559800 306120 561120 306160
rect 569280 306130 569380 306140
rect 569420 306240 569520 306250
rect 569420 306130 569520 306140
rect 569560 306240 569660 306250
rect 569560 306130 569660 306140
rect 569700 306240 569800 306250
rect 569700 306130 569800 306140
rect 569840 306240 569940 306250
rect 569840 306130 569940 306140
rect 569980 306240 570080 306250
rect 569980 306130 570080 306140
rect 559800 306020 559840 306120
rect 559940 306020 559980 306120
rect 560080 306020 560120 306120
rect 560220 306020 560260 306120
rect 560360 306020 560400 306120
rect 560500 306020 560540 306120
rect 560640 306020 560680 306120
rect 560780 306020 560820 306120
rect 560920 306020 560960 306120
rect 561060 306020 561120 306120
rect 559800 305980 561120 306020
rect 559800 305880 559840 305980
rect 559940 305880 559980 305980
rect 560080 305880 560120 305980
rect 560220 305880 560260 305980
rect 560360 305880 560400 305980
rect 560500 305880 560540 305980
rect 560640 305880 560680 305980
rect 560780 305880 560820 305980
rect 560920 305880 560960 305980
rect 561060 305880 561120 305980
rect 559800 305840 561120 305880
rect 569280 305980 569380 305990
rect 569280 305870 569380 305880
rect 569420 305980 569520 305990
rect 569420 305870 569520 305880
rect 569560 305980 569660 305990
rect 569560 305870 569660 305880
rect 569700 305980 569800 305990
rect 569700 305870 569800 305880
rect 569840 305980 569940 305990
rect 569840 305870 569940 305880
rect 569980 305980 570080 305990
rect 569980 305870 570080 305880
rect 9670 304320 9680 304380
rect 9740 304320 9750 304380
rect 9835 304320 9845 304380
rect 9905 304320 9915 304380
rect 10035 304320 10045 304380
rect 10105 304320 10115 304380
rect 10225 304320 10235 304380
rect 10295 304320 10305 304380
rect 10405 304320 10415 304380
rect 10475 304320 10485 304380
rect 10605 304320 10615 304380
rect 10675 304320 10685 304380
rect 10795 304320 10805 304380
rect 10865 304320 10875 304380
rect 10955 304320 10965 304380
rect 11025 304320 11035 304380
rect 11145 304320 11155 304380
rect 11215 304320 11225 304380
rect 11320 304320 11330 304380
rect 11390 304320 11400 304380
rect 11460 304320 11470 304380
rect 11530 304320 11540 304380
rect 9670 304120 9680 304180
rect 9740 304120 9750 304180
rect 9835 304120 9845 304180
rect 9905 304120 9915 304180
rect 10035 304120 10045 304180
rect 10105 304120 10115 304180
rect 10225 304120 10235 304180
rect 10295 304120 10305 304180
rect 10405 304120 10415 304180
rect 10475 304120 10485 304180
rect 10605 304120 10615 304180
rect 10675 304120 10685 304180
rect 10795 304120 10805 304180
rect 10865 304120 10875 304180
rect 10955 304120 10965 304180
rect 11025 304120 11035 304180
rect 11145 304120 11155 304180
rect 11215 304120 11225 304180
rect 11320 304120 11330 304180
rect 11390 304120 11400 304180
rect 11460 304120 11470 304180
rect 11530 304120 11540 304180
rect 9670 303920 9680 303980
rect 9740 303920 9750 303980
rect 9835 303920 9845 303980
rect 9905 303920 9915 303980
rect 10035 303920 10045 303980
rect 10105 303920 10115 303980
rect 10225 303920 10235 303980
rect 10295 303920 10305 303980
rect 10405 303920 10415 303980
rect 10475 303920 10485 303980
rect 10605 303920 10615 303980
rect 10675 303920 10685 303980
rect 10795 303920 10805 303980
rect 10865 303920 10875 303980
rect 10955 303920 10965 303980
rect 11025 303920 11035 303980
rect 11145 303920 11155 303980
rect 11215 303920 11225 303980
rect 11320 303920 11330 303980
rect 11390 303920 11400 303980
rect 11460 303920 11470 303980
rect 11530 303920 11540 303980
rect 9670 303730 9680 303790
rect 9740 303730 9750 303790
rect 9835 303730 9845 303790
rect 9905 303730 9915 303790
rect 10035 303730 10045 303790
rect 10105 303730 10115 303790
rect 10225 303730 10235 303790
rect 10295 303730 10305 303790
rect 10405 303730 10415 303790
rect 10475 303730 10485 303790
rect 10605 303730 10615 303790
rect 10675 303730 10685 303790
rect 10795 303730 10805 303790
rect 10865 303730 10875 303790
rect 10955 303730 10965 303790
rect 11025 303730 11035 303790
rect 11145 303730 11155 303790
rect 11215 303730 11225 303790
rect 11320 303730 11330 303790
rect 11390 303730 11400 303790
rect 11460 303730 11470 303790
rect 11530 303730 11540 303790
rect 9670 303530 9680 303590
rect 9740 303530 9750 303590
rect 9835 303530 9845 303590
rect 9905 303530 9915 303590
rect 10035 303530 10045 303590
rect 10105 303530 10115 303590
rect 10225 303530 10235 303590
rect 10295 303530 10305 303590
rect 10405 303530 10415 303590
rect 10475 303530 10485 303590
rect 10605 303530 10615 303590
rect 10675 303530 10685 303590
rect 10795 303530 10805 303590
rect 10865 303530 10875 303590
rect 10955 303530 10965 303590
rect 11025 303530 11035 303590
rect 11145 303530 11155 303590
rect 11215 303530 11225 303590
rect 11320 303530 11330 303590
rect 11390 303530 11400 303590
rect 11460 303530 11470 303590
rect 11530 303530 11540 303590
rect 9670 303340 9680 303400
rect 9740 303340 9750 303400
rect 9835 303330 9845 303390
rect 9905 303330 9915 303390
rect 10035 303330 10045 303390
rect 10105 303330 10115 303390
rect 10225 303330 10235 303390
rect 10295 303330 10305 303390
rect 10405 303330 10415 303390
rect 10475 303330 10485 303390
rect 10605 303330 10615 303390
rect 10675 303330 10685 303390
rect 10795 303330 10805 303390
rect 10865 303330 10875 303390
rect 10955 303330 10965 303390
rect 11025 303330 11035 303390
rect 11145 303330 11155 303390
rect 11215 303330 11225 303390
rect 11320 303330 11330 303390
rect 11390 303330 11400 303390
rect 11460 303330 11470 303390
rect 11530 303330 11540 303390
rect 14990 303120 15000 303260
rect 15140 303120 15150 303260
rect 15190 303120 15200 303260
rect 15340 303120 15350 303260
rect 559940 302120 560000 302130
rect 559940 302050 560000 302060
rect 560130 302120 560190 302130
rect 560130 302050 560190 302060
rect 560330 302120 560390 302130
rect 560330 302050 560390 302060
rect 560520 302120 560580 302130
rect 560520 302050 560580 302060
rect 560720 302120 560780 302130
rect 560720 302050 560780 302060
rect 560920 302120 560980 302130
rect 560920 302050 560980 302060
rect 569140 302120 569200 302130
rect 569140 302050 569200 302060
rect 569330 302120 569390 302130
rect 569330 302050 569390 302060
rect 569530 302120 569590 302130
rect 569530 302050 569590 302060
rect 569720 302120 569780 302130
rect 569720 302050 569780 302060
rect 569920 302120 569980 302130
rect 569920 302050 569980 302060
rect 570120 302120 570180 302130
rect 570120 302050 570180 302060
rect 559930 301955 559990 301965
rect 559930 301885 559990 301895
rect 560130 301955 560190 301965
rect 560130 301885 560190 301895
rect 560330 301955 560390 301965
rect 560330 301885 560390 301895
rect 560520 301955 560580 301965
rect 560520 301885 560580 301895
rect 560720 301955 560780 301965
rect 560720 301885 560780 301895
rect 560920 301955 560980 301965
rect 560920 301885 560980 301895
rect 569130 301955 569190 301965
rect 569130 301885 569190 301895
rect 569330 301955 569390 301965
rect 569330 301885 569390 301895
rect 569530 301955 569590 301965
rect 569530 301885 569590 301895
rect 569720 301955 569780 301965
rect 569720 301885 569780 301895
rect 569920 301955 569980 301965
rect 569920 301885 569980 301895
rect 570120 301955 570180 301965
rect 570120 301885 570180 301895
rect 559930 301755 559990 301765
rect 559930 301685 559990 301695
rect 560130 301755 560190 301765
rect 560130 301685 560190 301695
rect 560330 301755 560390 301765
rect 560330 301685 560390 301695
rect 560520 301755 560580 301765
rect 560520 301685 560580 301695
rect 560720 301755 560780 301765
rect 560720 301685 560780 301695
rect 560920 301755 560980 301765
rect 560920 301685 560980 301695
rect 569130 301755 569190 301765
rect 569130 301685 569190 301695
rect 569330 301755 569390 301765
rect 569330 301685 569390 301695
rect 569530 301755 569590 301765
rect 569530 301685 569590 301695
rect 569720 301755 569780 301765
rect 569720 301685 569780 301695
rect 569920 301755 569980 301765
rect 569920 301685 569980 301695
rect 570120 301755 570180 301765
rect 570120 301685 570180 301695
rect 559930 301565 559990 301575
rect 559930 301495 559990 301505
rect 560130 301565 560190 301575
rect 560130 301495 560190 301505
rect 560330 301565 560390 301575
rect 560330 301495 560390 301505
rect 560520 301565 560580 301575
rect 560520 301495 560580 301505
rect 560720 301565 560780 301575
rect 560720 301495 560780 301505
rect 560920 301565 560980 301575
rect 560920 301495 560980 301505
rect 569130 301565 569190 301575
rect 569130 301495 569190 301505
rect 569330 301565 569390 301575
rect 569330 301495 569390 301505
rect 569530 301565 569590 301575
rect 569530 301495 569590 301505
rect 569720 301565 569780 301575
rect 569720 301495 569780 301505
rect 569920 301565 569980 301575
rect 569920 301495 569980 301505
rect 570120 301565 570180 301575
rect 570120 301495 570180 301505
rect 559930 301385 559990 301395
rect 559930 301315 559990 301325
rect 560130 301385 560190 301395
rect 560130 301315 560190 301325
rect 560330 301385 560390 301395
rect 560330 301315 560390 301325
rect 560520 301385 560580 301395
rect 560520 301315 560580 301325
rect 560720 301385 560780 301395
rect 560720 301315 560780 301325
rect 560920 301385 560980 301395
rect 560920 301315 560980 301325
rect 569130 301385 569190 301395
rect 569130 301315 569190 301325
rect 569330 301385 569390 301395
rect 569330 301315 569390 301325
rect 569530 301385 569590 301395
rect 569530 301315 569590 301325
rect 569720 301385 569780 301395
rect 569720 301315 569780 301325
rect 569920 301385 569980 301395
rect 569920 301315 569980 301325
rect 570120 301385 570180 301395
rect 570120 301315 570180 301325
rect 559930 301185 559990 301195
rect 559930 301115 559990 301125
rect 560130 301185 560190 301195
rect 560130 301115 560190 301125
rect 560330 301185 560390 301195
rect 560330 301115 560390 301125
rect 560520 301185 560580 301195
rect 560520 301115 560580 301125
rect 560720 301185 560780 301195
rect 560720 301115 560780 301125
rect 560920 301185 560980 301195
rect 560920 301115 560980 301125
rect 569130 301185 569190 301195
rect 569130 301115 569190 301125
rect 569330 301185 569390 301195
rect 569330 301115 569390 301125
rect 569530 301185 569590 301195
rect 569530 301115 569590 301125
rect 569720 301185 569780 301195
rect 569720 301115 569780 301125
rect 569920 301185 569980 301195
rect 569920 301115 569980 301125
rect 570120 301185 570180 301195
rect 570120 301115 570180 301125
rect 559930 300995 559990 301005
rect 559930 300925 559990 300935
rect 560130 300995 560190 301005
rect 560130 300925 560190 300935
rect 560330 300995 560390 301005
rect 560330 300925 560390 300935
rect 560520 300995 560580 301005
rect 560520 300925 560580 300935
rect 560720 300995 560780 301005
rect 560720 300925 560780 300935
rect 560920 300995 560980 301005
rect 560920 300925 560980 300935
rect 569130 300995 569190 301005
rect 569130 300925 569190 300935
rect 569330 300995 569390 301005
rect 569330 300925 569390 300935
rect 569530 300995 569590 301005
rect 569530 300925 569590 300935
rect 569720 300995 569780 301005
rect 569720 300925 569780 300935
rect 569920 300995 569980 301005
rect 569920 300925 569980 300935
rect 570120 300995 570180 301005
rect 570120 300925 570180 300935
rect 559930 300835 559990 300845
rect 559930 300765 559990 300775
rect 560130 300835 560190 300845
rect 560130 300765 560190 300775
rect 560330 300835 560390 300845
rect 560330 300765 560390 300775
rect 560520 300835 560580 300845
rect 560520 300765 560580 300775
rect 560720 300835 560780 300845
rect 560720 300765 560780 300775
rect 560920 300835 560980 300845
rect 560920 300765 560980 300775
rect 569130 300835 569190 300845
rect 569130 300765 569190 300775
rect 569330 300835 569390 300845
rect 569330 300765 569390 300775
rect 569530 300835 569590 300845
rect 569530 300765 569590 300775
rect 569720 300835 569780 300845
rect 569720 300765 569780 300775
rect 569920 300835 569980 300845
rect 569920 300765 569980 300775
rect 570120 300835 570180 300845
rect 570120 300765 570180 300775
rect 559930 300645 559990 300655
rect 559930 300575 559990 300585
rect 560130 300645 560190 300655
rect 560130 300575 560190 300585
rect 560330 300645 560390 300655
rect 560330 300575 560390 300585
rect 560520 300645 560580 300655
rect 560520 300575 560580 300585
rect 560720 300645 560780 300655
rect 560720 300575 560780 300585
rect 560920 300645 560980 300655
rect 560920 300575 560980 300585
rect 569130 300645 569190 300655
rect 569130 300575 569190 300585
rect 569330 300645 569390 300655
rect 569330 300575 569390 300585
rect 569530 300645 569590 300655
rect 569530 300575 569590 300585
rect 569720 300645 569780 300655
rect 569720 300575 569780 300585
rect 569920 300645 569980 300655
rect 569920 300575 569980 300585
rect 570120 300645 570180 300655
rect 570120 300575 570180 300585
rect 559930 300470 559990 300480
rect 559930 300400 559990 300410
rect 560130 300470 560190 300480
rect 560130 300400 560190 300410
rect 560330 300470 560390 300480
rect 560330 300400 560390 300410
rect 560520 300470 560580 300480
rect 560520 300400 560580 300410
rect 560720 300470 560780 300480
rect 560720 300400 560780 300410
rect 560920 300470 560980 300480
rect 560920 300400 560980 300410
rect 569130 300470 569190 300480
rect 569130 300400 569190 300410
rect 569330 300470 569390 300480
rect 569330 300400 569390 300410
rect 569530 300470 569590 300480
rect 569530 300400 569590 300410
rect 569720 300470 569780 300480
rect 569720 300400 569780 300410
rect 569920 300470 569980 300480
rect 569920 300400 569980 300410
rect 570120 300470 570180 300480
rect 570120 300400 570180 300410
rect 559930 300330 559990 300340
rect 559930 300260 559990 300270
rect 560130 300330 560190 300340
rect 560130 300260 560190 300270
rect 560330 300330 560390 300340
rect 560330 300260 560390 300270
rect 560520 300330 560580 300340
rect 560520 300260 560580 300270
rect 560720 300330 560780 300340
rect 560720 300260 560780 300270
rect 560920 300330 560980 300340
rect 560920 300260 560980 300270
rect 569130 300330 569190 300340
rect 569130 300260 569190 300270
rect 569330 300330 569390 300340
rect 569330 300260 569390 300270
rect 569530 300330 569590 300340
rect 569530 300260 569590 300270
rect 569720 300330 569780 300340
rect 569720 300260 569780 300270
rect 569920 300330 569980 300340
rect 569920 300260 569980 300270
rect 570120 300330 570180 300340
rect 570120 300260 570180 300270
rect 537949 294962 538239 294982
rect 537949 294892 537969 294962
rect 538059 294892 538139 294962
rect 538229 294892 538239 294962
rect 537949 294852 538239 294892
rect 537949 294772 537969 294852
rect 538049 294772 538139 294852
rect 538219 294772 538239 294852
rect 540439 294962 540729 294982
rect 540439 294892 540459 294962
rect 540549 294892 540629 294962
rect 540719 294892 540729 294962
rect 540439 294852 540729 294892
rect 536679 294612 536969 294732
rect 537409 294722 537559 294772
rect 536679 294532 536699 294612
rect 536779 294532 536869 294612
rect 536949 294532 536969 294612
rect 537089 294682 537169 294692
rect 537089 294592 537169 294602
rect 537239 294682 537319 294692
rect 537239 294592 537319 294602
rect 537409 294652 537419 294722
rect 537549 294652 537559 294722
rect 14990 294060 15000 294200
rect 15140 294060 15150 294200
rect 15190 294060 15200 294200
rect 15340 294060 15350 294200
rect 536679 294072 536969 294532
rect 537409 294182 537559 294652
rect 536679 293992 536699 294072
rect 536779 293992 536869 294072
rect 536949 293992 536969 294072
rect 537089 294142 537169 294152
rect 537089 294052 537169 294062
rect 537239 294142 537319 294152
rect 537239 294052 537319 294062
rect 537409 294112 537419 294182
rect 537549 294112 537559 294182
rect 9670 293920 9680 293980
rect 9740 293920 9750 293980
rect 9835 293920 9845 293980
rect 9905 293920 9915 293980
rect 10035 293920 10045 293980
rect 10105 293920 10115 293980
rect 10225 293920 10235 293980
rect 10295 293920 10305 293980
rect 10405 293920 10415 293980
rect 10475 293920 10485 293980
rect 10605 293920 10615 293980
rect 10675 293920 10685 293980
rect 10795 293920 10805 293980
rect 10865 293920 10875 293980
rect 10955 293920 10965 293980
rect 11025 293920 11035 293980
rect 11145 293920 11155 293980
rect 11215 293920 11225 293980
rect 11320 293920 11330 293980
rect 11390 293920 11400 293980
rect 11460 293920 11470 293980
rect 11530 293920 11540 293980
rect 5730 293740 5740 293920
rect 5920 293740 5930 293920
rect 9670 293720 9680 293780
rect 9740 293720 9750 293780
rect 9835 293720 9845 293780
rect 9905 293720 9915 293780
rect 10035 293720 10045 293780
rect 10105 293720 10115 293780
rect 10225 293720 10235 293780
rect 10295 293720 10305 293780
rect 10405 293720 10415 293780
rect 10475 293720 10485 293780
rect 10605 293720 10615 293780
rect 10675 293720 10685 293780
rect 10795 293720 10805 293780
rect 10865 293720 10875 293780
rect 10955 293720 10965 293780
rect 11025 293720 11035 293780
rect 11145 293720 11155 293780
rect 11215 293720 11225 293780
rect 11320 293720 11330 293780
rect 11390 293720 11400 293780
rect 11460 293720 11470 293780
rect 11530 293720 11540 293780
rect 5730 293400 5740 293580
rect 5920 293400 5930 293580
rect 9670 293520 9680 293580
rect 9740 293520 9750 293580
rect 9835 293520 9845 293580
rect 9905 293520 9915 293580
rect 10035 293520 10045 293580
rect 10105 293520 10115 293580
rect 10225 293520 10235 293580
rect 10295 293520 10305 293580
rect 10405 293520 10415 293580
rect 10475 293520 10485 293580
rect 10605 293520 10615 293580
rect 10675 293520 10685 293580
rect 10795 293520 10805 293580
rect 10865 293520 10875 293580
rect 10955 293520 10965 293580
rect 11025 293520 11035 293580
rect 11145 293520 11155 293580
rect 11215 293520 11225 293580
rect 11320 293520 11330 293580
rect 11390 293520 11400 293580
rect 11460 293520 11470 293580
rect 11530 293520 11540 293580
rect 536679 293532 536969 293992
rect 537409 293642 537559 294112
rect 537949 294312 538239 294772
rect 537949 294232 537969 294312
rect 538049 294232 538139 294312
rect 538219 294232 538239 294312
rect 537949 293912 538239 294232
rect 537949 293842 537979 293912
rect 538069 293842 538119 293912
rect 538209 293842 538239 293912
rect 537949 293772 538239 293842
rect 537949 293692 537969 293772
rect 538049 293692 538139 293772
rect 538219 293692 538239 293772
rect 537949 293682 538239 293692
rect 538649 294722 538799 294782
rect 538649 294652 538659 294722
rect 538789 294652 538799 294722
rect 538649 294182 538799 294652
rect 538649 294112 538659 294182
rect 538789 294112 538799 294182
rect 536679 293452 536699 293532
rect 536779 293452 536869 293532
rect 536949 293452 536969 293532
rect 537089 293602 537169 293612
rect 537089 293512 537169 293522
rect 537239 293602 537319 293612
rect 537239 293512 537319 293522
rect 537409 293572 537419 293642
rect 537549 293572 537559 293642
rect 536679 293432 536969 293452
rect 9670 293330 9680 293390
rect 9740 293330 9750 293390
rect 9835 293330 9845 293390
rect 9905 293330 9915 293390
rect 10035 293330 10045 293390
rect 10105 293330 10115 293390
rect 10225 293330 10235 293390
rect 10295 293330 10305 293390
rect 10405 293330 10415 293390
rect 10475 293330 10485 293390
rect 10605 293330 10615 293390
rect 10675 293330 10685 293390
rect 10795 293330 10805 293390
rect 10865 293330 10875 293390
rect 10955 293330 10965 293390
rect 11025 293330 11035 293390
rect 11145 293330 11155 293390
rect 11215 293330 11225 293390
rect 11320 293330 11330 293390
rect 11390 293330 11400 293390
rect 11460 293330 11470 293390
rect 11530 293330 11540 293390
rect 5730 293060 5740 293240
rect 5920 293060 5930 293240
rect 9670 293130 9680 293190
rect 9740 293130 9750 293190
rect 9835 293130 9845 293190
rect 9905 293130 9915 293190
rect 10035 293130 10045 293190
rect 10105 293130 10115 293190
rect 10225 293130 10235 293190
rect 10295 293130 10305 293190
rect 10405 293130 10415 293190
rect 10475 293130 10485 293190
rect 10605 293130 10615 293190
rect 10675 293130 10685 293190
rect 10795 293130 10805 293190
rect 10865 293130 10875 293190
rect 10955 293130 10965 293190
rect 11025 293130 11035 293190
rect 11145 293130 11155 293190
rect 11215 293130 11225 293190
rect 11320 293130 11330 293190
rect 11390 293130 11400 293190
rect 11460 293130 11470 293190
rect 11530 293130 11540 293190
rect 537409 293102 537559 293572
rect 538649 293642 538799 294112
rect 538649 293572 538659 293642
rect 538789 293572 538799 293642
rect 537979 293382 538059 293392
rect 537979 293292 538059 293302
rect 538149 293382 538229 293392
rect 538149 293292 538229 293302
rect 537409 293032 537419 293102
rect 537549 293032 537559 293102
rect 9670 292940 9680 293000
rect 9740 292940 9750 293000
rect 536679 292992 536969 293022
rect 9835 292930 9845 292990
rect 9905 292930 9915 292990
rect 10035 292930 10045 292990
rect 10105 292930 10115 292990
rect 10225 292930 10235 292990
rect 10295 292930 10305 292990
rect 10405 292930 10415 292990
rect 10475 292930 10485 292990
rect 10605 292930 10615 292990
rect 10675 292930 10685 292990
rect 10795 292930 10805 292990
rect 10865 292930 10875 292990
rect 10955 292930 10965 292990
rect 11025 292930 11035 292990
rect 11145 292930 11155 292990
rect 11215 292930 11225 292990
rect 11320 292930 11330 292990
rect 11390 292930 11400 292990
rect 11460 292930 11470 292990
rect 11530 292930 11540 292990
rect 536679 292912 536699 292992
rect 536779 292912 536869 292992
rect 536949 292912 536969 292992
rect 14990 292720 15000 292860
rect 15140 292720 15150 292860
rect 15190 292720 15200 292860
rect 15340 292720 15350 292860
rect 536679 292412 536969 292912
rect 536679 292332 536699 292412
rect 536779 292332 536869 292412
rect 536949 292332 536969 292412
rect 530629 292132 530759 292142
rect 530629 291982 530759 291992
rect 530879 292132 531009 292142
rect 530879 291982 531009 291992
rect 536679 291802 536969 292332
rect 537409 292522 537559 293032
rect 537409 292452 537419 292522
rect 537549 292452 537559 292522
rect 537409 291942 537559 292452
rect 537959 293252 538249 293292
rect 537959 293172 537979 293252
rect 538059 293172 538149 293252
rect 538229 293172 538249 293252
rect 537959 292672 538249 293172
rect 538649 293102 538799 293572
rect 539199 294612 539489 294812
rect 540439 294772 540459 294852
rect 540539 294772 540629 294852
rect 540709 294772 540729 294852
rect 542899 294972 543189 295012
rect 542899 294892 542919 294972
rect 542999 294892 543089 294972
rect 543169 294892 543189 294972
rect 562290 294900 562300 295100
rect 562500 294900 562510 295100
rect 562690 294900 562700 295100
rect 562900 294900 562910 295100
rect 563090 294900 563100 295100
rect 563300 294900 563310 295100
rect 563490 294900 563500 295100
rect 563700 294900 563710 295100
rect 563890 294900 563900 295100
rect 564100 294900 564110 295100
rect 564290 294900 564300 295100
rect 564500 294900 564510 295100
rect 564690 294900 564700 295100
rect 564900 294900 564910 295100
rect 565090 294900 565100 295100
rect 565300 294900 565310 295100
rect 565490 294900 565500 295100
rect 565700 294900 565710 295100
rect 565890 294900 565900 295100
rect 566100 294900 566110 295100
rect 566290 294900 566300 295100
rect 566500 294900 566510 295100
rect 566690 294900 566700 295100
rect 566900 294900 566910 295100
rect 567090 294900 567100 295100
rect 567300 294900 567310 295100
rect 567490 294900 567500 295100
rect 567700 294900 567710 295100
rect 542899 294842 543189 294892
rect 539879 294722 540029 294772
rect 539199 294532 539219 294612
rect 539299 294532 539389 294612
rect 539469 294532 539489 294612
rect 539579 294682 539659 294692
rect 539579 294592 539659 294602
rect 539729 294682 539809 294692
rect 539729 294592 539809 294602
rect 539879 294652 539889 294722
rect 540019 294652 540029 294722
rect 539199 294072 539489 294532
rect 539879 294182 540029 294652
rect 539199 293992 539219 294072
rect 539299 293992 539389 294072
rect 539469 293992 539489 294072
rect 539579 294142 539659 294152
rect 539579 294052 539659 294062
rect 539729 294142 539809 294152
rect 539729 294052 539809 294062
rect 539879 294112 539889 294182
rect 540019 294112 540029 294182
rect 539199 293532 539489 293992
rect 539879 293642 540029 294112
rect 540439 294312 540729 294772
rect 540439 294232 540459 294312
rect 540539 294232 540629 294312
rect 540709 294232 540729 294312
rect 540439 293922 540729 294232
rect 540439 293912 540619 293922
rect 540439 293842 540459 293912
rect 540549 293852 540619 293912
rect 540709 293852 540729 293922
rect 540549 293842 540729 293852
rect 540439 293782 540729 293842
rect 540439 293702 540459 293782
rect 540539 293702 540629 293782
rect 540709 293702 540729 293782
rect 540439 293682 540729 293702
rect 541119 294722 541269 294772
rect 541119 294652 541129 294722
rect 541259 294652 541269 294722
rect 541119 294182 541269 294652
rect 541119 294112 541129 294182
rect 541259 294112 541269 294182
rect 539199 293452 539219 293532
rect 539299 293452 539389 293532
rect 539469 293452 539489 293532
rect 539579 293602 539659 293612
rect 539579 293512 539659 293522
rect 539729 293602 539809 293612
rect 539729 293512 539809 293522
rect 539879 293572 539889 293642
rect 540019 293572 540029 293642
rect 539199 293422 539489 293452
rect 538649 293032 538659 293102
rect 538789 293032 538799 293102
rect 539879 293102 540029 293572
rect 541119 293642 541269 294112
rect 541119 293572 541129 293642
rect 541259 293572 541269 293642
rect 540459 293382 540539 293392
rect 540629 293382 540709 293392
rect 538379 293002 538459 293012
rect 538379 292912 538459 292922
rect 538489 293002 538569 293012
rect 538489 292912 538569 292922
rect 537959 292592 537979 292672
rect 538059 292592 538149 292672
rect 538229 292592 538249 292672
rect 537959 292222 538249 292592
rect 538649 292522 538799 293032
rect 538649 292452 538659 292522
rect 538789 292452 538799 292522
rect 538379 292392 538459 292402
rect 538379 292302 538459 292312
rect 538489 292392 538569 292402
rect 538489 292302 538569 292312
rect 537959 292142 537979 292222
rect 538069 292142 538139 292222
rect 538229 292142 538249 292222
rect 537959 292092 538249 292142
rect 537959 292012 537979 292092
rect 538059 292012 538149 292092
rect 538229 292012 538249 292092
rect 537959 291992 538249 292012
rect 537409 291872 537419 291942
rect 537549 291872 537559 291942
rect 537409 291832 537559 291872
rect 538649 291942 538799 292452
rect 538649 291872 538659 291942
rect 538789 291872 538799 291942
rect 534849 291652 535139 291732
rect 536759 291722 536889 291802
rect 538359 291752 538589 291842
rect 538649 291792 538799 291872
rect 539181 292992 539513 293042
rect 539181 292912 539209 292992
rect 539289 292912 539379 292992
rect 539459 292912 539513 292992
rect 539181 292412 539513 292912
rect 539181 292332 539209 292412
rect 539289 292332 539379 292412
rect 539459 292332 539513 292412
rect 539181 291832 539513 292332
rect 539879 293032 539889 293102
rect 540019 293032 540029 293102
rect 539879 292522 540029 293032
rect 539879 292452 539899 292522
rect 539879 291942 540029 292452
rect 540439 293262 540729 293302
rect 540439 293182 540459 293262
rect 540539 293182 540629 293262
rect 540709 293182 540729 293262
rect 540439 292682 540729 293182
rect 541119 293102 541269 293572
rect 541689 294612 541979 294812
rect 542899 294762 542919 294842
rect 542999 294762 543089 294842
rect 543169 294762 543189 294842
rect 542359 294722 542509 294762
rect 541689 294532 541709 294612
rect 541789 294532 541879 294612
rect 541959 294532 541979 294612
rect 542059 294682 542139 294692
rect 542059 294592 542139 294602
rect 542209 294682 542289 294692
rect 542209 294592 542289 294602
rect 542359 294652 542369 294722
rect 542499 294652 542509 294722
rect 541689 294072 541979 294532
rect 542359 294432 542509 294652
rect 542349 294182 542509 294432
rect 541689 293992 541709 294072
rect 541789 293992 541879 294072
rect 541959 293992 541979 294072
rect 542059 294142 542139 294152
rect 542059 294052 542139 294062
rect 542209 294142 542289 294152
rect 542209 294052 542289 294062
rect 542349 294112 542369 294182
rect 542499 294112 542509 294182
rect 541689 293522 541979 293992
rect 542349 293642 542509 294112
rect 541689 293442 541709 293522
rect 541789 293442 541879 293522
rect 541959 293442 541979 293522
rect 542069 293602 542149 293612
rect 542069 293512 542149 293522
rect 542209 293602 542289 293612
rect 542209 293512 542289 293522
rect 542349 293572 542369 293642
rect 542499 293572 542509 293642
rect 542349 293532 542509 293572
rect 542899 294302 543189 294762
rect 542899 294222 542919 294302
rect 542999 294222 543089 294302
rect 543169 294222 543189 294302
rect 542899 293922 543189 294222
rect 542899 293852 542919 293922
rect 542999 293852 543089 293922
rect 543169 293852 543189 293922
rect 542899 293762 543189 293852
rect 542899 293682 542919 293762
rect 542999 293682 543089 293762
rect 543169 293682 543189 293762
rect 541689 293422 541979 293442
rect 541119 293032 541129 293102
rect 541259 293032 541269 293102
rect 542349 293102 542499 293532
rect 542899 293432 543189 293682
rect 543589 294722 543739 294752
rect 543589 294652 543599 294722
rect 543729 294652 543739 294722
rect 543589 294182 543739 294652
rect 543589 294112 543599 294182
rect 543729 294112 543739 294182
rect 543589 293642 543739 294112
rect 543589 293572 543599 293642
rect 543729 293572 543739 293642
rect 542919 293382 542999 293392
rect 543089 293382 543169 293392
rect 542349 293032 542359 293102
rect 542489 293032 542499 293102
rect 540789 293002 540869 293012
rect 540789 292912 540869 292922
rect 540899 293002 540979 293012
rect 540899 292912 540979 292922
rect 540439 292602 540459 292682
rect 540539 292602 540629 292682
rect 540709 292602 540729 292682
rect 540439 292212 540729 292602
rect 541119 292522 541269 293032
rect 541119 292452 541129 292522
rect 541259 292452 541269 292522
rect 540789 292412 540869 292422
rect 540789 292322 540869 292332
rect 540899 292412 540979 292422
rect 540899 292322 540979 292332
rect 540439 292142 540459 292212
rect 540539 292142 540629 292212
rect 540709 292142 540729 292212
rect 540439 292102 540729 292142
rect 540439 292022 540459 292102
rect 540539 292022 540629 292102
rect 540709 292022 540729 292102
rect 540439 292002 540729 292022
rect 539879 291872 539889 291942
rect 540019 291872 540029 291942
rect 539879 291842 540029 291872
rect 541119 291942 541269 292452
rect 541119 291872 541129 291942
rect 541259 291872 541269 291942
rect 541119 291842 541269 291872
rect 541679 292992 541969 293032
rect 541679 292912 541699 292992
rect 541779 292912 541869 292992
rect 541949 292912 541969 292992
rect 541679 292402 541969 292912
rect 541679 292322 541699 292402
rect 541779 292322 541869 292402
rect 541949 292322 541969 292402
rect 539181 291752 539209 291832
rect 539289 291752 539379 291832
rect 539459 291752 539513 291832
rect 536679 291712 536759 291722
rect 536889 291712 536969 291722
rect 539181 291694 539513 291752
rect 540789 291832 540869 291842
rect 540789 291742 540869 291752
rect 540899 291832 540979 291842
rect 540899 291742 540979 291752
rect 541679 291832 541969 292322
rect 542349 292522 542499 293032
rect 542349 292452 542359 292522
rect 542489 292452 542499 292522
rect 542349 291942 542499 292452
rect 542899 293252 543189 293302
rect 542899 293172 542919 293252
rect 542999 293172 543089 293252
rect 543169 293172 543189 293252
rect 542899 292672 543189 293172
rect 543589 293102 543739 293572
rect 544139 294612 544429 294882
rect 544139 294532 544159 294612
rect 544239 294532 544329 294612
rect 544409 294532 544429 294612
rect 544139 294062 544429 294532
rect 562290 294500 562300 294700
rect 562500 294500 562510 294700
rect 562690 294500 562700 294700
rect 562900 294500 562910 294700
rect 563090 294500 563100 294700
rect 563300 294500 563310 294700
rect 563490 294500 563500 294700
rect 563700 294500 563710 294700
rect 563890 294500 563900 294700
rect 564100 294500 564110 294700
rect 564290 294500 564300 294700
rect 564500 294500 564510 294700
rect 564690 294500 564700 294700
rect 564900 294500 564910 294700
rect 565090 294500 565100 294700
rect 565300 294500 565310 294700
rect 565490 294500 565500 294700
rect 565700 294500 565710 294700
rect 565890 294500 565900 294700
rect 566100 294500 566110 294700
rect 566290 294500 566300 294700
rect 566500 294500 566510 294700
rect 566690 294500 566700 294700
rect 566900 294500 566910 294700
rect 567090 294500 567100 294700
rect 567300 294500 567310 294700
rect 567490 294500 567500 294700
rect 567700 294500 567710 294700
rect 562290 294100 562300 294300
rect 562500 294100 562510 294300
rect 562690 294100 562700 294300
rect 562900 294100 562910 294300
rect 563090 294100 563100 294300
rect 563300 294100 563310 294300
rect 563490 294100 563500 294300
rect 563700 294100 563710 294300
rect 563890 294100 563900 294300
rect 564100 294100 564110 294300
rect 564290 294100 564300 294300
rect 564500 294100 564510 294300
rect 564690 294100 564700 294300
rect 564900 294100 564910 294300
rect 565090 294100 565100 294300
rect 565300 294100 565310 294300
rect 565490 294100 565500 294300
rect 565700 294100 565710 294300
rect 565890 294100 565900 294300
rect 566100 294100 566110 294300
rect 566290 294100 566300 294300
rect 566500 294100 566510 294300
rect 566690 294100 566700 294300
rect 566900 294100 566910 294300
rect 567090 294100 567100 294300
rect 567300 294100 567310 294300
rect 567490 294100 567500 294300
rect 567700 294100 567710 294300
rect 544139 293982 544159 294062
rect 544239 293982 544329 294062
rect 544409 293982 544429 294062
rect 544139 293532 544429 293982
rect 562290 293700 562300 293900
rect 562500 293700 562510 293900
rect 562690 293700 562700 293900
rect 562900 293700 562910 293900
rect 563090 293700 563100 293900
rect 563300 293700 563310 293900
rect 563490 293700 563500 293900
rect 563700 293700 563710 293900
rect 563890 293700 563900 293900
rect 564100 293700 564110 293900
rect 564290 293700 564300 293900
rect 564500 293700 564510 293900
rect 564690 293700 564700 293900
rect 564900 293700 564910 293900
rect 565090 293700 565100 293900
rect 565300 293700 565310 293900
rect 565490 293700 565500 293900
rect 565700 293700 565710 293900
rect 565890 293700 565900 293900
rect 566100 293700 566110 293900
rect 566290 293700 566300 293900
rect 566500 293700 566510 293900
rect 566690 293700 566700 293900
rect 566900 293700 566910 293900
rect 567090 293700 567100 293900
rect 567300 293700 567310 293900
rect 567490 293700 567500 293900
rect 567700 293700 567710 293900
rect 544139 293452 544159 293532
rect 544239 293452 544329 293532
rect 544409 293452 544429 293532
rect 544139 293442 544429 293452
rect 562290 293300 562300 293500
rect 562500 293300 562510 293500
rect 562690 293300 562700 293500
rect 562900 293300 562910 293500
rect 563090 293300 563100 293500
rect 563300 293300 563310 293500
rect 563490 293300 563500 293500
rect 563700 293300 563710 293500
rect 563890 293300 563900 293500
rect 564100 293300 564110 293500
rect 564290 293300 564300 293500
rect 564500 293300 564510 293500
rect 564690 293300 564700 293500
rect 564900 293300 564910 293500
rect 565090 293300 565100 293500
rect 565300 293300 565310 293500
rect 565490 293300 565500 293500
rect 565700 293300 565710 293500
rect 565890 293300 565900 293500
rect 566100 293300 566110 293500
rect 566290 293300 566300 293500
rect 566500 293300 566510 293500
rect 566690 293300 566700 293500
rect 566900 293300 566910 293500
rect 567090 293300 567100 293500
rect 567300 293300 567310 293500
rect 567490 293300 567500 293500
rect 567700 293300 567710 293500
rect 543589 293032 543599 293102
rect 543729 293032 543739 293102
rect 543249 292992 543329 293002
rect 543249 292902 543329 292912
rect 543359 292992 543439 293002
rect 543359 292902 543439 292912
rect 542899 292592 542919 292672
rect 542999 292592 543089 292672
rect 543169 292592 543189 292672
rect 542899 292212 543189 292592
rect 543589 292522 543739 293032
rect 543589 292452 543599 292522
rect 543729 292452 543739 292522
rect 543249 292412 543329 292422
rect 543249 292322 543329 292332
rect 543359 292412 543439 292422
rect 543359 292322 543439 292332
rect 542899 292142 542919 292212
rect 542999 292142 543089 292212
rect 543169 292142 543189 292212
rect 542899 292092 543189 292142
rect 542899 292012 542919 292092
rect 542999 292012 543089 292092
rect 543169 292012 543189 292092
rect 542899 292002 543189 292012
rect 542349 291872 542359 291942
rect 542489 291872 542499 291942
rect 542349 291832 542499 291872
rect 543589 291942 543739 292452
rect 543589 291872 543599 291942
rect 543729 291872 543739 291942
rect 543589 291842 543739 291872
rect 544169 292992 544459 293082
rect 544169 292912 544189 292992
rect 544269 292912 544359 292992
rect 544439 292912 544459 292992
rect 544169 292412 544459 292912
rect 544169 292332 544189 292412
rect 544269 292332 544359 292412
rect 544439 292332 544459 292412
rect 543249 291832 543329 291842
rect 541679 291752 541699 291832
rect 541779 291752 541869 291832
rect 541949 291752 541969 291832
rect 541679 291732 541969 291752
rect 543249 291742 543329 291752
rect 543359 291832 543439 291842
rect 543359 291742 543439 291752
rect 544169 291832 544459 292332
rect 550129 292302 550259 292312
rect 550129 292152 550259 292162
rect 550389 292302 550519 292312
rect 550389 292152 550519 292162
rect 544169 291752 544189 291832
rect 544269 291752 544359 291832
rect 544439 291752 544459 291832
rect 544169 291732 544459 291752
rect 534849 291542 534869 291652
rect 534959 291542 535029 291652
rect 535119 291542 535139 291652
rect 544779 291602 545069 291642
rect 534849 291282 535139 291542
rect 536099 291562 536409 291582
rect 536179 291482 536329 291562
rect 534929 291202 535059 291282
rect 533080 290940 533140 290950
rect 533080 290870 533140 290880
rect 533180 290940 533240 290950
rect 533180 290870 533240 290880
rect 533280 290940 533340 290950
rect 533280 290870 533340 290880
rect 533060 290820 533360 290840
rect 533060 290760 533080 290820
rect 533140 290760 533180 290820
rect 533240 290760 533280 290820
rect 533340 290760 533360 290820
rect 533060 290720 533360 290760
rect 533060 290660 533080 290720
rect 533140 290660 533180 290720
rect 533240 290660 533280 290720
rect 533340 290660 533360 290720
rect 533060 290580 533360 290660
rect 533060 290520 533080 290580
rect 533140 290520 533180 290580
rect 533240 290520 533280 290580
rect 533340 290520 533360 290580
rect 533060 290480 533360 290520
rect 533060 290420 533080 290480
rect 533140 290420 533180 290480
rect 533240 290420 533280 290480
rect 533340 290420 533360 290480
rect 533060 290380 533360 290420
rect 533060 290320 533080 290380
rect 533140 290320 533180 290380
rect 533240 290320 533280 290380
rect 533340 290320 533360 290380
rect 533060 290280 533360 290320
rect 533060 290220 533080 290280
rect 533140 290220 533180 290280
rect 533240 290220 533280 290280
rect 533340 290220 533360 290280
rect 533060 290180 533360 290220
rect 534849 290742 535139 291202
rect 534929 290662 535059 290742
rect 534849 290202 535139 290662
rect 534929 290122 535059 290202
rect 534849 289662 535139 290122
rect 535569 291402 535719 291432
rect 535569 291332 535579 291402
rect 535709 291332 535719 291402
rect 535569 290872 535719 291332
rect 535569 290802 535579 290872
rect 535709 290802 535719 290872
rect 535569 290322 535719 290802
rect 535569 290252 535579 290322
rect 535709 290252 535719 290322
rect 535569 289782 535719 290252
rect 536099 291142 536409 291482
rect 538629 291552 538919 291582
rect 538629 291472 538649 291552
rect 538729 291472 538819 291552
rect 538899 291472 538919 291552
rect 536099 291062 536119 291142
rect 536209 291062 536299 291142
rect 536389 291062 536409 291142
rect 536099 291022 536409 291062
rect 536179 290942 536329 291022
rect 536099 290482 536409 290942
rect 536179 290402 536329 290482
rect 536099 290072 536409 290402
rect 536099 290062 536299 290072
rect 536099 289982 536119 290062
rect 536209 289992 536299 290062
rect 536389 289992 536409 290072
rect 536209 289982 536409 289992
rect 536099 289932 536409 289982
rect 536179 289852 536329 289932
rect 536099 289842 536409 289852
rect 536809 291402 536959 291442
rect 536809 291332 536819 291402
rect 536949 291332 536959 291402
rect 536809 290862 536959 291332
rect 538039 291402 538189 291432
rect 538039 291332 538049 291402
rect 538179 291332 538189 291402
rect 536809 290792 536819 290862
rect 536949 290792 536959 290862
rect 536809 290322 536959 290792
rect 536809 290252 536819 290322
rect 536949 290252 536959 290322
rect 535569 289712 535579 289782
rect 535709 289712 535719 289782
rect 535569 289672 535719 289712
rect 536809 289782 536959 290252
rect 536809 289712 536819 289782
rect 536949 289712 536959 289782
rect 534929 289582 535059 289662
rect 534849 289572 535139 289582
rect 531759 289252 531849 289262
rect 531759 289112 531849 289122
rect 531969 289252 532059 289262
rect 531969 289112 532059 289122
rect 536809 289132 536959 289712
rect 537319 291282 537639 291312
rect 537319 291202 537329 291282
rect 537409 291202 537549 291282
rect 537629 291202 537639 291282
rect 537319 290742 537639 291202
rect 537319 290662 537329 290742
rect 537409 290662 537549 290742
rect 537629 290662 537639 290742
rect 537319 290202 537639 290662
rect 537399 290122 537559 290202
rect 537319 289732 537639 290122
rect 538039 290862 538189 291332
rect 538039 290792 538049 290862
rect 538179 290792 538189 290862
rect 538039 290322 538189 290792
rect 538039 290252 538049 290322
rect 538179 290252 538189 290322
rect 538039 289782 538189 290252
rect 538629 291142 538919 291472
rect 541099 291552 541389 291592
rect 541099 291472 541109 291552
rect 541189 291472 541299 291552
rect 541379 291472 541389 291552
rect 538629 291062 538649 291142
rect 538739 291062 538809 291142
rect 538899 291062 538919 291142
rect 538629 291022 538919 291062
rect 538629 291012 538819 291022
rect 538629 290932 538649 291012
rect 538729 290942 538819 291012
rect 538899 290942 538919 291022
rect 538729 290932 538919 290942
rect 538629 290472 538919 290932
rect 538629 290392 538639 290472
rect 538719 290392 538809 290472
rect 538889 290392 538919 290472
rect 538629 290062 538919 290392
rect 538629 289982 538649 290062
rect 538739 289982 538809 290062
rect 538899 289982 538919 290062
rect 538629 289942 538919 289982
rect 538709 289862 538819 289942
rect 538899 289862 538919 289942
rect 538629 289832 538919 289862
rect 539279 291402 539429 291432
rect 539279 291332 539289 291402
rect 539419 291332 539429 291402
rect 540519 291402 540669 291422
rect 539279 290862 539429 291332
rect 539279 290792 539289 290862
rect 539419 290792 539429 290862
rect 539279 290322 539429 290792
rect 539279 290252 539289 290322
rect 539419 290252 539429 290322
rect 537319 289652 537729 289732
rect 537399 289572 537559 289652
rect 537639 289572 537729 289652
rect 537319 289472 537729 289572
rect 536809 289062 536819 289132
rect 536949 289062 536959 289132
rect 536809 289052 536959 289062
rect 536759 288862 536849 288872
rect 536899 288862 536989 288872
rect 536849 288782 536899 288852
rect 536759 288632 536989 288782
rect 536849 288552 536899 288632
rect 536759 286582 536989 288552
rect 537069 288372 537339 288382
rect 537069 288292 537089 288372
rect 537169 288292 537239 288372
rect 537319 288292 537339 288372
rect 537089 288282 537169 288292
rect 537239 288282 537319 288292
rect 537539 288172 537729 289472
rect 538039 289712 538049 289782
rect 538179 289712 538189 289782
rect 538039 289122 538189 289712
rect 539279 289782 539429 290252
rect 539279 289712 539289 289782
rect 539419 289712 539429 289782
rect 538039 289052 538049 289122
rect 538179 289052 538189 289122
rect 538039 289002 538189 289052
rect 538379 289132 538459 289142
rect 538379 289042 538459 289052
rect 538489 289132 538569 289142
rect 538489 289042 538569 289052
rect 539279 289122 539429 289712
rect 539279 289052 539289 289122
rect 539419 289052 539429 289122
rect 539279 288962 539429 289052
rect 539849 291282 540139 291372
rect 539849 291202 539859 291282
rect 539939 291202 540039 291282
rect 540119 291202 540139 291282
rect 539849 290742 540139 291202
rect 539849 290662 539859 290742
rect 539939 290662 540049 290742
rect 540129 290662 540139 290742
rect 539849 290202 540139 290662
rect 539849 290122 539859 290202
rect 539939 290122 540039 290202
rect 540119 290122 540139 290202
rect 539849 289662 540139 290122
rect 539849 289582 539859 289662
rect 539939 289582 540049 289662
rect 540129 289582 540139 289662
rect 538279 288772 538389 288782
rect 538279 288652 538389 288662
rect 539139 288772 539249 288782
rect 539139 288652 539249 288662
rect 539579 288392 539659 288402
rect 539579 288302 539659 288312
rect 539729 288392 539809 288402
rect 539729 288302 539809 288312
rect 537449 288142 537759 288172
rect 537449 288062 537539 288142
rect 537619 288062 537649 288142
rect 537729 288062 537759 288142
rect 539849 288112 540139 289582
rect 540519 291332 540529 291402
rect 540659 291332 540669 291402
rect 540519 290862 540669 291332
rect 540519 290792 540529 290862
rect 540659 290792 540669 290862
rect 540519 290322 540669 290792
rect 540519 290252 540529 290322
rect 540659 290252 540669 290322
rect 540519 289782 540669 290252
rect 541099 291142 541389 291472
rect 543549 291552 543839 291582
rect 543549 291472 543559 291552
rect 543639 291472 543749 291552
rect 543829 291472 543839 291552
rect 541099 291062 541119 291142
rect 541209 291062 541279 291142
rect 541369 291062 541389 291142
rect 541099 291022 541389 291062
rect 541099 290942 541109 291022
rect 541189 290942 541299 291022
rect 541379 290942 541389 291022
rect 541099 290472 541389 290942
rect 541099 290392 541109 290472
rect 541189 290392 541289 290472
rect 541369 290392 541389 290472
rect 541099 290062 541389 290392
rect 541099 289982 541119 290062
rect 541209 289982 541279 290062
rect 541369 289982 541389 290062
rect 541099 289932 541389 289982
rect 541099 289852 541109 289932
rect 541189 289852 541299 289932
rect 541379 289852 541389 289932
rect 541099 289842 541389 289852
rect 541749 291402 541899 291432
rect 541749 291332 541759 291402
rect 541889 291332 541899 291402
rect 542989 291402 543139 291452
rect 541749 290862 541899 291332
rect 541749 290792 541759 290862
rect 541889 290792 541899 290862
rect 541749 290322 541899 290792
rect 541749 290252 541759 290322
rect 541889 290252 541899 290322
rect 540519 289712 540529 289782
rect 540659 289712 540669 289782
rect 540519 289122 540669 289712
rect 541749 289782 541899 290252
rect 541749 289712 541759 289782
rect 541889 289712 541899 289782
rect 540519 289052 540529 289122
rect 540659 289052 540669 289122
rect 540519 288982 540669 289052
rect 540789 289132 540869 289142
rect 540789 289042 540869 289052
rect 540899 289132 540979 289142
rect 540899 289042 540979 289052
rect 541749 289122 541899 289712
rect 542309 291272 542599 291372
rect 542309 291192 542319 291272
rect 542399 291192 542499 291272
rect 542579 291192 542599 291272
rect 542309 290732 542599 291192
rect 542309 290652 542319 290732
rect 542399 290652 542499 290732
rect 542579 290652 542599 290732
rect 542309 290192 542599 290652
rect 542309 290112 542329 290192
rect 542409 290112 542499 290192
rect 542579 290112 542599 290192
rect 542309 289752 542599 290112
rect 542989 291332 542999 291402
rect 543129 291332 543139 291402
rect 542989 290862 543139 291332
rect 542989 290792 542999 290862
rect 543129 290792 543139 290862
rect 542989 290322 543139 290792
rect 542989 290252 542999 290322
rect 543129 290252 543139 290322
rect 542989 289782 543139 290252
rect 542309 289652 542609 289752
rect 542309 289572 542319 289652
rect 542399 289572 542509 289652
rect 542589 289572 542609 289652
rect 542309 289552 542609 289572
rect 541749 289052 541759 289122
rect 541889 289052 541899 289122
rect 541749 289042 541899 289052
rect 541769 288882 541859 288892
rect 541909 288882 541999 288892
rect 541859 288802 541909 288882
rect 540349 288772 540459 288782
rect 540349 288652 540459 288662
rect 541199 288772 541309 288782
rect 541199 288652 541309 288662
rect 539849 288062 539949 288112
rect 537449 288042 537759 288062
rect 540029 288062 540139 288112
rect 541769 288622 541999 288802
rect 541859 288542 541909 288622
rect 538719 287962 538799 287992
rect 537459 287782 537539 287812
rect 537459 287692 537539 287702
rect 537459 287652 537719 287692
rect 537459 287562 537569 287652
rect 537679 287562 537719 287652
rect 537459 287522 537719 287562
rect 537459 287162 537539 287522
rect 537459 287072 537539 287082
rect 538109 287342 538319 287362
rect 538199 287262 538229 287342
rect 536849 286502 536899 286582
rect 536759 285962 536989 286502
rect 538109 286742 538319 287262
rect 538719 287342 538799 287882
rect 539949 287492 540029 288032
rect 539949 287402 540029 287412
rect 541129 287962 541209 287992
rect 538719 287252 538799 287262
rect 540559 287342 540769 287362
rect 540649 287262 540679 287342
rect 538199 286662 538229 286742
rect 537509 286452 537629 286462
rect 537509 286342 537629 286352
rect 538109 286142 538319 286662
rect 539339 286912 539429 286942
rect 538729 286452 538849 286462
rect 538729 286342 538849 286352
rect 539339 286312 539429 286832
rect 540559 286742 540769 287262
rect 541129 287342 541209 287882
rect 541129 287252 541209 287262
rect 540649 286662 540679 286742
rect 539939 286452 540059 286462
rect 539939 286342 540059 286352
rect 539339 286222 539429 286232
rect 540559 286196 540769 286662
rect 541769 286582 541999 288542
rect 542059 288392 542139 288402
rect 542059 288302 542139 288312
rect 542199 288392 542279 288402
rect 542199 288302 542279 288312
rect 542389 288132 542609 289552
rect 542989 289712 542999 289782
rect 543129 289712 543139 289782
rect 542989 289142 543139 289712
rect 543549 291142 543839 291472
rect 544779 291522 544799 291602
rect 544879 291522 544969 291602
rect 545049 291522 545069 291602
rect 543549 291062 543569 291142
rect 543659 291062 543729 291142
rect 543819 291062 543839 291142
rect 543549 291012 543839 291062
rect 543549 290932 543559 291012
rect 543639 290932 543749 291012
rect 543829 290932 543839 291012
rect 543549 290472 543839 290932
rect 543549 290392 543559 290472
rect 543639 290392 543749 290472
rect 543829 290392 543839 290472
rect 543549 290062 543839 290392
rect 543549 289982 543569 290062
rect 543659 289982 543729 290062
rect 543819 289982 543839 290062
rect 543549 289932 543839 289982
rect 543549 289852 543559 289932
rect 543639 289852 543749 289932
rect 543829 289852 543839 289932
rect 543549 289602 543839 289852
rect 544219 291402 544369 291442
rect 544219 291332 544229 291402
rect 544359 291332 544369 291402
rect 544219 290862 544369 291332
rect 544219 290792 544229 290862
rect 544359 290792 544369 290862
rect 544219 290322 544369 290792
rect 544219 290252 544229 290322
rect 544359 290252 544369 290322
rect 544219 289782 544369 290252
rect 544219 289712 544229 289782
rect 544359 289712 544369 289782
rect 542989 289072 542999 289142
rect 543129 289072 543139 289142
rect 542989 289012 543139 289072
rect 543249 289142 543329 289152
rect 543249 289052 543329 289062
rect 543359 289142 543439 289152
rect 543359 289052 543439 289062
rect 544219 289122 544369 289712
rect 544779 291272 545069 291522
rect 546049 291552 546339 291572
rect 546049 291472 546069 291552
rect 546149 291472 546239 291552
rect 546319 291472 546339 291552
rect 544779 291192 544799 291272
rect 544879 291192 544969 291272
rect 545049 291192 545069 291272
rect 544779 290732 545069 291192
rect 544779 290652 544799 290732
rect 544879 290652 544969 290732
rect 545049 290652 545069 290732
rect 544779 290192 545069 290652
rect 544779 290112 544799 290192
rect 544879 290112 544969 290192
rect 545049 290112 545069 290192
rect 544779 289642 545069 290112
rect 545459 291402 545609 291442
rect 545459 291332 545469 291402
rect 545599 291332 545609 291402
rect 545459 290862 545609 291332
rect 545459 290792 545469 290862
rect 545599 290792 545609 290862
rect 545459 290322 545609 290792
rect 545459 290252 545469 290322
rect 545599 290252 545609 290322
rect 545459 289782 545609 290252
rect 546049 291142 546339 291472
rect 546049 291062 546069 291142
rect 546159 291062 546229 291142
rect 546319 291062 546339 291142
rect 546049 291012 546339 291062
rect 546049 290932 546069 291012
rect 546149 290932 546239 291012
rect 546319 290932 546339 291012
rect 546049 290472 546339 290932
rect 546049 290392 546069 290472
rect 546149 290392 546239 290472
rect 546319 290392 546339 290472
rect 546049 290062 546339 290392
rect 546049 289982 546069 290062
rect 546159 289982 546229 290062
rect 546319 289982 546339 290062
rect 546049 289922 546339 289982
rect 546049 289842 546069 289922
rect 546149 289842 546239 289922
rect 546319 289842 546339 289922
rect 546049 289822 546339 289842
rect 545459 289712 545469 289782
rect 545599 289712 545609 289782
rect 545459 289682 545609 289712
rect 544779 289562 544799 289642
rect 544879 289562 544969 289642
rect 545049 289562 545069 289642
rect 544779 289552 545069 289562
rect 549069 289242 549139 289252
rect 549069 289142 549139 289152
rect 549229 289242 549299 289252
rect 549229 289142 549299 289152
rect 544219 289052 544229 289122
rect 544359 289052 544369 289122
rect 544219 289012 544369 289052
rect 542769 288772 542879 288782
rect 542769 288652 542879 288662
rect 543649 288772 543759 288782
rect 572740 288704 572750 288764
rect 572810 288704 572820 288764
rect 572880 288704 572890 288764
rect 572950 288704 572960 288764
rect 573055 288704 573065 288764
rect 573125 288704 573135 288764
rect 573245 288704 573255 288764
rect 573315 288704 573325 288764
rect 573405 288704 573415 288764
rect 573475 288704 573485 288764
rect 573595 288704 573605 288764
rect 573665 288704 573675 288764
rect 573795 288704 573805 288764
rect 573865 288704 573875 288764
rect 573975 288704 573985 288764
rect 574045 288704 574055 288764
rect 574165 288704 574175 288764
rect 574235 288704 574245 288764
rect 574365 288704 574375 288764
rect 574435 288704 574445 288764
rect 574530 288694 574540 288754
rect 574600 288694 574610 288754
rect 543649 288652 543759 288662
rect 578360 288600 578440 288610
rect 572740 288504 572750 288564
rect 572810 288504 572820 288564
rect 572880 288504 572890 288564
rect 572950 288504 572960 288564
rect 573055 288504 573065 288564
rect 573125 288504 573135 288564
rect 573245 288504 573255 288564
rect 573315 288504 573325 288564
rect 573405 288504 573415 288564
rect 573475 288504 573485 288564
rect 573595 288504 573605 288564
rect 573665 288504 573675 288564
rect 573795 288504 573805 288564
rect 573865 288504 573875 288564
rect 573975 288504 573985 288564
rect 574045 288504 574055 288564
rect 574165 288504 574175 288564
rect 574235 288504 574245 288564
rect 574365 288504 574375 288564
rect 574435 288504 574445 288564
rect 574530 288504 574540 288564
rect 574600 288504 574610 288564
rect 578360 288510 578440 288520
rect 578540 288600 578620 288610
rect 578540 288510 578620 288520
rect 578360 288440 578440 288450
rect 572740 288304 572750 288364
rect 572810 288304 572820 288364
rect 572880 288304 572890 288364
rect 572950 288304 572960 288364
rect 573055 288304 573065 288364
rect 573125 288304 573135 288364
rect 573245 288304 573255 288364
rect 573315 288304 573325 288364
rect 573405 288304 573415 288364
rect 573475 288304 573485 288364
rect 573595 288304 573605 288364
rect 573665 288304 573675 288364
rect 573795 288304 573805 288364
rect 573865 288304 573875 288364
rect 573975 288304 573985 288364
rect 574045 288304 574055 288364
rect 574165 288304 574175 288364
rect 574235 288304 574245 288364
rect 574365 288304 574375 288364
rect 574435 288304 574445 288364
rect 574530 288304 574540 288364
rect 574600 288304 574610 288364
rect 578360 288350 578440 288360
rect 578540 288440 578620 288450
rect 578540 288350 578620 288360
rect 578360 288280 578440 288290
rect 578360 288190 578440 288200
rect 578540 288280 578620 288290
rect 578540 288190 578620 288200
rect 542389 288052 542399 288132
rect 542479 288052 542519 288132
rect 542599 288052 542609 288132
rect 543549 288122 543839 288132
rect 543549 288082 543599 288122
rect 542389 288042 542609 288052
rect 543679 288082 543839 288122
rect 572740 288114 572750 288174
rect 572810 288114 572820 288174
rect 572880 288114 572890 288174
rect 572950 288114 572960 288174
rect 573055 288114 573065 288174
rect 573125 288114 573135 288174
rect 573245 288114 573255 288174
rect 573315 288114 573325 288174
rect 573405 288114 573415 288174
rect 573475 288114 573485 288174
rect 573595 288114 573605 288174
rect 573665 288114 573675 288174
rect 573795 288114 573805 288174
rect 573865 288114 573875 288174
rect 573975 288114 573985 288174
rect 574045 288114 574055 288174
rect 574165 288114 574175 288174
rect 574235 288114 574245 288174
rect 574365 288114 574375 288174
rect 574435 288114 574445 288174
rect 574530 288114 574540 288174
rect 574600 288114 574610 288174
rect 578360 288100 578440 288110
rect 542349 287782 542429 287812
rect 542349 287692 542429 287702
rect 542349 287652 542619 287692
rect 542349 287562 542479 287652
rect 542589 287562 542619 287652
rect 542349 287522 542619 287562
rect 542349 287162 542429 287522
rect 543599 287502 543679 288042
rect 578360 288010 578440 288020
rect 578540 288100 578620 288110
rect 578540 288010 578620 288020
rect 572740 287914 572750 287974
rect 572810 287914 572820 287974
rect 572880 287914 572890 287974
rect 572950 287914 572960 287974
rect 573055 287914 573065 287974
rect 573125 287914 573135 287974
rect 573245 287914 573255 287974
rect 573315 287914 573325 287974
rect 573405 287914 573415 287974
rect 573475 287914 573485 287974
rect 573595 287914 573605 287974
rect 573665 287914 573675 287974
rect 573795 287914 573805 287974
rect 573865 287914 573875 287974
rect 573975 287914 573985 287974
rect 574045 287914 574055 287974
rect 574165 287914 574175 287974
rect 574235 287914 574245 287974
rect 574365 287914 574375 287974
rect 574435 287914 574445 287974
rect 574530 287914 574540 287974
rect 574600 287914 574610 287974
rect 578360 287940 578440 287950
rect 578360 287850 578440 287860
rect 578540 287940 578620 287950
rect 578540 287850 578620 287860
rect 572740 287714 572750 287774
rect 572810 287714 572820 287774
rect 572880 287714 572890 287774
rect 572950 287714 572960 287774
rect 573055 287714 573065 287774
rect 573125 287714 573135 287774
rect 573245 287714 573255 287774
rect 573315 287714 573325 287774
rect 573405 287714 573415 287774
rect 573475 287714 573485 287774
rect 573595 287714 573605 287774
rect 573665 287714 573675 287774
rect 573795 287714 573805 287774
rect 573865 287714 573875 287774
rect 573975 287714 573985 287774
rect 574045 287714 574055 287774
rect 574165 287714 574175 287774
rect 574235 287714 574245 287774
rect 574365 287714 574375 287774
rect 574435 287714 574445 287774
rect 574530 287714 574540 287774
rect 574600 287714 574610 287774
rect 543599 287412 543679 287422
rect 542349 287072 542429 287082
rect 542989 287342 543199 287362
rect 543079 287262 543109 287342
rect 541859 286502 541909 286582
rect 541159 286452 541279 286462
rect 541159 286342 541279 286352
rect 538199 286062 538229 286142
rect 538109 286052 538319 286062
rect 540390 286146 540790 286196
rect 540390 286056 540420 286146
rect 540508 286142 540790 286146
rect 540508 286062 540559 286142
rect 540649 286062 540679 286142
rect 540769 286062 540790 286142
rect 540508 286056 540790 286062
rect 536849 285882 536899 285962
rect 536759 285872 536989 285882
rect 537384 285478 537544 285488
rect 537384 285308 537544 285318
rect 538444 285478 538604 285488
rect 538444 285308 538604 285318
rect 539904 285478 540064 285488
rect 539904 285308 540064 285318
rect 538864 285088 538884 285158
rect 538954 285088 539104 285158
rect 539174 285088 539194 285158
rect 537384 284898 537544 284908
rect 537384 284728 537544 284738
rect 538444 284898 538604 284908
rect 538444 284728 538604 284738
rect 538864 284568 539194 285088
rect 539904 284898 540064 284908
rect 539904 284728 540064 284738
rect 538864 284498 538884 284568
rect 538954 284498 539104 284568
rect 539174 284498 539194 284568
rect 538864 283308 539194 284498
rect 540390 284420 540790 286056
rect 541769 285982 541999 286502
rect 542989 286742 543199 287262
rect 543079 286662 543109 286742
rect 542389 286442 542509 286452
rect 542389 286332 542509 286342
rect 542989 286142 543199 286662
rect 544219 286932 544309 286962
rect 543599 286452 543719 286462
rect 543599 286342 543719 286352
rect 544219 286332 544309 286852
rect 544219 286242 544309 286252
rect 543079 286062 543109 286142
rect 542989 286052 543199 286062
rect 557700 286200 557900 286210
rect 557700 285990 557900 286000
rect 558100 286200 558300 286210
rect 558100 285990 558300 286000
rect 558500 286200 558700 286210
rect 558500 285990 558700 286000
rect 558900 286200 559100 286210
rect 558900 285990 559100 286000
rect 559300 286200 559500 286210
rect 559300 285990 559500 286000
rect 541859 285902 541909 285982
rect 541769 285892 541999 285902
rect 557700 285800 557900 285810
rect 557700 285590 557900 285600
rect 558100 285800 558300 285810
rect 558100 285590 558300 285600
rect 558500 285800 558700 285810
rect 558500 285590 558700 285600
rect 558900 285800 559100 285810
rect 558900 285590 559100 285600
rect 559300 285800 559500 285810
rect 559300 285590 559500 285600
rect 541124 285478 541284 285488
rect 541124 285308 541284 285318
rect 542604 285478 542764 285488
rect 542604 285308 542764 285318
rect 543604 285478 543764 285488
rect 543604 285308 543764 285318
rect 557700 285400 557900 285410
rect 557700 285190 557900 285200
rect 558100 285400 558300 285410
rect 558100 285190 558300 285200
rect 558500 285400 558700 285410
rect 558500 285190 558700 285200
rect 558900 285400 559100 285410
rect 558900 285190 559100 285200
rect 559300 285400 559500 285410
rect 559300 285190 559500 285200
rect 542044 285158 542394 285168
rect 542044 285088 542064 285158
rect 542134 285088 542304 285158
rect 542374 285088 542394 285158
rect 541124 284898 541284 284908
rect 541124 284728 541284 284738
rect 542044 284568 542394 285088
rect 557700 285000 557900 285010
rect 542604 284898 542764 284908
rect 542604 284728 542764 284738
rect 543604 284898 543764 284908
rect 557700 284790 557900 284800
rect 558100 285000 558300 285010
rect 558100 284790 558300 284800
rect 558500 285000 558700 285010
rect 558500 284790 558700 284800
rect 558900 285000 559100 285010
rect 558900 284790 559100 284800
rect 559300 285000 559500 285010
rect 559300 284790 559500 284800
rect 543604 284728 543764 284738
rect 542044 284498 542064 284568
rect 542134 284498 542304 284568
rect 542374 284498 542394 284568
rect 540024 284408 540244 284418
rect 540024 284338 540044 284408
rect 540114 284338 540154 284408
rect 540224 284338 540244 284408
rect 540024 283838 540244 284338
rect 540390 284360 540440 284420
rect 540500 284360 540540 284420
rect 540600 284360 540640 284420
rect 540700 284360 540790 284420
rect 540390 284320 540790 284360
rect 540390 284260 540440 284320
rect 540500 284260 540540 284320
rect 540600 284260 540640 284320
rect 540700 284260 540790 284320
rect 540390 284220 540790 284260
rect 540390 284160 540440 284220
rect 540500 284160 540540 284220
rect 540600 284160 540640 284220
rect 540700 284160 540790 284220
rect 540390 284120 540790 284160
rect 540390 284060 540440 284120
rect 540500 284060 540540 284120
rect 540600 284060 540640 284120
rect 540700 284060 540790 284120
rect 540390 283926 540790 284060
rect 540390 283866 540410 283926
rect 540470 283866 540510 283926
rect 540570 283866 540610 283926
rect 540670 283866 540710 283926
rect 540770 283866 540790 283926
rect 540390 283846 540790 283866
rect 540964 284408 541184 284428
rect 540964 284338 540984 284408
rect 541054 284338 541094 284408
rect 541164 284338 541184 284408
rect 540964 283848 541184 284338
rect 540024 283768 540044 283838
rect 540114 283768 540154 283838
rect 540224 283768 540244 283838
rect 539764 283518 539984 283528
rect 539764 283358 539984 283368
rect 538864 283238 538884 283308
rect 538954 283238 539094 283308
rect 539164 283238 539194 283308
rect 538864 283218 539194 283238
rect 538864 283148 538884 283218
rect 538954 283148 539094 283218
rect 539164 283148 539194 283218
rect 537404 282958 537584 282968
rect 537404 282818 537584 282828
rect 538544 282958 538724 282968
rect 538544 282818 538724 282828
rect 538864 282788 539194 283148
rect 540024 283088 540244 283768
rect 540964 283778 540984 283848
rect 541054 283778 541094 283848
rect 541164 283778 541184 283848
rect 540284 283518 540504 283528
rect 540284 283358 540504 283368
rect 540704 283518 540924 283528
rect 540704 283358 540924 283368
rect 540024 283018 540044 283088
rect 540114 283018 540154 283088
rect 540224 283018 540244 283088
rect 539524 282968 539704 282978
rect 539524 282828 539704 282838
rect 538864 282718 538884 282788
rect 538954 282718 539104 282788
rect 539174 282718 539194 282788
rect 538864 282708 539194 282718
rect 540024 282638 540244 283018
rect 540964 283088 541184 283778
rect 541254 283518 541474 283528
rect 541254 283358 541474 283368
rect 540964 283018 540984 283088
rect 541054 283018 541094 283088
rect 541164 283018 541184 283088
rect 540294 282968 540474 282978
rect 540294 282828 540474 282838
rect 540734 282968 540914 282978
rect 540734 282828 540914 282838
rect 540024 282568 540044 282638
rect 540114 282568 540154 282638
rect 540224 282568 540244 282638
rect 540024 282498 540244 282568
rect 540964 282638 541184 283018
rect 542044 283328 542394 284498
rect 557700 284600 557900 284610
rect 557700 284390 557900 284400
rect 558100 284600 558300 284610
rect 558100 284390 558300 284400
rect 558500 284600 558700 284610
rect 558500 284390 558700 284400
rect 558900 284600 559100 284610
rect 558900 284390 559100 284400
rect 559300 284600 559500 284610
rect 559300 284390 559500 284400
rect 557700 284200 557900 284210
rect 557700 283990 557900 284000
rect 558100 284200 558300 284210
rect 558100 283990 558300 284000
rect 558500 284200 558700 284210
rect 558500 283990 558700 284000
rect 558900 284200 559100 284210
rect 558900 283990 559100 284000
rect 559300 284200 559500 284210
rect 559300 283990 559500 284000
rect 557700 283800 557900 283810
rect 557700 283590 557900 283600
rect 558100 283800 558300 283810
rect 558100 283590 558300 283600
rect 558500 283800 558700 283810
rect 558500 283590 558700 283600
rect 558900 283800 559100 283810
rect 558900 283590 559100 283600
rect 559300 283800 559500 283810
rect 559300 283590 559500 283600
rect 542044 283258 542064 283328
rect 542134 283258 542304 283328
rect 542374 283258 542394 283328
rect 542044 283238 542394 283258
rect 542044 283168 542064 283238
rect 542134 283168 542304 283238
rect 542374 283168 542394 283238
rect 557700 283400 557900 283410
rect 557700 283190 557900 283200
rect 558100 283400 558300 283410
rect 558100 283190 558300 283200
rect 558500 283400 558700 283410
rect 558500 283190 558700 283200
rect 558900 283400 559100 283410
rect 558900 283190 559100 283200
rect 559300 283400 559500 283410
rect 559300 283190 559500 283200
rect 541454 282958 541634 282968
rect 541454 282818 541634 282828
rect 542044 282788 542394 283168
rect 557700 283000 557900 283010
rect 542524 282968 542704 282978
rect 542524 282828 542704 282838
rect 543524 282968 543704 282978
rect 543524 282828 543704 282838
rect 557700 282790 557900 282800
rect 558100 283000 558300 283010
rect 558100 282790 558300 282800
rect 558500 283000 558700 283010
rect 558500 282790 558700 282800
rect 558900 283000 559100 283010
rect 558900 282790 559100 282800
rect 559300 283000 559500 283010
rect 559300 282790 559500 282800
rect 542044 282718 542064 282788
rect 542134 282718 542304 282788
rect 542374 282718 542394 282788
rect 542044 282688 542394 282718
rect 540964 282568 540984 282638
rect 541054 282568 541094 282638
rect 541164 282568 541184 282638
rect 540964 282508 541184 282568
rect 557700 282600 557900 282610
rect 557700 282390 557900 282400
rect 558100 282600 558300 282610
rect 558100 282390 558300 282400
rect 558500 282600 558700 282610
rect 558500 282390 558700 282400
rect 558900 282600 559100 282610
rect 558900 282390 559100 282400
rect 559300 282600 559500 282610
rect 559300 282390 559500 282400
rect 567900 281300 568100 281310
rect 572760 281224 572770 281284
rect 572830 281224 572840 281284
rect 572900 281224 572910 281284
rect 572970 281224 572980 281284
rect 573075 281224 573085 281284
rect 573145 281224 573155 281284
rect 573265 281224 573275 281284
rect 573335 281224 573345 281284
rect 573425 281224 573435 281284
rect 573495 281224 573505 281284
rect 573615 281224 573625 281284
rect 573685 281224 573695 281284
rect 573815 281224 573825 281284
rect 573885 281224 573895 281284
rect 573995 281224 574005 281284
rect 574065 281224 574075 281284
rect 574185 281224 574195 281284
rect 574255 281224 574265 281284
rect 574385 281224 574395 281284
rect 574455 281224 574465 281284
rect 574550 281214 574560 281274
rect 574620 281214 574630 281274
rect 567900 281090 568100 281100
rect 537364 281058 537484 281068
rect 537364 280928 537484 280938
rect 543734 281058 543854 281068
rect 572760 281024 572770 281084
rect 572830 281024 572840 281084
rect 572900 281024 572910 281084
rect 572970 281024 572980 281084
rect 573075 281024 573085 281084
rect 573145 281024 573155 281084
rect 573265 281024 573275 281084
rect 573335 281024 573345 281084
rect 573425 281024 573435 281084
rect 573495 281024 573505 281084
rect 573615 281024 573625 281084
rect 573685 281024 573695 281084
rect 573815 281024 573825 281084
rect 573885 281024 573895 281084
rect 573995 281024 574005 281084
rect 574065 281024 574075 281084
rect 574185 281024 574195 281084
rect 574255 281024 574265 281084
rect 574385 281024 574395 281084
rect 574455 281024 574465 281084
rect 574550 281024 574560 281084
rect 574620 281024 574630 281084
rect 543734 280928 543854 280938
rect 567900 281000 568100 281010
rect 572760 280824 572770 280884
rect 572830 280824 572840 280884
rect 572900 280824 572910 280884
rect 572970 280824 572980 280884
rect 573075 280824 573085 280884
rect 573145 280824 573155 280884
rect 573265 280824 573275 280884
rect 573335 280824 573345 280884
rect 573425 280824 573435 280884
rect 573495 280824 573505 280884
rect 573615 280824 573625 280884
rect 573685 280824 573695 280884
rect 573815 280824 573825 280884
rect 573885 280824 573895 280884
rect 573995 280824 574005 280884
rect 574065 280824 574075 280884
rect 574185 280824 574195 280884
rect 574255 280824 574265 280884
rect 574385 280824 574395 280884
rect 574455 280824 574465 280884
rect 574550 280824 574560 280884
rect 574620 280824 574630 280884
rect 567900 280790 568100 280800
rect 567900 280700 568100 280710
rect 13060 280500 13280 280520
rect 13060 280430 13190 280500
rect 13260 280430 13280 280500
rect 572760 280634 572770 280694
rect 572830 280634 572840 280694
rect 572900 280634 572910 280694
rect 572970 280634 572980 280694
rect 573075 280634 573085 280694
rect 573145 280634 573155 280694
rect 573265 280634 573275 280694
rect 573335 280634 573345 280694
rect 573425 280634 573435 280694
rect 573495 280634 573505 280694
rect 573615 280634 573625 280694
rect 573685 280634 573695 280694
rect 573815 280634 573825 280694
rect 573885 280634 573895 280694
rect 573995 280634 574005 280694
rect 574065 280634 574075 280694
rect 574185 280634 574195 280694
rect 574255 280634 574265 280694
rect 574385 280634 574395 280694
rect 574455 280634 574465 280694
rect 574550 280634 574560 280694
rect 574620 280634 574630 280694
rect 567900 280490 568100 280500
rect 572760 280434 572770 280494
rect 572830 280434 572840 280494
rect 572900 280434 572910 280494
rect 572970 280434 572980 280494
rect 573075 280434 573085 280494
rect 573145 280434 573155 280494
rect 573265 280434 573275 280494
rect 573335 280434 573345 280494
rect 573425 280434 573435 280494
rect 573495 280434 573505 280494
rect 573615 280434 573625 280494
rect 573685 280434 573695 280494
rect 573815 280434 573825 280494
rect 573885 280434 573895 280494
rect 573995 280434 574005 280494
rect 574065 280434 574075 280494
rect 574185 280434 574195 280494
rect 574255 280434 574265 280494
rect 574385 280434 574395 280494
rect 574455 280434 574465 280494
rect 574550 280434 574560 280494
rect 574620 280434 574630 280494
rect 13060 280390 13280 280430
rect 13060 280320 13080 280390
rect 13150 280320 13280 280390
rect 13060 280300 13280 280320
rect 567900 280400 568100 280410
rect 572760 280234 572770 280294
rect 572830 280234 572840 280294
rect 572900 280234 572910 280294
rect 572970 280234 572980 280294
rect 573075 280234 573085 280294
rect 573145 280234 573155 280294
rect 573265 280234 573275 280294
rect 573335 280234 573345 280294
rect 573425 280234 573435 280294
rect 573495 280234 573505 280294
rect 573615 280234 573625 280294
rect 573685 280234 573695 280294
rect 573815 280234 573825 280294
rect 573885 280234 573895 280294
rect 573995 280234 574005 280294
rect 574065 280234 574075 280294
rect 574185 280234 574195 280294
rect 574255 280234 574265 280294
rect 574385 280234 574395 280294
rect 574455 280234 574465 280294
rect 574550 280234 574560 280294
rect 574620 280234 574630 280294
rect 567900 280190 568100 280200
rect 14530 278370 14540 278550
rect 14640 278370 14650 278550
rect 14530 277950 14540 278130
rect 14640 277950 14650 278130
rect 537364 278058 537484 278068
rect 537364 277928 537484 277938
rect 543734 278058 543854 278068
rect 543734 277928 543854 277938
rect 30980 276140 45120 276160
rect 30980 275900 31020 276140
rect 31260 275900 32740 276140
rect 32980 275900 34460 276140
rect 34700 275900 35940 276140
rect 36180 275900 37660 276140
rect 37900 275900 39260 276140
rect 39500 275900 40980 276140
rect 41220 275900 42580 276140
rect 42820 275900 44300 276140
rect 44540 275900 44780 276140
rect 45020 275900 45120 276140
rect 30980 275880 45120 275900
rect 12830 275780 12840 275850
rect 12910 275780 12920 275850
rect 13070 275780 13080 275850
rect 13150 275780 13160 275850
rect 13440 275700 20920 275730
rect 13440 275630 13450 275700
rect 13520 275630 13690 275700
rect 13760 275630 14060 275700
rect 14130 275630 20670 275700
rect 20740 275630 20830 275700
rect 20900 275630 20920 275700
rect 13440 275600 20920 275630
rect 12830 275470 12840 275540
rect 12910 275470 12920 275540
rect 13070 275470 13080 275540
rect 13150 275470 13160 275540
rect 13440 275310 13450 275380
rect 13520 275310 13530 275380
rect 13680 275310 13690 275380
rect 13760 275310 13770 275380
rect 12830 275150 12840 275220
rect 12910 275150 12920 275220
rect 13070 275150 13080 275220
rect 13150 275150 13160 275220
rect 17690 275200 17700 275300
rect 17800 275200 17810 275300
rect 17990 275200 18000 275300
rect 18200 275200 18210 275300
rect 18390 275200 18400 275300
rect 18500 275200 18510 275300
rect 13440 274990 13450 275060
rect 13520 274990 13530 275060
rect 13680 274990 13690 275060
rect 13760 274990 13770 275060
rect 537364 275058 537484 275068
rect 20390 275020 27120 275040
rect 20390 274910 20510 275020
rect 20620 274910 21620 275020
rect 21730 274910 22030 275020
rect 22140 274910 23140 275020
rect 23250 274940 24880 275020
rect 24960 274980 27120 275020
rect 24960 274940 26960 274980
rect 23250 274910 26960 274940
rect 20390 274900 26960 274910
rect 27040 274900 27120 274980
rect 537364 274928 537484 274938
rect 543734 275058 543854 275068
rect 543734 274928 543854 274938
rect 12830 274830 12840 274900
rect 12910 274830 12920 274900
rect 13070 274830 13080 274900
rect 13150 274830 13160 274900
rect 20390 274880 27120 274900
rect 20390 274800 24880 274880
rect 24960 274860 27120 274880
rect 24960 274800 26960 274860
rect 20390 274780 26960 274800
rect 27040 274780 27120 274860
rect 20390 274770 27120 274780
rect 13440 274680 13450 274750
rect 13520 274680 13530 274750
rect 13680 274680 13690 274750
rect 13760 274680 13770 274750
rect 13840 274740 17990 274760
rect 13840 274720 17630 274740
rect 13840 274640 13860 274720
rect 13940 274640 15160 274720
rect 15240 274640 15340 274720
rect 15420 274640 17630 274720
rect 13840 274620 17630 274640
rect 17750 274620 17850 274740
rect 17970 274620 17990 274740
rect 20390 274660 20510 274770
rect 20620 274660 21620 274770
rect 21730 274660 22030 274770
rect 22140 274660 23140 274770
rect 23250 274740 27120 274770
rect 23250 274660 24880 274740
rect 24960 274660 26960 274740
rect 27040 274660 27120 274740
rect 20390 274640 27120 274660
rect 13840 274600 17990 274620
rect 12830 274520 12840 274590
rect 12910 274520 12920 274590
rect 13070 274520 13080 274590
rect 13150 274520 13160 274590
rect 18170 274500 22440 274520
rect 13440 274360 13450 274430
rect 13520 274360 13530 274430
rect 13680 274360 13690 274430
rect 13760 274360 13770 274430
rect 18170 274380 18190 274500
rect 18310 274380 18410 274500
rect 18530 274380 19150 274500
rect 19270 274380 19370 274500
rect 19490 274490 22440 274500
rect 19490 274420 22180 274490
rect 22250 274420 22360 274490
rect 22430 274420 22440 274490
rect 19490 274380 22440 274420
rect 18170 274360 22440 274380
rect 15140 274280 15150 274350
rect 15220 274280 15230 274350
rect 15350 274280 15360 274350
rect 15430 274280 15440 274350
rect 16680 274280 16690 274350
rect 16760 274280 16770 274350
rect 16890 274280 16900 274350
rect 16970 274280 16980 274350
rect 12830 274200 12840 274270
rect 12910 274200 12920 274270
rect 13070 274200 13080 274270
rect 13150 274200 13160 274270
rect 14500 274120 14510 274190
rect 14580 274120 14590 274190
rect 14710 274120 14720 274190
rect 14790 274120 14800 274190
rect 16050 274120 16060 274190
rect 16130 274120 16140 274190
rect 16260 274120 16270 274190
rect 16340 274120 16350 274190
rect 20650 274170 20660 274240
rect 20730 274170 20740 274240
rect 20830 274170 20840 274240
rect 20910 274170 20920 274240
rect 22840 274160 22850 274230
rect 22920 274160 22930 274230
rect 23020 274160 23030 274230
rect 23100 274160 23110 274230
rect 13440 274040 13450 274110
rect 13520 274040 13530 274110
rect 13680 274040 13690 274110
rect 13760 274040 13770 274110
rect 15140 273970 15150 274040
rect 15220 273970 15230 274040
rect 15350 273970 15360 274040
rect 15430 273970 15440 274040
rect 16680 274030 20070 274060
rect 16680 273960 16690 274030
rect 16760 273960 16900 274030
rect 16970 273960 19720 274030
rect 19790 273960 19970 274030
rect 20040 273960 20070 274030
rect 12830 273890 12840 273960
rect 12910 273890 12920 273960
rect 13070 273890 13080 273960
rect 13150 273890 13160 273960
rect 16680 273930 20070 273960
rect 21320 273910 21330 273980
rect 21400 273910 21410 273980
rect 21500 273910 21510 273980
rect 21580 273910 21590 273980
rect 22170 273910 22180 273980
rect 22250 273910 22260 273980
rect 22350 273910 22360 273980
rect 22430 273910 22440 273980
rect 14500 273810 14510 273880
rect 14580 273810 14590 273880
rect 14710 273810 14720 273880
rect 14790 273810 14800 273880
rect 16050 273810 16060 273880
rect 16130 273810 16140 273880
rect 16260 273810 16270 273880
rect 16340 273810 16350 273880
rect 13440 273730 13450 273800
rect 13520 273730 13530 273800
rect 13680 273730 13690 273800
rect 13760 273730 13770 273800
rect 15140 273650 15150 273720
rect 15220 273650 15230 273720
rect 15350 273650 15360 273720
rect 15430 273650 15440 273720
rect 16680 273650 16690 273720
rect 16760 273650 16770 273720
rect 16890 273650 16900 273720
rect 16970 273650 16980 273720
rect 20650 273650 20660 273720
rect 20730 273650 20740 273720
rect 20830 273650 20840 273720
rect 20910 273650 20920 273720
rect 22840 273650 22850 273720
rect 22920 273650 22930 273720
rect 23020 273650 23030 273720
rect 23100 273650 23110 273720
rect 12830 273570 12840 273640
rect 12910 273570 12920 273640
rect 13070 273570 13080 273640
rect 13150 273570 13160 273640
rect 26070 273590 26080 273670
rect 26160 273590 26170 273670
rect 26210 273590 26220 273670
rect 26300 273590 26310 273670
rect 14500 273490 14510 273560
rect 14580 273490 14590 273560
rect 14710 273490 14720 273560
rect 14790 273490 14800 273560
rect 13440 273410 13450 273480
rect 13520 273410 13530 273480
rect 13680 273410 13690 273480
rect 13760 273410 13770 273480
rect 15140 273330 15150 273400
rect 15220 273330 15230 273400
rect 15350 273330 15360 273400
rect 15430 273330 15440 273400
rect 12350 273060 12360 273330
rect 12630 273060 12640 273330
rect 12830 273250 12840 273320
rect 12910 273250 12920 273320
rect 13070 273250 13080 273320
rect 13150 273250 13160 273320
rect 13440 273100 13450 273170
rect 13520 273100 13530 273170
rect 13680 273100 13690 273170
rect 13760 273100 13770 273170
rect 13990 273060 14000 273330
rect 14270 273060 14280 273330
rect 15600 273280 15610 273540
rect 15870 273280 15880 273540
rect 16050 273490 16060 273560
rect 16130 273490 16140 273560
rect 16260 273490 16270 273560
rect 16340 273490 16350 273560
rect 16680 273330 16690 273400
rect 16760 273330 16770 273400
rect 16890 273330 16900 273400
rect 16970 273330 16980 273400
rect 21320 273390 21330 273460
rect 21400 273390 21410 273460
rect 21500 273390 21510 273460
rect 21580 273390 21590 273460
rect 22170 273390 22180 273460
rect 22250 273390 22260 273460
rect 22350 273390 22360 273460
rect 22430 273390 22440 273460
rect 24390 273390 24400 273470
rect 24480 273390 24490 273470
rect 25220 273380 25640 273400
rect 25850 273390 25860 273470
rect 25940 273390 25950 273470
rect 26720 273460 29380 273480
rect 25220 273310 25230 273380
rect 25300 273310 25560 273380
rect 25630 273310 25640 273380
rect 26720 273360 26730 273460
rect 26830 273440 29380 273460
rect 26830 273380 29310 273440
rect 29370 273380 29380 273440
rect 26830 273360 29380 273380
rect 26720 273340 29380 273360
rect 25220 273290 25640 273310
rect 14500 273180 14510 273250
rect 14580 273180 14590 273250
rect 14710 273180 14720 273250
rect 14790 273180 14800 273250
rect 16050 273170 16060 273240
rect 16130 273170 16140 273240
rect 16260 273170 16270 273240
rect 16340 273170 16350 273240
rect 18170 273170 18180 273240
rect 18250 273170 18260 273240
rect 18460 273170 18470 273240
rect 18540 273170 18550 273240
rect 19690 273170 19700 273240
rect 19770 273170 19780 273240
rect 19980 273170 19990 273240
rect 20060 273170 20070 273240
rect 24870 273210 28260 273220
rect 20650 273130 20660 273200
rect 20730 273130 20740 273200
rect 20830 273130 20840 273200
rect 20910 273130 20920 273200
rect 22840 273130 22850 273200
rect 22920 273130 22930 273200
rect 23020 273130 23030 273200
rect 23100 273130 23110 273200
rect 24870 273130 24880 273210
rect 24960 273130 28170 273210
rect 28250 273130 28260 273210
rect 24870 273120 28260 273130
rect 28360 273100 28370 273190
rect 28460 273100 28470 273190
rect 29710 273180 30890 273200
rect 29710 273120 29720 273180
rect 29780 273120 30490 273180
rect 30550 273120 30610 273180
rect 30670 273120 30730 273180
rect 30790 273120 30890 273180
rect 29710 273100 30890 273120
rect 15140 273020 15150 273090
rect 15220 273020 15230 273090
rect 15350 273020 15360 273090
rect 15430 273020 15440 273090
rect 16680 273020 16690 273090
rect 16760 273020 16770 273090
rect 16890 273020 16900 273090
rect 16970 273020 16980 273090
rect 17610 273010 17620 273080
rect 17690 273010 17700 273080
rect 17900 273010 17910 273080
rect 17980 273010 17990 273080
rect 19130 273010 19140 273080
rect 19210 273010 19220 273080
rect 19420 273010 19430 273080
rect 19500 273010 19510 273080
rect 28570 273050 29010 273060
rect 12830 272940 12840 273010
rect 12910 272940 12920 273010
rect 13070 272940 13080 273010
rect 13150 272940 13160 273010
rect 14500 272860 14510 272930
rect 14580 272860 14590 272930
rect 14710 272860 14720 272930
rect 14790 272860 14800 272930
rect 16050 272860 16060 272930
rect 16130 272860 16140 272930
rect 16260 272860 16270 272930
rect 16340 272860 16350 272930
rect 18170 272850 18180 272920
rect 18250 272850 18260 272920
rect 18460 272850 18470 272920
rect 18540 272850 18550 272920
rect 19690 272850 19700 272920
rect 19770 272850 19780 272920
rect 19980 272850 19990 272920
rect 20060 272850 20070 272920
rect 21320 272880 21330 272950
rect 21400 272880 21410 272950
rect 21500 272880 21510 272950
rect 21580 272880 21590 272950
rect 22170 272870 22180 272940
rect 22250 272870 22260 272940
rect 22350 272870 22360 272940
rect 22430 272870 22440 272940
rect 24390 272870 24400 272950
rect 24480 272870 24490 272950
rect 25850 272870 25860 272950
rect 25940 272870 25950 272950
rect 27460 272890 27470 273010
rect 27590 272890 27600 273010
rect 28570 272990 28580 273050
rect 28640 272990 28940 273050
rect 29000 272990 29010 273050
rect 28570 272980 29010 272990
rect 29300 272860 29310 272920
rect 29370 272860 29380 272920
rect 13440 272780 13450 272850
rect 13520 272780 13530 272850
rect 13680 272780 13690 272850
rect 13760 272780 13770 272850
rect 15140 272700 15150 272770
rect 15220 272700 15230 272770
rect 15350 272700 15360 272770
rect 15430 272700 15440 272770
rect 16680 272700 16690 272770
rect 16760 272700 16770 272770
rect 16890 272700 16900 272770
rect 16970 272700 16980 272770
rect 17610 272690 17620 272760
rect 17690 272690 17700 272760
rect 17900 272690 17910 272760
rect 17980 272690 17990 272760
rect 12830 272620 12840 272690
rect 12910 272620 12920 272690
rect 13070 272620 13080 272690
rect 13150 272620 13160 272690
rect 14500 272540 14510 272610
rect 14580 272540 14590 272610
rect 14710 272540 14720 272610
rect 14790 272540 14800 272610
rect 16050 272540 16060 272610
rect 16130 272540 16140 272610
rect 16260 272540 16270 272610
rect 16340 272540 16350 272610
rect 18170 272530 18180 272600
rect 18250 272530 18260 272600
rect 18460 272530 18470 272600
rect 18540 272530 18550 272600
rect 13440 272460 13450 272530
rect 13520 272460 13530 272530
rect 13680 272460 13690 272530
rect 13760 272460 13770 272530
rect 18700 272520 18710 272780
rect 18970 272520 18980 272780
rect 19130 272690 19140 272760
rect 19210 272690 19220 272760
rect 19420 272690 19430 272760
rect 19500 272690 19510 272760
rect 19690 272530 19700 272600
rect 19770 272530 19780 272600
rect 19980 272530 19990 272600
rect 20060 272530 20070 272600
rect 20220 272520 20230 272780
rect 20490 272520 20500 272780
rect 20650 272620 20660 272690
rect 20730 272620 20740 272690
rect 20830 272620 20840 272690
rect 20910 272620 20920 272690
rect 21740 272530 21750 272780
rect 22000 272530 22010 272780
rect 22840 272620 22850 272690
rect 22920 272620 22930 272690
rect 23020 272620 23030 272690
rect 23100 272620 23110 272690
rect 23270 272530 23280 272780
rect 23530 272530 23540 272780
rect 25220 272690 25640 272710
rect 24870 272610 24880 272690
rect 24960 272610 24970 272690
rect 25220 272620 25230 272690
rect 25300 272620 25560 272690
rect 25630 272620 25640 272690
rect 25220 272600 25640 272620
rect 26720 272670 27250 272680
rect 26720 272600 26730 272670
rect 26800 272600 27170 272670
rect 27240 272600 27250 272670
rect 26720 272590 27250 272600
rect 27630 272670 28210 272680
rect 27630 272600 27640 272670
rect 27710 272600 28170 272670
rect 28240 272600 28250 272670
rect 27630 272590 28210 272600
rect 28360 272590 28370 272680
rect 28460 272590 28470 272680
rect 28740 272580 28750 272670
rect 28840 272580 28850 272670
rect 29710 272610 29720 272670
rect 29780 272610 29790 272670
rect 30180 272580 30190 272670
rect 30280 272580 30290 272670
rect 15140 272390 15150 272460
rect 15220 272390 15230 272460
rect 15350 272390 15360 272460
rect 15430 272390 15440 272460
rect 16680 272380 16690 272450
rect 16760 272380 16770 272450
rect 16890 272380 16900 272450
rect 16970 272380 16980 272450
rect 17610 272380 17620 272450
rect 17690 272380 17700 272450
rect 17900 272380 17910 272450
rect 17980 272380 17990 272450
rect 19130 272380 19140 272450
rect 19210 272380 19220 272450
rect 19420 272380 19430 272450
rect 19500 272380 19510 272450
rect 12830 272310 12840 272380
rect 12910 272310 12920 272380
rect 13070 272310 13080 272380
rect 13150 272310 13160 272380
rect 21320 272360 21330 272430
rect 21400 272360 21410 272430
rect 21500 272360 21510 272430
rect 21580 272360 21590 272430
rect 22170 272360 22180 272430
rect 22250 272360 22260 272430
rect 22350 272360 22360 272430
rect 22430 272360 22440 272430
rect 24390 272350 24400 272430
rect 24480 272350 24490 272430
rect 25850 272350 25860 272430
rect 25940 272350 25950 272430
rect 12350 272010 12360 272280
rect 12630 272010 12640 272280
rect 13440 272150 13450 272220
rect 13520 272150 13530 272220
rect 13680 272150 13690 272220
rect 13760 272150 13770 272220
rect 12830 271990 12840 272060
rect 12910 271990 12920 272060
rect 13070 271990 13080 272060
rect 13150 271990 13160 272060
rect 13990 272010 14000 272280
rect 14270 272010 14280 272280
rect 14500 272230 14510 272300
rect 14580 272230 14590 272300
rect 14710 272230 14720 272300
rect 14790 272230 14800 272300
rect 16050 272230 16060 272300
rect 16130 272230 16140 272300
rect 16260 272230 16270 272300
rect 16340 272230 16350 272300
rect 18170 272220 18180 272290
rect 18250 272220 18260 272290
rect 18460 272220 18470 272290
rect 18540 272220 18550 272290
rect 19690 272220 19700 272290
rect 19770 272220 19780 272290
rect 19980 272220 19990 272290
rect 20060 272220 20070 272290
rect 27470 272270 27480 272390
rect 27600 272270 27610 272390
rect 29300 272350 29310 272410
rect 29370 272350 29380 272410
rect 28570 272280 29010 272290
rect 28570 272220 28580 272280
rect 28640 272220 28940 272280
rect 29000 272220 29010 272280
rect 28570 272210 29010 272220
rect 24870 272170 28260 272180
rect 15140 272070 15150 272140
rect 15220 272070 15230 272140
rect 15350 272070 15360 272140
rect 15430 272070 15440 272140
rect 16680 272070 16690 272140
rect 16760 272070 16770 272140
rect 16890 272070 16900 272140
rect 16970 272070 16980 272140
rect 17610 272060 17620 272130
rect 17690 272060 17700 272130
rect 17900 272060 17910 272130
rect 17980 272060 17990 272130
rect 19130 272060 19140 272130
rect 19210 272060 19220 272130
rect 19420 272060 19430 272130
rect 19500 272060 19510 272130
rect 20650 272100 20660 272170
rect 20730 272100 20740 272170
rect 20830 272100 20840 272170
rect 20910 272100 20920 272170
rect 22840 272100 22850 272170
rect 22920 272100 22930 272170
rect 23020 272100 23030 272170
rect 23100 272100 23110 272170
rect 24870 272090 24880 272170
rect 24960 272090 28170 272170
rect 28250 272090 28260 272170
rect 24870 272080 28260 272090
rect 28360 272070 28370 272160
rect 28460 272070 28470 272160
rect 29710 272150 30890 272170
rect 29710 272090 29720 272150
rect 29780 272090 30490 272150
rect 30550 272090 30610 272150
rect 30670 272090 30730 272150
rect 30790 272090 30890 272150
rect 29710 272070 30890 272090
rect 537364 272058 537484 272068
rect 14500 271910 14510 271980
rect 14580 271910 14590 271980
rect 14710 271910 14720 271980
rect 14790 271910 14800 271980
rect 13440 271830 13450 271900
rect 13520 271830 13530 271900
rect 13680 271830 13690 271900
rect 13760 271830 13770 271900
rect 15140 271750 15150 271820
rect 15220 271750 15230 271820
rect 15350 271750 15360 271820
rect 15430 271750 15440 271820
rect 15600 271780 15610 272040
rect 15870 271780 15880 272040
rect 25220 271990 25640 272010
rect 16050 271910 16060 271980
rect 16130 271910 16140 271980
rect 16260 271910 16270 271980
rect 16340 271910 16350 271980
rect 25220 271920 25230 271990
rect 25300 271920 25560 271990
rect 25630 271920 25640 271990
rect 21320 271840 21330 271910
rect 21400 271840 21410 271910
rect 21500 271840 21510 271910
rect 21580 271840 21590 271910
rect 22170 271840 22180 271910
rect 22250 271840 22260 271910
rect 22350 271840 22360 271910
rect 22430 271840 22440 271910
rect 24390 271840 24400 271920
rect 24480 271840 24490 271920
rect 25220 271900 25640 271920
rect 25850 271840 25860 271920
rect 25940 271840 25950 271920
rect 26720 271910 29380 271930
rect 537364 271928 537484 271938
rect 543734 272058 543854 272068
rect 543734 271928 543854 271938
rect 16680 271750 16690 271820
rect 16760 271750 16770 271820
rect 16890 271750 16900 271820
rect 16970 271750 16980 271820
rect 26720 271810 26730 271910
rect 26830 271890 29380 271910
rect 26830 271830 29310 271890
rect 29370 271830 29380 271890
rect 26830 271810 29380 271830
rect 26720 271790 29380 271810
rect 12830 271670 12840 271740
rect 12910 271670 12920 271740
rect 13070 271670 13080 271740
rect 13150 271670 13160 271740
rect 14500 271590 14510 271660
rect 14580 271590 14590 271660
rect 14710 271590 14720 271660
rect 14790 271590 14800 271660
rect 16050 271590 16060 271660
rect 16130 271590 16140 271660
rect 16260 271590 16270 271660
rect 16340 271590 16350 271660
rect 20650 271590 20660 271660
rect 20730 271590 20740 271660
rect 20830 271590 20840 271660
rect 20910 271590 20920 271660
rect 22840 271580 22850 271650
rect 22920 271580 22930 271650
rect 23020 271580 23030 271650
rect 23100 271580 23110 271650
rect 26070 271630 26080 271710
rect 26160 271630 26170 271710
rect 26210 271630 26220 271710
rect 26300 271630 26310 271710
rect 13440 271510 13450 271580
rect 13520 271510 13530 271580
rect 13680 271510 13690 271580
rect 13760 271510 13770 271580
rect 16680 271510 20070 271540
rect 15140 271440 15150 271510
rect 15220 271440 15230 271510
rect 15350 271440 15360 271510
rect 15430 271440 15440 271510
rect 16680 271440 16690 271510
rect 16760 271440 16900 271510
rect 16970 271440 19720 271510
rect 19790 271440 19970 271510
rect 20040 271440 20070 271510
rect 12830 271360 12840 271430
rect 12910 271360 12920 271430
rect 13070 271360 13080 271430
rect 13150 271360 13160 271430
rect 16680 271410 20070 271440
rect 14500 271280 14510 271350
rect 14580 271280 14590 271350
rect 14710 271280 14720 271350
rect 14790 271280 14800 271350
rect 16050 271280 16060 271350
rect 16130 271280 16140 271350
rect 16260 271280 16270 271350
rect 16340 271280 16350 271350
rect 21320 271330 21330 271400
rect 21400 271330 21410 271400
rect 21500 271330 21510 271400
rect 21580 271330 21590 271400
rect 22170 271330 22180 271400
rect 22250 271330 22260 271400
rect 22350 271330 22360 271400
rect 22430 271330 22440 271400
rect 13440 271200 13450 271270
rect 13520 271200 13530 271270
rect 13680 271200 13690 271270
rect 13760 271200 13770 271270
rect 15140 271120 15150 271190
rect 15220 271120 15230 271190
rect 15350 271120 15360 271190
rect 15430 271120 15440 271190
rect 16680 271120 16690 271190
rect 16760 271120 16770 271190
rect 16890 271120 16900 271190
rect 16970 271120 16980 271190
rect 12830 271040 12840 271110
rect 12910 271040 12920 271110
rect 13070 271040 13080 271110
rect 13150 271040 13160 271110
rect 20650 271070 20660 271140
rect 20730 271070 20740 271140
rect 20830 271070 20840 271140
rect 20910 271070 20920 271140
rect 22840 271070 22850 271140
rect 22920 271070 22930 271140
rect 23020 271070 23030 271140
rect 23100 271070 23110 271140
rect 14500 270960 14510 271030
rect 14580 270960 14590 271030
rect 14710 270960 14720 271030
rect 14790 270960 14800 271030
rect 16050 270960 16060 271030
rect 16130 270960 16140 271030
rect 16260 270960 16270 271030
rect 16340 270960 16350 271030
rect 13440 270880 13450 270950
rect 13520 270880 13530 270950
rect 13680 270880 13690 270950
rect 13760 270880 13770 270950
rect 18170 270920 22440 270940
rect 18170 270800 18190 270920
rect 18310 270800 18410 270920
rect 18530 270800 19150 270920
rect 19270 270800 19370 270920
rect 19490 270880 22440 270920
rect 19490 270810 22180 270880
rect 22250 270810 22360 270880
rect 22430 270810 22440 270880
rect 19490 270800 22440 270810
rect 12830 270720 12840 270790
rect 12910 270720 12920 270790
rect 13070 270720 13080 270790
rect 13150 270720 13160 270790
rect 18170 270780 22440 270800
rect 13840 270680 17990 270700
rect 13840 270660 17630 270680
rect 13440 270570 13450 270640
rect 13520 270570 13530 270640
rect 13680 270570 13690 270640
rect 13760 270570 13770 270640
rect 13840 270580 13860 270660
rect 13940 270580 15160 270660
rect 15240 270580 15340 270660
rect 15420 270580 17630 270660
rect 13840 270560 17630 270580
rect 17750 270560 17850 270680
rect 17970 270560 17990 270680
rect 13840 270540 17990 270560
rect 20390 270620 24980 270640
rect 20390 270510 20510 270620
rect 20620 270510 21620 270620
rect 21730 270510 22030 270620
rect 22140 270510 23140 270620
rect 23250 270540 24880 270620
rect 24960 270540 24980 270620
rect 23250 270510 24980 270540
rect 20390 270480 24980 270510
rect 12830 270410 12840 270480
rect 12910 270410 12920 270480
rect 13070 270410 13080 270480
rect 13150 270410 13160 270480
rect 20390 270400 24880 270480
rect 24960 270400 24980 270480
rect 20390 270370 24980 270400
rect 13440 270250 13450 270320
rect 13520 270250 13530 270320
rect 13680 270250 13690 270320
rect 13760 270250 13770 270320
rect 20390 270260 20510 270370
rect 20620 270260 21620 270370
rect 21730 270260 22030 270370
rect 22140 270260 23140 270370
rect 23250 270340 24980 270370
rect 23250 270260 24880 270340
rect 24960 270260 24980 270340
rect 20390 270240 24980 270260
rect 12830 270090 12840 270160
rect 12910 270090 12920 270160
rect 13070 270090 13080 270160
rect 13150 270090 13160 270160
rect 19290 270000 19300 270100
rect 19400 270000 19410 270100
rect 19490 270000 19500 270100
rect 19700 270000 19710 270100
rect 19790 270000 19800 270100
rect 19900 270000 19910 270100
rect 13440 269930 13450 270000
rect 13520 269930 13530 270000
rect 13680 269930 13690 270000
rect 13760 269930 13770 270000
rect 12830 269780 12840 269850
rect 12910 269780 12920 269850
rect 13070 269780 13080 269850
rect 13150 269780 13160 269850
rect 13440 269690 20920 269720
rect 13440 269620 13450 269690
rect 13520 269620 13690 269690
rect 13760 269620 14060 269690
rect 14130 269620 20670 269690
rect 20740 269620 20830 269690
rect 20900 269620 20920 269690
rect 13440 269590 20920 269620
rect 12830 269460 12840 269530
rect 12910 269460 12920 269530
rect 13070 269460 13080 269530
rect 13150 269460 13160 269530
rect 30980 269440 45120 269460
rect 30980 269200 31020 269440
rect 31260 269200 32740 269440
rect 32980 269200 34460 269440
rect 34700 269200 35940 269440
rect 36180 269200 37660 269440
rect 37900 269200 39260 269440
rect 39500 269200 40980 269440
rect 41220 269200 42580 269440
rect 42820 269200 44300 269440
rect 44540 269200 44780 269440
rect 45020 269200 45120 269440
rect 30980 269180 45120 269200
rect 537364 269058 537484 269068
rect 537364 268928 537484 268938
rect 543734 269058 543854 269068
rect 543734 268928 543854 268938
rect 44690 268300 44700 268600
rect 45000 268300 45010 268600
rect 44690 267800 44700 268100
rect 45000 267800 45010 268100
rect 542294 267738 543464 267748
rect 537744 267728 538914 267738
rect 44690 267300 44700 267600
rect 45000 267300 45010 267600
rect 537744 267308 538914 267318
rect 539254 267728 540424 267738
rect 539254 267308 540424 267318
rect 540774 267728 541944 267738
rect 542294 267318 543464 267328
rect 540774 267308 541944 267318
rect 14530 267120 14540 267300
rect 14640 267120 14650 267300
rect 14530 266700 14540 266880
rect 14640 266700 14650 266880
rect 44690 266800 44700 267100
rect 45000 266800 45010 267100
rect 44690 266300 44700 266600
rect 45000 266300 45010 266600
rect 44690 265800 44700 266100
rect 45000 265800 45010 266100
rect 44690 265300 44700 265600
rect 45000 265300 45010 265600
rect 13060 265000 13280 265020
rect 13060 264930 13080 265000
rect 13150 264930 13280 265000
rect 13060 264890 13280 264930
rect 13060 264820 13190 264890
rect 13260 264820 13280 264890
rect 13060 264800 13280 264820
rect 44690 264800 44700 265100
rect 45000 264800 45010 265100
rect 44690 264300 44700 264600
rect 45000 264300 45010 264600
rect 44690 263800 44700 264100
rect 45000 263800 45010 264100
rect 44690 263300 44700 263600
rect 45000 263300 45010 263600
rect 44690 262800 44700 263100
rect 45000 262800 45010 263100
rect 44690 262300 44700 262600
rect 45000 262300 45010 262600
rect 44690 261800 44700 262100
rect 45000 261800 45010 262100
rect 44690 261300 44700 261600
rect 45000 261300 45010 261600
rect 44690 260800 44700 261100
rect 45000 260800 45010 261100
rect 14970 252460 14980 252580
rect 15100 252460 15110 252580
rect 15150 252460 15160 252580
rect 15280 252460 15290 252580
rect 15330 252460 15340 252580
rect 15460 252460 15470 252580
rect 15510 252460 15520 252580
rect 15640 252460 15650 252580
rect 15690 252460 15700 252580
rect 15820 252460 15830 252580
rect 9670 252320 9680 252380
rect 9740 252320 9750 252380
rect 9835 252320 9845 252380
rect 9905 252320 9915 252380
rect 10035 252320 10045 252380
rect 10105 252320 10115 252380
rect 10225 252320 10235 252380
rect 10295 252320 10305 252380
rect 10405 252320 10415 252380
rect 10475 252320 10485 252380
rect 10605 252320 10615 252380
rect 10675 252320 10685 252380
rect 10795 252320 10805 252380
rect 10865 252320 10875 252380
rect 10955 252320 10965 252380
rect 11025 252320 11035 252380
rect 11145 252320 11155 252380
rect 11215 252320 11225 252380
rect 11320 252320 11330 252380
rect 11390 252320 11400 252380
rect 11460 252320 11470 252380
rect 11530 252320 11540 252380
rect 5810 252200 5820 252320
rect 5940 252200 5950 252320
rect 9670 252120 9680 252180
rect 9740 252120 9750 252180
rect 9835 252120 9845 252180
rect 9905 252120 9915 252180
rect 10035 252120 10045 252180
rect 10105 252120 10115 252180
rect 10225 252120 10235 252180
rect 10295 252120 10305 252180
rect 10405 252120 10415 252180
rect 10475 252120 10485 252180
rect 10605 252120 10615 252180
rect 10675 252120 10685 252180
rect 10795 252120 10805 252180
rect 10865 252120 10875 252180
rect 10955 252120 10965 252180
rect 11025 252120 11035 252180
rect 11145 252120 11155 252180
rect 11215 252120 11225 252180
rect 11320 252120 11330 252180
rect 11390 252120 11400 252180
rect 11460 252120 11470 252180
rect 11530 252120 11540 252180
rect 5810 252000 5820 252120
rect 5940 252000 5950 252120
rect 9670 251920 9680 251980
rect 9740 251920 9750 251980
rect 9835 251920 9845 251980
rect 9905 251920 9915 251980
rect 10035 251920 10045 251980
rect 10105 251920 10115 251980
rect 10225 251920 10235 251980
rect 10295 251920 10305 251980
rect 10405 251920 10415 251980
rect 10475 251920 10485 251980
rect 10605 251920 10615 251980
rect 10675 251920 10685 251980
rect 10795 251920 10805 251980
rect 10865 251920 10875 251980
rect 10955 251920 10965 251980
rect 11025 251920 11035 251980
rect 11145 251920 11155 251980
rect 11215 251920 11225 251980
rect 11320 251920 11330 251980
rect 11390 251920 11400 251980
rect 11460 251920 11470 251980
rect 11530 251920 11540 251980
rect 5810 251800 5820 251920
rect 5940 251800 5950 251920
rect 9670 251730 9680 251790
rect 9740 251730 9750 251790
rect 9835 251730 9845 251790
rect 9905 251730 9915 251790
rect 10035 251730 10045 251790
rect 10105 251730 10115 251790
rect 10225 251730 10235 251790
rect 10295 251730 10305 251790
rect 10405 251730 10415 251790
rect 10475 251730 10485 251790
rect 10605 251730 10615 251790
rect 10675 251730 10685 251790
rect 10795 251730 10805 251790
rect 10865 251730 10875 251790
rect 10955 251730 10965 251790
rect 11025 251730 11035 251790
rect 11145 251730 11155 251790
rect 11215 251730 11225 251790
rect 11320 251730 11330 251790
rect 11390 251730 11400 251790
rect 11460 251730 11470 251790
rect 11530 251730 11540 251790
rect 5810 251600 5820 251720
rect 5940 251600 5950 251720
rect 9670 251530 9680 251590
rect 9740 251530 9750 251590
rect 9835 251530 9845 251590
rect 9905 251530 9915 251590
rect 10035 251530 10045 251590
rect 10105 251530 10115 251590
rect 10225 251530 10235 251590
rect 10295 251530 10305 251590
rect 10405 251530 10415 251590
rect 10475 251530 10485 251590
rect 10605 251530 10615 251590
rect 10675 251530 10685 251590
rect 10795 251530 10805 251590
rect 10865 251530 10875 251590
rect 10955 251530 10965 251590
rect 11025 251530 11035 251590
rect 11145 251530 11155 251590
rect 11215 251530 11225 251590
rect 11320 251530 11330 251590
rect 11390 251530 11400 251590
rect 11460 251530 11470 251590
rect 11530 251530 11540 251590
rect 5810 251400 5820 251520
rect 5940 251400 5950 251520
rect 9670 251340 9680 251400
rect 9740 251340 9750 251400
rect 9835 251330 9845 251390
rect 9905 251330 9915 251390
rect 10035 251330 10045 251390
rect 10105 251330 10115 251390
rect 10225 251330 10235 251390
rect 10295 251330 10305 251390
rect 10405 251330 10415 251390
rect 10475 251330 10485 251390
rect 10605 251330 10615 251390
rect 10675 251330 10685 251390
rect 10795 251330 10805 251390
rect 10865 251330 10875 251390
rect 10955 251330 10965 251390
rect 11025 251330 11035 251390
rect 11145 251330 11155 251390
rect 11215 251330 11225 251390
rect 11320 251330 11330 251390
rect 11390 251330 11400 251390
rect 11460 251330 11470 251390
rect 11530 251330 11540 251390
rect 9670 241920 9680 241980
rect 9740 241920 9750 241980
rect 9835 241920 9845 241980
rect 9905 241920 9915 241980
rect 10035 241920 10045 241980
rect 10105 241920 10115 241980
rect 10225 241920 10235 241980
rect 10295 241920 10305 241980
rect 10405 241920 10415 241980
rect 10475 241920 10485 241980
rect 10605 241920 10615 241980
rect 10675 241920 10685 241980
rect 10795 241920 10805 241980
rect 10865 241920 10875 241980
rect 10955 241920 10965 241980
rect 11025 241920 11035 241980
rect 11145 241920 11155 241980
rect 11215 241920 11225 241980
rect 11320 241920 11330 241980
rect 11390 241920 11400 241980
rect 11460 241920 11470 241980
rect 11530 241920 11540 241980
rect 16090 241800 16100 242000
rect 16300 241800 16310 242000
rect 9670 241720 9680 241780
rect 9740 241720 9750 241780
rect 9835 241720 9845 241780
rect 9905 241720 9915 241780
rect 10035 241720 10045 241780
rect 10105 241720 10115 241780
rect 10225 241720 10235 241780
rect 10295 241720 10305 241780
rect 10405 241720 10415 241780
rect 10475 241720 10485 241780
rect 10605 241720 10615 241780
rect 10675 241720 10685 241780
rect 10795 241720 10805 241780
rect 10865 241720 10875 241780
rect 10955 241720 10965 241780
rect 11025 241720 11035 241780
rect 11145 241720 11155 241780
rect 11215 241720 11225 241780
rect 11320 241720 11330 241780
rect 11390 241720 11400 241780
rect 11460 241720 11470 241780
rect 11530 241720 11540 241780
rect 9670 241520 9680 241580
rect 9740 241520 9750 241580
rect 9835 241520 9845 241580
rect 9905 241520 9915 241580
rect 10035 241520 10045 241580
rect 10105 241520 10115 241580
rect 10225 241520 10235 241580
rect 10295 241520 10305 241580
rect 10405 241520 10415 241580
rect 10475 241520 10485 241580
rect 10605 241520 10615 241580
rect 10675 241520 10685 241580
rect 10795 241520 10805 241580
rect 10865 241520 10875 241580
rect 10955 241520 10965 241580
rect 11025 241520 11035 241580
rect 11145 241520 11155 241580
rect 11215 241520 11225 241580
rect 11320 241520 11330 241580
rect 11390 241520 11400 241580
rect 11460 241520 11470 241580
rect 11530 241520 11540 241580
rect 16090 241500 16100 241700
rect 16300 241500 16310 241700
rect 9670 241330 9680 241390
rect 9740 241330 9750 241390
rect 9835 241330 9845 241390
rect 9905 241330 9915 241390
rect 10035 241330 10045 241390
rect 10105 241330 10115 241390
rect 10225 241330 10235 241390
rect 10295 241330 10305 241390
rect 10405 241330 10415 241390
rect 10475 241330 10485 241390
rect 10605 241330 10615 241390
rect 10675 241330 10685 241390
rect 10795 241330 10805 241390
rect 10865 241330 10875 241390
rect 10955 241330 10965 241390
rect 11025 241330 11035 241390
rect 11145 241330 11155 241390
rect 11215 241330 11225 241390
rect 11320 241330 11330 241390
rect 11390 241330 11400 241390
rect 11460 241330 11470 241390
rect 11530 241330 11540 241390
rect 16090 241200 16100 241400
rect 16300 241200 16310 241400
rect 9670 241130 9680 241190
rect 9740 241130 9750 241190
rect 9835 241130 9845 241190
rect 9905 241130 9915 241190
rect 10035 241130 10045 241190
rect 10105 241130 10115 241190
rect 10225 241130 10235 241190
rect 10295 241130 10305 241190
rect 10405 241130 10415 241190
rect 10475 241130 10485 241190
rect 10605 241130 10615 241190
rect 10675 241130 10685 241190
rect 10795 241130 10805 241190
rect 10865 241130 10875 241190
rect 10955 241130 10965 241190
rect 11025 241130 11035 241190
rect 11145 241130 11155 241190
rect 11215 241130 11225 241190
rect 11320 241130 11330 241190
rect 11390 241130 11400 241190
rect 11460 241130 11470 241190
rect 11530 241130 11540 241190
rect 9670 240940 9680 241000
rect 9740 240940 9750 241000
rect 9835 240930 9845 240990
rect 9905 240930 9915 240990
rect 10035 240930 10045 240990
rect 10105 240930 10115 240990
rect 10225 240930 10235 240990
rect 10295 240930 10305 240990
rect 10405 240930 10415 240990
rect 10475 240930 10485 240990
rect 10605 240930 10615 240990
rect 10675 240930 10685 240990
rect 10795 240930 10805 240990
rect 10865 240930 10875 240990
rect 10955 240930 10965 240990
rect 11025 240930 11035 240990
rect 11145 240930 11155 240990
rect 11215 240930 11225 240990
rect 11320 240930 11330 240990
rect 11390 240930 11400 240990
rect 11460 240930 11470 240990
rect 11530 240930 11540 240990
rect 16090 240900 16100 241100
rect 16300 240900 16310 241100
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 23400 702060 23520 702180
rect 23600 702060 23720 702180
rect 23800 702060 23920 702180
rect 24000 702060 24120 702180
rect 24200 702060 24320 702180
rect 65060 702080 65240 702260
rect 65400 702080 65580 702260
rect 65740 702080 65920 702260
rect 573280 702140 573380 702240
rect 573420 702140 573520 702240
rect 573560 702140 573660 702240
rect 573700 702140 573800 702240
rect 573840 702140 573940 702240
rect 573980 702140 574080 702240
rect 563840 702020 563940 702120
rect 563980 702020 564080 702120
rect 564120 702020 564220 702120
rect 564260 702020 564360 702120
rect 564400 702020 564500 702120
rect 564540 702020 564640 702120
rect 564680 702020 564780 702120
rect 564820 702020 564920 702120
rect 564960 702020 565060 702120
rect 563840 701880 563940 701980
rect 563980 701880 564080 701980
rect 564120 701880 564220 701980
rect 564260 701880 564360 701980
rect 564400 701880 564500 701980
rect 564540 701880 564640 701980
rect 564680 701880 564780 701980
rect 564820 701880 564920 701980
rect 564960 701880 565060 701980
rect 573280 701880 573380 701980
rect 573420 701880 573520 701980
rect 573560 701880 573660 701980
rect 573700 701880 573800 701980
rect 573840 701880 573940 701980
rect 573980 701880 574080 701980
rect 24460 692900 24580 693020
rect 64720 692860 64860 693000
rect 66060 692860 66200 693000
rect 75120 692860 75260 693000
rect 24460 692720 24580 692840
rect 24460 692540 24580 692660
rect 64720 692660 64860 692800
rect 66060 692660 66200 692800
rect 75120 692660 75260 692800
rect 24460 692360 24580 692480
rect 24460 692180 24580 692300
rect 12900 691700 13100 691900
rect 13200 691700 13400 691900
rect 13500 691700 13700 691900
rect 13800 691700 14000 691900
rect 566300 690900 566500 691100
rect 566700 690900 566900 691100
rect 567100 690900 567300 691100
rect 567500 690900 567700 691100
rect 567900 690900 568100 691100
rect 568300 690900 568500 691100
rect 568700 690900 568900 691100
rect 569100 690900 569300 691100
rect 569500 690900 569700 691100
rect 569900 690900 570100 691100
rect 570300 690900 570500 691100
rect 570700 690900 570900 691100
rect 571100 690900 571300 691100
rect 571500 690900 571700 691100
rect 566300 690500 566500 690700
rect 566700 690500 566900 690700
rect 567100 690500 567300 690700
rect 567500 690500 567700 690700
rect 567900 690500 568100 690700
rect 568300 690500 568500 690700
rect 568700 690500 568900 690700
rect 569100 690500 569300 690700
rect 569500 690500 569700 690700
rect 569900 690500 570100 690700
rect 570300 690500 570500 690700
rect 570700 690500 570900 690700
rect 571100 690500 571300 690700
rect 571500 690500 571700 690700
rect 47200 690200 47300 690300
rect 566300 690100 566500 690300
rect 566700 690100 566900 690300
rect 567100 690100 567300 690300
rect 567500 690100 567700 690300
rect 567900 690100 568100 690300
rect 568300 690100 568500 690300
rect 568700 690100 568900 690300
rect 569100 690100 569300 690300
rect 569500 690100 569700 690300
rect 569900 690100 570100 690300
rect 570300 690100 570500 690300
rect 570700 690100 570900 690300
rect 571100 690100 571300 690300
rect 571500 690100 571700 690300
rect 47200 689800 47300 690000
rect 566300 689700 566500 689900
rect 566700 689700 566900 689900
rect 567100 689700 567300 689900
rect 567500 689700 567700 689900
rect 567900 689700 568100 689900
rect 568300 689700 568500 689900
rect 568700 689700 568900 689900
rect 569100 689700 569300 689900
rect 569500 689700 569700 689900
rect 569900 689700 570100 689900
rect 570300 689700 570500 689900
rect 570700 689700 570900 689900
rect 571100 689700 571300 689900
rect 571500 689700 571700 689900
rect 47200 689500 47300 689600
rect 566300 689300 566500 689500
rect 566700 689300 566900 689500
rect 567100 689300 567300 689500
rect 567500 689300 567700 689500
rect 567900 689300 568100 689500
rect 568300 689300 568500 689500
rect 568700 689300 568900 689500
rect 569100 689300 569300 689500
rect 569500 689300 569700 689500
rect 569900 689300 570100 689500
rect 570300 689300 570500 689500
rect 570700 689300 570900 689500
rect 571100 689300 571300 689500
rect 571500 689300 571700 689500
rect 42000 688600 42100 688700
rect 42000 688300 42100 688500
rect 42000 688100 42100 688200
rect 42260 683040 42340 683120
rect 42400 683040 42480 683120
rect 42540 683040 42620 683120
rect 582360 684520 582440 684600
rect 582540 684520 582620 684600
rect 582360 684360 582440 684440
rect 582540 684360 582620 684440
rect 582360 684200 582440 684280
rect 582540 684200 582620 684280
rect 582360 684020 582440 684100
rect 582540 684020 582620 684100
rect 582360 683860 582440 683940
rect 582540 683860 582620 683940
rect 46660 683040 46740 683120
rect 46800 683040 46880 683120
rect 46940 683040 47020 683120
rect 561700 682000 561900 682200
rect 562100 682000 562300 682200
rect 562500 682000 562700 682200
rect 562900 682000 563100 682200
rect 563300 682000 563500 682200
rect 561700 681600 561900 681800
rect 562100 681600 562300 681800
rect 562500 681600 562700 681800
rect 562900 681600 563100 681800
rect 563300 681600 563500 681800
rect 561700 681200 561900 681400
rect 562100 681200 562300 681400
rect 562500 681200 562700 681400
rect 562900 681200 563100 681400
rect 563300 681200 563500 681400
rect 561700 680800 561900 681000
rect 562100 680800 562300 681000
rect 562500 680800 562700 681000
rect 562900 680800 563100 681000
rect 563300 680800 563500 681000
rect 561700 680400 561900 680600
rect 562100 680400 562300 680600
rect 562500 680400 562700 680600
rect 562900 680400 563100 680600
rect 563300 680400 563500 680600
rect 561700 680000 561900 680200
rect 562100 680000 562300 680200
rect 562500 680000 562700 680200
rect 562900 680000 563100 680200
rect 563300 680000 563500 680200
rect 561700 679600 561900 679800
rect 562100 679600 562300 679800
rect 562500 679600 562700 679800
rect 562900 679600 563100 679800
rect 563300 679600 563500 679800
rect 561700 679200 561900 679400
rect 562100 679200 562300 679400
rect 562500 679200 562700 679400
rect 562900 679200 563100 679400
rect 563300 679200 563500 679400
rect 561700 678800 561900 679000
rect 562100 678800 562300 679000
rect 562500 678800 562700 679000
rect 562900 678800 563100 679000
rect 563300 678800 563500 679000
rect 561700 678400 561900 678600
rect 562100 678400 562300 678600
rect 562500 678400 562700 678600
rect 562900 678400 563100 678600
rect 563300 678400 563500 678600
rect 571900 677100 572100 677300
rect 571900 676800 572100 677000
rect 571900 676500 572100 676700
rect 571900 676200 572100 676400
rect 32800 663000 33100 663300
rect 33300 663000 33600 663300
rect 33800 663000 34100 663300
rect 34300 663000 34600 663300
rect 34800 663000 35100 663300
rect 35300 663000 35600 663300
rect 35800 663000 36100 663300
rect 36300 663000 36600 663300
rect 36800 663000 37100 663300
rect 37300 663000 37600 663300
rect 37800 663000 38100 663300
rect 38300 663000 38600 663300
rect 38800 663000 39100 663300
rect 39300 663000 39600 663300
rect 39800 663000 40100 663300
rect 40300 663000 40600 663300
rect 281080 352580 281140 352640
rect 281180 352580 281240 352640
rect 294760 352600 294820 352660
rect 294860 352600 294920 352660
rect 281080 352480 281140 352540
rect 281180 352480 281240 352540
rect 294760 352500 294820 352560
rect 294860 352500 294920 352560
rect 281060 351020 281120 351080
rect 281160 351020 281220 351080
rect 281060 350920 281120 350980
rect 281160 350920 281220 350980
rect 294760 350860 294820 350920
rect 294860 350860 294920 350920
rect 294760 350760 294820 350820
rect 294860 350760 294920 350820
rect 281060 349320 281120 349380
rect 281160 349320 281220 349380
rect 281060 349220 281120 349280
rect 281160 349220 281220 349280
rect 294760 349160 294820 349220
rect 294860 349160 294920 349220
rect 294760 349060 294820 349120
rect 294860 349060 294920 349120
rect 281040 347620 281100 347680
rect 281140 347620 281200 347680
rect 281040 347520 281100 347580
rect 281140 347520 281200 347580
rect 294760 347460 294820 347520
rect 294860 347460 294920 347520
rect 294760 347360 294820 347420
rect 294860 347360 294920 347420
rect 281060 345920 281120 345980
rect 281160 345920 281220 345980
rect 281060 345820 281120 345880
rect 281160 345820 281220 345880
rect 294760 345760 294820 345820
rect 294860 345760 294920 345820
rect 294760 345660 294820 345720
rect 294860 345660 294920 345720
rect 281060 344200 281120 344260
rect 281160 344200 281220 344260
rect 281060 344100 281120 344160
rect 281160 344100 281220 344160
rect 294800 343900 295100 344200
rect 281040 342500 281100 342560
rect 281140 342500 281200 342560
rect 281040 342400 281100 342460
rect 281140 342400 281200 342460
rect 294760 342360 294820 342420
rect 294860 342360 294920 342420
rect 294760 342260 294820 342320
rect 294860 342260 294920 342320
rect 281060 340660 281120 340720
rect 281160 340660 281220 340720
rect 281060 340560 281120 340620
rect 281160 340560 281220 340620
rect 288300 340500 288600 340800
rect 569280 306140 569380 306240
rect 569420 306140 569520 306240
rect 569560 306140 569660 306240
rect 569700 306140 569800 306240
rect 569840 306140 569940 306240
rect 569980 306140 570080 306240
rect 559840 306020 559940 306120
rect 559980 306020 560080 306120
rect 560120 306020 560220 306120
rect 560260 306020 560360 306120
rect 560400 306020 560500 306120
rect 560540 306020 560640 306120
rect 560680 306020 560780 306120
rect 560820 306020 560920 306120
rect 560960 306020 561060 306120
rect 559840 305880 559940 305980
rect 559980 305880 560080 305980
rect 560120 305880 560220 305980
rect 560260 305880 560360 305980
rect 560400 305880 560500 305980
rect 560540 305880 560640 305980
rect 560680 305880 560780 305980
rect 560820 305880 560920 305980
rect 560960 305880 561060 305980
rect 569280 305880 569380 305980
rect 569420 305880 569520 305980
rect 569560 305880 569660 305980
rect 569700 305880 569800 305980
rect 569840 305880 569940 305980
rect 569980 305880 570080 305980
rect 9680 304320 9740 304380
rect 9845 304320 9905 304380
rect 10045 304320 10105 304380
rect 10235 304320 10295 304380
rect 10415 304320 10475 304380
rect 10615 304320 10675 304380
rect 10805 304320 10865 304380
rect 10965 304320 11025 304380
rect 11155 304320 11215 304380
rect 11330 304320 11390 304380
rect 11470 304320 11530 304380
rect 9680 304120 9740 304180
rect 9845 304120 9905 304180
rect 10045 304120 10105 304180
rect 10235 304120 10295 304180
rect 10415 304120 10475 304180
rect 10615 304120 10675 304180
rect 10805 304120 10865 304180
rect 10965 304120 11025 304180
rect 11155 304120 11215 304180
rect 11330 304120 11390 304180
rect 11470 304120 11530 304180
rect 9680 303920 9740 303980
rect 9845 303920 9905 303980
rect 10045 303920 10105 303980
rect 10235 303920 10295 303980
rect 10415 303920 10475 303980
rect 10615 303920 10675 303980
rect 10805 303920 10865 303980
rect 10965 303920 11025 303980
rect 11155 303920 11215 303980
rect 11330 303920 11390 303980
rect 11470 303920 11530 303980
rect 9680 303730 9740 303790
rect 9845 303730 9905 303790
rect 10045 303730 10105 303790
rect 10235 303730 10295 303790
rect 10415 303730 10475 303790
rect 10615 303730 10675 303790
rect 10805 303730 10865 303790
rect 10965 303730 11025 303790
rect 11155 303730 11215 303790
rect 11330 303730 11390 303790
rect 11470 303730 11530 303790
rect 9680 303530 9740 303590
rect 9845 303530 9905 303590
rect 10045 303530 10105 303590
rect 10235 303530 10295 303590
rect 10415 303530 10475 303590
rect 10615 303530 10675 303590
rect 10805 303530 10865 303590
rect 10965 303530 11025 303590
rect 11155 303530 11215 303590
rect 11330 303530 11390 303590
rect 11470 303530 11530 303590
rect 9680 303340 9740 303400
rect 9845 303330 9905 303390
rect 10045 303330 10105 303390
rect 10235 303330 10295 303390
rect 10415 303330 10475 303390
rect 10615 303330 10675 303390
rect 10805 303330 10865 303390
rect 10965 303330 11025 303390
rect 11155 303330 11215 303390
rect 11330 303330 11390 303390
rect 11470 303330 11530 303390
rect 15000 303120 15140 303260
rect 15200 303120 15340 303260
rect 559940 302060 560000 302120
rect 560130 302060 560190 302120
rect 560330 302060 560390 302120
rect 560520 302060 560580 302120
rect 560720 302060 560780 302120
rect 560920 302060 560980 302120
rect 569140 302060 569200 302120
rect 569330 302060 569390 302120
rect 569530 302060 569590 302120
rect 569720 302060 569780 302120
rect 569920 302060 569980 302120
rect 570120 302060 570180 302120
rect 559930 301895 559990 301955
rect 560130 301895 560190 301955
rect 560330 301895 560390 301955
rect 560520 301895 560580 301955
rect 560720 301895 560780 301955
rect 560920 301895 560980 301955
rect 569130 301895 569190 301955
rect 569330 301895 569390 301955
rect 569530 301895 569590 301955
rect 569720 301895 569780 301955
rect 569920 301895 569980 301955
rect 570120 301895 570180 301955
rect 559930 301695 559990 301755
rect 560130 301695 560190 301755
rect 560330 301695 560390 301755
rect 560520 301695 560580 301755
rect 560720 301695 560780 301755
rect 560920 301695 560980 301755
rect 569130 301695 569190 301755
rect 569330 301695 569390 301755
rect 569530 301695 569590 301755
rect 569720 301695 569780 301755
rect 569920 301695 569980 301755
rect 570120 301695 570180 301755
rect 559930 301505 559990 301565
rect 560130 301505 560190 301565
rect 560330 301505 560390 301565
rect 560520 301505 560580 301565
rect 560720 301505 560780 301565
rect 560920 301505 560980 301565
rect 569130 301505 569190 301565
rect 569330 301505 569390 301565
rect 569530 301505 569590 301565
rect 569720 301505 569780 301565
rect 569920 301505 569980 301565
rect 570120 301505 570180 301565
rect 559930 301325 559990 301385
rect 560130 301325 560190 301385
rect 560330 301325 560390 301385
rect 560520 301325 560580 301385
rect 560720 301325 560780 301385
rect 560920 301325 560980 301385
rect 569130 301325 569190 301385
rect 569330 301325 569390 301385
rect 569530 301325 569590 301385
rect 569720 301325 569780 301385
rect 569920 301325 569980 301385
rect 570120 301325 570180 301385
rect 559930 301125 559990 301185
rect 560130 301125 560190 301185
rect 560330 301125 560390 301185
rect 560520 301125 560580 301185
rect 560720 301125 560780 301185
rect 560920 301125 560980 301185
rect 569130 301125 569190 301185
rect 569330 301125 569390 301185
rect 569530 301125 569590 301185
rect 569720 301125 569780 301185
rect 569920 301125 569980 301185
rect 570120 301125 570180 301185
rect 559930 300935 559990 300995
rect 560130 300935 560190 300995
rect 560330 300935 560390 300995
rect 560520 300935 560580 300995
rect 560720 300935 560780 300995
rect 560920 300935 560980 300995
rect 569130 300935 569190 300995
rect 569330 300935 569390 300995
rect 569530 300935 569590 300995
rect 569720 300935 569780 300995
rect 569920 300935 569980 300995
rect 570120 300935 570180 300995
rect 559930 300775 559990 300835
rect 560130 300775 560190 300835
rect 560330 300775 560390 300835
rect 560520 300775 560580 300835
rect 560720 300775 560780 300835
rect 560920 300775 560980 300835
rect 569130 300775 569190 300835
rect 569330 300775 569390 300835
rect 569530 300775 569590 300835
rect 569720 300775 569780 300835
rect 569920 300775 569980 300835
rect 570120 300775 570180 300835
rect 559930 300585 559990 300645
rect 560130 300585 560190 300645
rect 560330 300585 560390 300645
rect 560520 300585 560580 300645
rect 560720 300585 560780 300645
rect 560920 300585 560980 300645
rect 569130 300585 569190 300645
rect 569330 300585 569390 300645
rect 569530 300585 569590 300645
rect 569720 300585 569780 300645
rect 569920 300585 569980 300645
rect 570120 300585 570180 300645
rect 559930 300410 559990 300470
rect 560130 300410 560190 300470
rect 560330 300410 560390 300470
rect 560520 300410 560580 300470
rect 560720 300410 560780 300470
rect 560920 300410 560980 300470
rect 569130 300410 569190 300470
rect 569330 300410 569390 300470
rect 569530 300410 569590 300470
rect 569720 300410 569780 300470
rect 569920 300410 569980 300470
rect 570120 300410 570180 300470
rect 559930 300270 559990 300330
rect 560130 300270 560190 300330
rect 560330 300270 560390 300330
rect 560520 300270 560580 300330
rect 560720 300270 560780 300330
rect 560920 300270 560980 300330
rect 569130 300270 569190 300330
rect 569330 300270 569390 300330
rect 569530 300270 569590 300330
rect 569720 300270 569780 300330
rect 569920 300270 569980 300330
rect 570120 300270 570180 300330
rect 537969 294892 538059 294962
rect 538139 294892 538229 294962
rect 540459 294892 540549 294962
rect 540629 294892 540719 294962
rect 537089 294602 537169 294682
rect 537239 294602 537319 294682
rect 15000 294060 15140 294200
rect 15200 294060 15340 294200
rect 537089 294062 537169 294142
rect 537239 294062 537319 294142
rect 9680 293920 9740 293980
rect 9845 293920 9905 293980
rect 10045 293920 10105 293980
rect 10235 293920 10295 293980
rect 10415 293920 10475 293980
rect 10615 293920 10675 293980
rect 10805 293920 10865 293980
rect 10965 293920 11025 293980
rect 11155 293920 11215 293980
rect 11330 293920 11390 293980
rect 11470 293920 11530 293980
rect 5740 293740 5920 293920
rect 9680 293720 9740 293780
rect 9845 293720 9905 293780
rect 10045 293720 10105 293780
rect 10235 293720 10295 293780
rect 10415 293720 10475 293780
rect 10615 293720 10675 293780
rect 10805 293720 10865 293780
rect 10965 293720 11025 293780
rect 11155 293720 11215 293780
rect 11330 293720 11390 293780
rect 11470 293720 11530 293780
rect 5740 293400 5920 293580
rect 9680 293520 9740 293580
rect 9845 293520 9905 293580
rect 10045 293520 10105 293580
rect 10235 293520 10295 293580
rect 10415 293520 10475 293580
rect 10615 293520 10675 293580
rect 10805 293520 10865 293580
rect 10965 293520 11025 293580
rect 11155 293520 11215 293580
rect 11330 293520 11390 293580
rect 11470 293520 11530 293580
rect 537979 293842 538069 293912
rect 538119 293842 538209 293912
rect 537089 293522 537169 293602
rect 537239 293522 537319 293602
rect 9680 293330 9740 293390
rect 9845 293330 9905 293390
rect 10045 293330 10105 293390
rect 10235 293330 10295 293390
rect 10415 293330 10475 293390
rect 10615 293330 10675 293390
rect 10805 293330 10865 293390
rect 10965 293330 11025 293390
rect 11155 293330 11215 293390
rect 11330 293330 11390 293390
rect 11470 293330 11530 293390
rect 5740 293060 5920 293240
rect 9680 293130 9740 293190
rect 9845 293130 9905 293190
rect 10045 293130 10105 293190
rect 10235 293130 10295 293190
rect 10415 293130 10475 293190
rect 10615 293130 10675 293190
rect 10805 293130 10865 293190
rect 10965 293130 11025 293190
rect 11155 293130 11215 293190
rect 11330 293130 11390 293190
rect 11470 293130 11530 293190
rect 537979 293302 538059 293382
rect 538149 293302 538229 293382
rect 9680 292940 9740 293000
rect 9845 292930 9905 292990
rect 10045 292930 10105 292990
rect 10235 292930 10295 292990
rect 10415 292930 10475 292990
rect 10615 292930 10675 292990
rect 10805 292930 10865 292990
rect 10965 292930 11025 292990
rect 11155 292930 11215 292990
rect 11330 292930 11390 292990
rect 11470 292930 11530 292990
rect 15000 292720 15140 292860
rect 15200 292720 15340 292860
rect 530629 291992 530759 292132
rect 530879 291992 531009 292132
rect 542919 294892 542999 294972
rect 543089 294892 543169 294972
rect 562300 294900 562500 295100
rect 562700 294900 562900 295100
rect 563100 294900 563300 295100
rect 563500 294900 563700 295100
rect 563900 294900 564100 295100
rect 564300 294900 564500 295100
rect 564700 294900 564900 295100
rect 565100 294900 565300 295100
rect 565500 294900 565700 295100
rect 565900 294900 566100 295100
rect 566300 294900 566500 295100
rect 566700 294900 566900 295100
rect 567100 294900 567300 295100
rect 567500 294900 567700 295100
rect 539579 294602 539659 294682
rect 539729 294602 539809 294682
rect 539579 294062 539659 294142
rect 539729 294062 539809 294142
rect 540459 293842 540549 293912
rect 540619 293852 540709 293922
rect 539579 293522 539659 293602
rect 539729 293522 539809 293602
rect 540459 293302 540539 293382
rect 540629 293302 540709 293382
rect 538379 292922 538459 293002
rect 538489 292922 538569 293002
rect 538379 292312 538459 292392
rect 538489 292312 538569 292392
rect 537979 292142 538069 292222
rect 538139 292142 538229 292222
rect 542059 294602 542139 294682
rect 542209 294602 542289 294682
rect 542059 294062 542139 294142
rect 542209 294062 542289 294142
rect 542069 293522 542149 293602
rect 542209 293522 542289 293602
rect 542919 293852 542999 293922
rect 543089 293852 543169 293922
rect 542919 293302 542999 293382
rect 543089 293302 543169 293382
rect 540789 292922 540869 293002
rect 540899 292922 540979 293002
rect 540789 292332 540869 292412
rect 540899 292332 540979 292412
rect 540459 292142 540539 292212
rect 540629 292142 540709 292212
rect 540789 291752 540869 291832
rect 540899 291752 540979 291832
rect 562300 294500 562500 294700
rect 562700 294500 562900 294700
rect 563100 294500 563300 294700
rect 563500 294500 563700 294700
rect 563900 294500 564100 294700
rect 564300 294500 564500 294700
rect 564700 294500 564900 294700
rect 565100 294500 565300 294700
rect 565500 294500 565700 294700
rect 565900 294500 566100 294700
rect 566300 294500 566500 294700
rect 566700 294500 566900 294700
rect 567100 294500 567300 294700
rect 567500 294500 567700 294700
rect 562300 294100 562500 294300
rect 562700 294100 562900 294300
rect 563100 294100 563300 294300
rect 563500 294100 563700 294300
rect 563900 294100 564100 294300
rect 564300 294100 564500 294300
rect 564700 294100 564900 294300
rect 565100 294100 565300 294300
rect 565500 294100 565700 294300
rect 565900 294100 566100 294300
rect 566300 294100 566500 294300
rect 566700 294100 566900 294300
rect 567100 294100 567300 294300
rect 567500 294100 567700 294300
rect 562300 293700 562500 293900
rect 562700 293700 562900 293900
rect 563100 293700 563300 293900
rect 563500 293700 563700 293900
rect 563900 293700 564100 293900
rect 564300 293700 564500 293900
rect 564700 293700 564900 293900
rect 565100 293700 565300 293900
rect 565500 293700 565700 293900
rect 565900 293700 566100 293900
rect 566300 293700 566500 293900
rect 566700 293700 566900 293900
rect 567100 293700 567300 293900
rect 567500 293700 567700 293900
rect 562300 293300 562500 293500
rect 562700 293300 562900 293500
rect 563100 293300 563300 293500
rect 563500 293300 563700 293500
rect 563900 293300 564100 293500
rect 564300 293300 564500 293500
rect 564700 293300 564900 293500
rect 565100 293300 565300 293500
rect 565500 293300 565700 293500
rect 565900 293300 566100 293500
rect 566300 293300 566500 293500
rect 566700 293300 566900 293500
rect 567100 293300 567300 293500
rect 567500 293300 567700 293500
rect 543249 292912 543329 292992
rect 543359 292912 543439 292992
rect 543249 292332 543329 292412
rect 543359 292332 543439 292412
rect 542919 292142 542999 292212
rect 543089 292142 543169 292212
rect 543249 291752 543329 291832
rect 543359 291752 543439 291832
rect 550129 292162 550259 292302
rect 550389 292162 550519 292302
rect 534869 291542 534959 291652
rect 535029 291542 535119 291652
rect 533080 290880 533140 290940
rect 533180 290880 533240 290940
rect 533280 290880 533340 290940
rect 533080 290760 533140 290820
rect 533180 290760 533240 290820
rect 533280 290760 533340 290820
rect 533080 290660 533140 290720
rect 533180 290660 533240 290720
rect 533280 290660 533340 290720
rect 533080 290520 533140 290580
rect 533180 290520 533240 290580
rect 533280 290520 533340 290580
rect 533080 290420 533140 290480
rect 533180 290420 533240 290480
rect 533280 290420 533340 290480
rect 533080 290320 533140 290380
rect 533180 290320 533240 290380
rect 533280 290320 533340 290380
rect 533080 290220 533140 290280
rect 533180 290220 533240 290280
rect 533280 290220 533340 290280
rect 536119 291062 536209 291142
rect 536299 291062 536389 291142
rect 536119 289982 536209 290062
rect 536299 289992 536389 290072
rect 531759 289122 531849 289252
rect 531969 289122 532059 289252
rect 538649 291062 538739 291142
rect 538809 291062 538899 291142
rect 538649 289982 538739 290062
rect 538809 289982 538899 290062
rect 537089 288292 537169 288372
rect 537239 288292 537319 288372
rect 538379 289052 538459 289132
rect 538489 289052 538569 289132
rect 538279 288662 538389 288772
rect 539139 288662 539249 288772
rect 539579 288312 539659 288392
rect 539729 288312 539809 288392
rect 541119 291062 541209 291142
rect 541279 291062 541369 291142
rect 541119 289982 541209 290062
rect 541279 289982 541369 290062
rect 540789 289052 540869 289132
rect 540899 289052 540979 289132
rect 540349 288662 540459 288772
rect 541199 288662 541309 288772
rect 537569 287562 537679 287652
rect 537509 286352 537629 286452
rect 538729 286352 538849 286452
rect 539939 286352 540059 286452
rect 542059 288312 542139 288392
rect 542199 288312 542279 288392
rect 544799 291522 544879 291602
rect 544969 291522 545049 291602
rect 543569 291062 543659 291142
rect 543729 291062 543819 291142
rect 543569 289982 543659 290062
rect 543729 289982 543819 290062
rect 543249 289062 543329 289142
rect 543359 289062 543439 289142
rect 546069 291062 546159 291142
rect 546229 291062 546319 291142
rect 546069 289982 546159 290062
rect 546229 289982 546319 290062
rect 549069 289152 549139 289242
rect 549229 289152 549299 289242
rect 542769 288662 542879 288772
rect 543649 288662 543759 288772
rect 572750 288704 572810 288764
rect 572890 288704 572950 288764
rect 573065 288704 573125 288764
rect 573255 288704 573315 288764
rect 573415 288704 573475 288764
rect 573605 288704 573665 288764
rect 573805 288704 573865 288764
rect 573985 288704 574045 288764
rect 574175 288704 574235 288764
rect 574375 288704 574435 288764
rect 574540 288694 574600 288754
rect 572750 288504 572810 288564
rect 572890 288504 572950 288564
rect 573065 288504 573125 288564
rect 573255 288504 573315 288564
rect 573415 288504 573475 288564
rect 573605 288504 573665 288564
rect 573805 288504 573865 288564
rect 573985 288504 574045 288564
rect 574175 288504 574235 288564
rect 574375 288504 574435 288564
rect 574540 288504 574600 288564
rect 578360 288520 578440 288600
rect 578540 288520 578620 288600
rect 572750 288304 572810 288364
rect 572890 288304 572950 288364
rect 573065 288304 573125 288364
rect 573255 288304 573315 288364
rect 573415 288304 573475 288364
rect 573605 288304 573665 288364
rect 573805 288304 573865 288364
rect 573985 288304 574045 288364
rect 574175 288304 574235 288364
rect 574375 288304 574435 288364
rect 574540 288304 574600 288364
rect 578360 288360 578440 288440
rect 578540 288360 578620 288440
rect 578360 288200 578440 288280
rect 578540 288200 578620 288280
rect 572750 288114 572810 288174
rect 572890 288114 572950 288174
rect 573065 288114 573125 288174
rect 573255 288114 573315 288174
rect 573415 288114 573475 288174
rect 573605 288114 573665 288174
rect 573805 288114 573865 288174
rect 573985 288114 574045 288174
rect 574175 288114 574235 288174
rect 574375 288114 574435 288174
rect 574540 288114 574600 288174
rect 542479 287562 542589 287652
rect 578360 288020 578440 288100
rect 578540 288020 578620 288100
rect 572750 287914 572810 287974
rect 572890 287914 572950 287974
rect 573065 287914 573125 287974
rect 573255 287914 573315 287974
rect 573415 287914 573475 287974
rect 573605 287914 573665 287974
rect 573805 287914 573865 287974
rect 573985 287914 574045 287974
rect 574175 287914 574235 287974
rect 574375 287914 574435 287974
rect 574540 287914 574600 287974
rect 578360 287860 578440 287940
rect 578540 287860 578620 287940
rect 572750 287714 572810 287774
rect 572890 287714 572950 287774
rect 573065 287714 573125 287774
rect 573255 287714 573315 287774
rect 573415 287714 573475 287774
rect 573605 287714 573665 287774
rect 573805 287714 573865 287774
rect 573985 287714 574045 287774
rect 574175 287714 574235 287774
rect 574375 287714 574435 287774
rect 574540 287714 574600 287774
rect 541159 286352 541279 286452
rect 537384 285318 537544 285478
rect 538444 285318 538604 285478
rect 539904 285318 540064 285478
rect 537384 284738 537544 284898
rect 538444 284738 538604 284898
rect 539904 284738 540064 284898
rect 543599 286352 543719 286452
rect 557700 286000 557900 286200
rect 558100 286000 558300 286200
rect 558500 286000 558700 286200
rect 558900 286000 559100 286200
rect 559300 286000 559500 286200
rect 557700 285600 557900 285800
rect 558100 285600 558300 285800
rect 558500 285600 558700 285800
rect 558900 285600 559100 285800
rect 559300 285600 559500 285800
rect 541124 285318 541284 285478
rect 542604 285318 542764 285478
rect 543604 285318 543764 285478
rect 557700 285200 557900 285400
rect 558100 285200 558300 285400
rect 558500 285200 558700 285400
rect 558900 285200 559100 285400
rect 559300 285200 559500 285400
rect 541124 284738 541284 284898
rect 542604 284738 542764 284898
rect 543604 284738 543764 284898
rect 557700 284800 557900 285000
rect 558100 284800 558300 285000
rect 558500 284800 558700 285000
rect 558900 284800 559100 285000
rect 559300 284800 559500 285000
rect 540440 284360 540500 284420
rect 540540 284360 540600 284420
rect 540640 284360 540700 284420
rect 540440 284260 540500 284320
rect 540540 284260 540600 284320
rect 540640 284260 540700 284320
rect 540440 284160 540500 284220
rect 540540 284160 540600 284220
rect 540640 284160 540700 284220
rect 540440 284060 540500 284120
rect 540540 284060 540600 284120
rect 540640 284060 540700 284120
rect 539764 283368 539984 283518
rect 537404 282828 537584 282958
rect 538544 282828 538724 282958
rect 540284 283368 540504 283518
rect 540704 283368 540924 283518
rect 539524 282838 539704 282968
rect 541254 283368 541474 283518
rect 540294 282838 540474 282968
rect 540734 282838 540914 282968
rect 557700 284400 557900 284600
rect 558100 284400 558300 284600
rect 558500 284400 558700 284600
rect 558900 284400 559100 284600
rect 559300 284400 559500 284600
rect 557700 284000 557900 284200
rect 558100 284000 558300 284200
rect 558500 284000 558700 284200
rect 558900 284000 559100 284200
rect 559300 284000 559500 284200
rect 557700 283600 557900 283800
rect 558100 283600 558300 283800
rect 558500 283600 558700 283800
rect 558900 283600 559100 283800
rect 559300 283600 559500 283800
rect 557700 283200 557900 283400
rect 558100 283200 558300 283400
rect 558500 283200 558700 283400
rect 558900 283200 559100 283400
rect 559300 283200 559500 283400
rect 541454 282828 541634 282958
rect 542524 282838 542704 282968
rect 543524 282838 543704 282968
rect 557700 282800 557900 283000
rect 558100 282800 558300 283000
rect 558500 282800 558700 283000
rect 558900 282800 559100 283000
rect 559300 282800 559500 283000
rect 557700 282400 557900 282600
rect 558100 282400 558300 282600
rect 558500 282400 558700 282600
rect 558900 282400 559100 282600
rect 559300 282400 559500 282600
rect 567900 281100 568100 281300
rect 572770 281224 572830 281284
rect 572910 281224 572970 281284
rect 573085 281224 573145 281284
rect 573275 281224 573335 281284
rect 573435 281224 573495 281284
rect 573625 281224 573685 281284
rect 573825 281224 573885 281284
rect 574005 281224 574065 281284
rect 574195 281224 574255 281284
rect 574395 281224 574455 281284
rect 574560 281214 574620 281274
rect 537364 280938 537484 281058
rect 543734 280938 543854 281058
rect 572770 281024 572830 281084
rect 572910 281024 572970 281084
rect 573085 281024 573145 281084
rect 573275 281024 573335 281084
rect 573435 281024 573495 281084
rect 573625 281024 573685 281084
rect 573825 281024 573885 281084
rect 574005 281024 574065 281084
rect 574195 281024 574255 281084
rect 574395 281024 574455 281084
rect 574560 281024 574620 281084
rect 567900 280800 568100 281000
rect 572770 280824 572830 280884
rect 572910 280824 572970 280884
rect 573085 280824 573145 280884
rect 573275 280824 573335 280884
rect 573435 280824 573495 280884
rect 573625 280824 573685 280884
rect 573825 280824 573885 280884
rect 574005 280824 574065 280884
rect 574195 280824 574255 280884
rect 574395 280824 574455 280884
rect 574560 280824 574620 280884
rect 13190 280430 13260 280500
rect 567900 280500 568100 280700
rect 572770 280634 572830 280694
rect 572910 280634 572970 280694
rect 573085 280634 573145 280694
rect 573275 280634 573335 280694
rect 573435 280634 573495 280694
rect 573625 280634 573685 280694
rect 573825 280634 573885 280694
rect 574005 280634 574065 280694
rect 574195 280634 574255 280694
rect 574395 280634 574455 280694
rect 574560 280634 574620 280694
rect 572770 280434 572830 280494
rect 572910 280434 572970 280494
rect 573085 280434 573145 280494
rect 573275 280434 573335 280494
rect 573435 280434 573495 280494
rect 573625 280434 573685 280494
rect 573825 280434 573885 280494
rect 574005 280434 574065 280494
rect 574195 280434 574255 280494
rect 574395 280434 574455 280494
rect 574560 280434 574620 280494
rect 13080 280320 13150 280390
rect 567900 280200 568100 280400
rect 572770 280234 572830 280294
rect 572910 280234 572970 280294
rect 573085 280234 573145 280294
rect 573275 280234 573335 280294
rect 573435 280234 573495 280294
rect 573625 280234 573685 280294
rect 573825 280234 573885 280294
rect 574005 280234 574065 280294
rect 574195 280234 574255 280294
rect 574395 280234 574455 280294
rect 574560 280234 574620 280294
rect 14540 278370 14640 278550
rect 14540 277950 14640 278130
rect 537364 277938 537484 278058
rect 543734 277938 543854 278058
rect 31020 275900 31260 276140
rect 32740 275900 32980 276140
rect 34460 275900 34700 276140
rect 35940 275900 36180 276140
rect 37660 275900 37900 276140
rect 39260 275900 39500 276140
rect 40980 275900 41220 276140
rect 42580 275900 42820 276140
rect 44300 275900 44540 276140
rect 12840 275780 12910 275850
rect 13080 275780 13150 275850
rect 13450 275630 13520 275700
rect 13690 275630 13760 275700
rect 14060 275630 14130 275700
rect 20670 275630 20740 275700
rect 20830 275630 20900 275700
rect 12840 275470 12910 275540
rect 13080 275470 13150 275540
rect 13450 275310 13520 275380
rect 13690 275310 13760 275380
rect 12840 275150 12910 275220
rect 13080 275150 13150 275220
rect 17700 275200 17800 275300
rect 18000 275200 18200 275300
rect 18400 275200 18500 275300
rect 13450 274990 13520 275060
rect 13690 274990 13760 275060
rect 24880 274940 24960 275020
rect 26960 274900 27040 274980
rect 537364 274938 537484 275058
rect 543734 274938 543854 275058
rect 12840 274830 12910 274900
rect 13080 274830 13150 274900
rect 24880 274800 24960 274880
rect 26960 274780 27040 274860
rect 13450 274680 13520 274750
rect 13690 274680 13760 274750
rect 15160 274640 15240 274720
rect 15340 274640 15420 274720
rect 17630 274620 17750 274740
rect 17850 274620 17970 274740
rect 24880 274660 24960 274740
rect 26960 274660 27040 274740
rect 12840 274520 12910 274590
rect 13080 274520 13150 274590
rect 13450 274360 13520 274430
rect 13690 274360 13760 274430
rect 18190 274380 18310 274500
rect 18410 274380 18530 274500
rect 19150 274380 19270 274500
rect 19370 274380 19490 274500
rect 22180 274420 22250 274490
rect 22360 274420 22430 274490
rect 15150 274280 15220 274350
rect 15360 274280 15430 274350
rect 16690 274280 16760 274350
rect 16900 274280 16970 274350
rect 12840 274200 12910 274270
rect 13080 274200 13150 274270
rect 14510 274120 14580 274190
rect 14720 274120 14790 274190
rect 16060 274120 16130 274190
rect 16270 274120 16340 274190
rect 20660 274170 20730 274240
rect 20840 274170 20910 274240
rect 22850 274160 22920 274230
rect 23030 274160 23100 274230
rect 13450 274040 13520 274110
rect 13690 274040 13760 274110
rect 15150 273970 15220 274040
rect 15360 273970 15430 274040
rect 16690 273960 16760 274030
rect 16900 273960 16970 274030
rect 19720 273960 19790 274030
rect 19970 273960 20040 274030
rect 12840 273890 12910 273960
rect 13080 273890 13150 273960
rect 21330 273910 21400 273980
rect 21510 273910 21580 273980
rect 22180 273910 22250 273980
rect 22360 273910 22430 273980
rect 14510 273810 14580 273880
rect 14720 273810 14790 273880
rect 16060 273810 16130 273880
rect 16270 273810 16340 273880
rect 13450 273730 13520 273800
rect 13690 273730 13760 273800
rect 15150 273650 15220 273720
rect 15360 273650 15430 273720
rect 16690 273650 16760 273720
rect 16900 273650 16970 273720
rect 20660 273650 20730 273720
rect 20840 273650 20910 273720
rect 22850 273650 22920 273720
rect 23030 273650 23100 273720
rect 12840 273570 12910 273640
rect 13080 273570 13150 273640
rect 26080 273590 26160 273670
rect 26220 273590 26300 273670
rect 14510 273490 14580 273560
rect 14720 273490 14790 273560
rect 13450 273410 13520 273480
rect 13690 273410 13760 273480
rect 15150 273330 15220 273400
rect 15360 273330 15430 273400
rect 12360 273060 12630 273330
rect 12840 273250 12910 273320
rect 13080 273250 13150 273320
rect 13450 273100 13520 273170
rect 13690 273100 13760 273170
rect 14000 273060 14270 273330
rect 15610 273280 15870 273540
rect 16060 273490 16130 273560
rect 16270 273490 16340 273560
rect 16690 273330 16760 273400
rect 16900 273330 16970 273400
rect 21330 273390 21400 273460
rect 21510 273390 21580 273460
rect 22180 273390 22250 273460
rect 22360 273390 22430 273460
rect 24400 273390 24480 273470
rect 25860 273390 25940 273470
rect 29310 273380 29370 273440
rect 14510 273180 14580 273250
rect 14720 273180 14790 273250
rect 16060 273170 16130 273240
rect 16270 273170 16340 273240
rect 18180 273170 18250 273240
rect 18470 273170 18540 273240
rect 19700 273170 19770 273240
rect 19990 273170 20060 273240
rect 20660 273130 20730 273200
rect 20840 273130 20910 273200
rect 22850 273130 22920 273200
rect 23030 273130 23100 273200
rect 24880 273130 24960 273210
rect 28370 273100 28460 273190
rect 29720 273120 29780 273180
rect 15150 273020 15220 273090
rect 15360 273020 15430 273090
rect 16690 273020 16760 273090
rect 16900 273020 16970 273090
rect 17620 273010 17690 273080
rect 17910 273010 17980 273080
rect 19140 273010 19210 273080
rect 19430 273010 19500 273080
rect 12840 272940 12910 273010
rect 13080 272940 13150 273010
rect 14510 272860 14580 272930
rect 14720 272860 14790 272930
rect 16060 272860 16130 272930
rect 16270 272860 16340 272930
rect 18180 272850 18250 272920
rect 18470 272850 18540 272920
rect 19700 272850 19770 272920
rect 19990 272850 20060 272920
rect 21330 272880 21400 272950
rect 21510 272880 21580 272950
rect 22180 272870 22250 272940
rect 22360 272870 22430 272940
rect 24400 272870 24480 272950
rect 25860 272870 25940 272950
rect 27470 272890 27590 273010
rect 29310 272860 29370 272920
rect 13450 272780 13520 272850
rect 13690 272780 13760 272850
rect 15150 272700 15220 272770
rect 15360 272700 15430 272770
rect 16690 272700 16760 272770
rect 16900 272700 16970 272770
rect 17620 272690 17690 272760
rect 17910 272690 17980 272760
rect 12840 272620 12910 272690
rect 13080 272620 13150 272690
rect 14510 272540 14580 272610
rect 14720 272540 14790 272610
rect 16060 272540 16130 272610
rect 16270 272540 16340 272610
rect 18180 272530 18250 272600
rect 18470 272530 18540 272600
rect 13450 272460 13520 272530
rect 13690 272460 13760 272530
rect 18710 272520 18970 272780
rect 19140 272690 19210 272760
rect 19430 272690 19500 272760
rect 19700 272530 19770 272600
rect 19990 272530 20060 272600
rect 20230 272520 20490 272780
rect 20660 272620 20730 272690
rect 20840 272620 20910 272690
rect 21750 272530 22000 272780
rect 22850 272620 22920 272690
rect 23030 272620 23100 272690
rect 23280 272530 23530 272780
rect 24880 272610 24960 272690
rect 28370 272590 28460 272680
rect 28750 272580 28840 272670
rect 29720 272610 29780 272670
rect 30190 272580 30280 272670
rect 15150 272390 15220 272460
rect 15360 272390 15430 272460
rect 16690 272380 16760 272450
rect 16900 272380 16970 272450
rect 17620 272380 17690 272450
rect 17910 272380 17980 272450
rect 19140 272380 19210 272450
rect 19430 272380 19500 272450
rect 12840 272310 12910 272380
rect 13080 272310 13150 272380
rect 21330 272360 21400 272430
rect 21510 272360 21580 272430
rect 22180 272360 22250 272430
rect 22360 272360 22430 272430
rect 24400 272350 24480 272430
rect 25860 272350 25940 272430
rect 12360 272010 12630 272280
rect 13450 272150 13520 272220
rect 13690 272150 13760 272220
rect 12840 271990 12910 272060
rect 13080 271990 13150 272060
rect 14000 272010 14270 272280
rect 14510 272230 14580 272300
rect 14720 272230 14790 272300
rect 16060 272230 16130 272300
rect 16270 272230 16340 272300
rect 18180 272220 18250 272290
rect 18470 272220 18540 272290
rect 19700 272220 19770 272290
rect 19990 272220 20060 272290
rect 27480 272270 27600 272390
rect 29310 272350 29370 272410
rect 15150 272070 15220 272140
rect 15360 272070 15430 272140
rect 16690 272070 16760 272140
rect 16900 272070 16970 272140
rect 17620 272060 17690 272130
rect 17910 272060 17980 272130
rect 19140 272060 19210 272130
rect 19430 272060 19500 272130
rect 20660 272100 20730 272170
rect 20840 272100 20910 272170
rect 22850 272100 22920 272170
rect 23030 272100 23100 272170
rect 24880 272090 24960 272170
rect 28370 272070 28460 272160
rect 29720 272090 29780 272150
rect 14510 271910 14580 271980
rect 14720 271910 14790 271980
rect 13450 271830 13520 271900
rect 13690 271830 13760 271900
rect 15150 271750 15220 271820
rect 15360 271750 15430 271820
rect 15610 271780 15870 272040
rect 16060 271910 16130 271980
rect 16270 271910 16340 271980
rect 537364 271938 537484 272058
rect 21330 271840 21400 271910
rect 21510 271840 21580 271910
rect 22180 271840 22250 271910
rect 22360 271840 22430 271910
rect 24400 271840 24480 271920
rect 25860 271840 25940 271920
rect 543734 271938 543854 272058
rect 16690 271750 16760 271820
rect 16900 271750 16970 271820
rect 29310 271830 29370 271890
rect 12840 271670 12910 271740
rect 13080 271670 13150 271740
rect 14510 271590 14580 271660
rect 14720 271590 14790 271660
rect 16060 271590 16130 271660
rect 16270 271590 16340 271660
rect 20660 271590 20730 271660
rect 20840 271590 20910 271660
rect 22850 271580 22920 271650
rect 23030 271580 23100 271650
rect 26080 271630 26160 271710
rect 26220 271630 26300 271710
rect 13450 271510 13520 271580
rect 13690 271510 13760 271580
rect 15150 271440 15220 271510
rect 15360 271440 15430 271510
rect 16690 271440 16760 271510
rect 16900 271440 16970 271510
rect 19720 271440 19790 271510
rect 19970 271440 20040 271510
rect 12840 271360 12910 271430
rect 13080 271360 13150 271430
rect 14510 271280 14580 271350
rect 14720 271280 14790 271350
rect 16060 271280 16130 271350
rect 16270 271280 16340 271350
rect 21330 271330 21400 271400
rect 21510 271330 21580 271400
rect 22180 271330 22250 271400
rect 22360 271330 22430 271400
rect 13450 271200 13520 271270
rect 13690 271200 13760 271270
rect 15150 271120 15220 271190
rect 15360 271120 15430 271190
rect 16690 271120 16760 271190
rect 16900 271120 16970 271190
rect 12840 271040 12910 271110
rect 13080 271040 13150 271110
rect 20660 271070 20730 271140
rect 20840 271070 20910 271140
rect 22850 271070 22920 271140
rect 23030 271070 23100 271140
rect 14510 270960 14580 271030
rect 14720 270960 14790 271030
rect 16060 270960 16130 271030
rect 16270 270960 16340 271030
rect 13450 270880 13520 270950
rect 13690 270880 13760 270950
rect 18190 270800 18310 270920
rect 18410 270800 18530 270920
rect 19150 270800 19270 270920
rect 19370 270800 19490 270920
rect 22180 270810 22250 270880
rect 22360 270810 22430 270880
rect 12840 270720 12910 270790
rect 13080 270720 13150 270790
rect 13450 270570 13520 270640
rect 13690 270570 13760 270640
rect 15160 270580 15240 270660
rect 15340 270580 15420 270660
rect 17630 270560 17750 270680
rect 17850 270560 17970 270680
rect 24880 270540 24960 270620
rect 12840 270410 12910 270480
rect 13080 270410 13150 270480
rect 24880 270400 24960 270480
rect 13450 270250 13520 270320
rect 13690 270250 13760 270320
rect 24880 270260 24960 270340
rect 12840 270090 12910 270160
rect 13080 270090 13150 270160
rect 19300 270000 19400 270100
rect 19500 270000 19700 270100
rect 19800 270000 19900 270100
rect 13450 269930 13520 270000
rect 13690 269930 13760 270000
rect 12840 269780 12910 269850
rect 13080 269780 13150 269850
rect 13450 269620 13520 269690
rect 13690 269620 13760 269690
rect 14060 269620 14130 269690
rect 20670 269620 20740 269690
rect 20830 269620 20900 269690
rect 12840 269460 12910 269530
rect 13080 269460 13150 269530
rect 31020 269200 31260 269440
rect 32740 269200 32980 269440
rect 34460 269200 34700 269440
rect 35940 269200 36180 269440
rect 37660 269200 37900 269440
rect 39260 269200 39500 269440
rect 40980 269200 41220 269440
rect 42580 269200 42820 269440
rect 44300 269200 44540 269440
rect 537364 268938 537484 269058
rect 543734 268938 543854 269058
rect 44700 268300 45000 268600
rect 44700 267800 45000 268100
rect 44700 267300 45000 267600
rect 537744 267318 538914 267728
rect 539254 267318 540424 267728
rect 540774 267318 541944 267728
rect 542294 267328 543464 267738
rect 14540 267120 14640 267300
rect 14540 266700 14640 266880
rect 44700 266800 45000 267100
rect 44700 266300 45000 266600
rect 44700 265800 45000 266100
rect 44700 265300 45000 265600
rect 13080 264930 13150 265000
rect 13190 264820 13260 264890
rect 44700 264800 45000 265100
rect 44700 264300 45000 264600
rect 44700 263800 45000 264100
rect 44700 263300 45000 263600
rect 44700 262800 45000 263100
rect 44700 262300 45000 262600
rect 44700 261800 45000 262100
rect 44700 261300 45000 261600
rect 44700 260800 45000 261100
rect 14980 252460 15100 252580
rect 15160 252460 15280 252580
rect 15340 252460 15460 252580
rect 15520 252460 15640 252580
rect 15700 252460 15820 252580
rect 9680 252320 9740 252380
rect 9845 252320 9905 252380
rect 10045 252320 10105 252380
rect 10235 252320 10295 252380
rect 10415 252320 10475 252380
rect 10615 252320 10675 252380
rect 10805 252320 10865 252380
rect 10965 252320 11025 252380
rect 11155 252320 11215 252380
rect 11330 252320 11390 252380
rect 11470 252320 11530 252380
rect 5820 252200 5940 252320
rect 9680 252120 9740 252180
rect 9845 252120 9905 252180
rect 10045 252120 10105 252180
rect 10235 252120 10295 252180
rect 10415 252120 10475 252180
rect 10615 252120 10675 252180
rect 10805 252120 10865 252180
rect 10965 252120 11025 252180
rect 11155 252120 11215 252180
rect 11330 252120 11390 252180
rect 11470 252120 11530 252180
rect 5820 252000 5940 252120
rect 9680 251920 9740 251980
rect 9845 251920 9905 251980
rect 10045 251920 10105 251980
rect 10235 251920 10295 251980
rect 10415 251920 10475 251980
rect 10615 251920 10675 251980
rect 10805 251920 10865 251980
rect 10965 251920 11025 251980
rect 11155 251920 11215 251980
rect 11330 251920 11390 251980
rect 11470 251920 11530 251980
rect 5820 251800 5940 251920
rect 9680 251730 9740 251790
rect 9845 251730 9905 251790
rect 10045 251730 10105 251790
rect 10235 251730 10295 251790
rect 10415 251730 10475 251790
rect 10615 251730 10675 251790
rect 10805 251730 10865 251790
rect 10965 251730 11025 251790
rect 11155 251730 11215 251790
rect 11330 251730 11390 251790
rect 11470 251730 11530 251790
rect 5820 251600 5940 251720
rect 9680 251530 9740 251590
rect 9845 251530 9905 251590
rect 10045 251530 10105 251590
rect 10235 251530 10295 251590
rect 10415 251530 10475 251590
rect 10615 251530 10675 251590
rect 10805 251530 10865 251590
rect 10965 251530 11025 251590
rect 11155 251530 11215 251590
rect 11330 251530 11390 251590
rect 11470 251530 11530 251590
rect 5820 251400 5940 251520
rect 9680 251340 9740 251400
rect 9845 251330 9905 251390
rect 10045 251330 10105 251390
rect 10235 251330 10295 251390
rect 10415 251330 10475 251390
rect 10615 251330 10675 251390
rect 10805 251330 10865 251390
rect 10965 251330 11025 251390
rect 11155 251330 11215 251390
rect 11330 251330 11390 251390
rect 11470 251330 11530 251390
rect 9680 241920 9740 241980
rect 9845 241920 9905 241980
rect 10045 241920 10105 241980
rect 10235 241920 10295 241980
rect 10415 241920 10475 241980
rect 10615 241920 10675 241980
rect 10805 241920 10865 241980
rect 10965 241920 11025 241980
rect 11155 241920 11215 241980
rect 11330 241920 11390 241980
rect 11470 241920 11530 241980
rect 16100 241800 16300 242000
rect 9680 241720 9740 241780
rect 9845 241720 9905 241780
rect 10045 241720 10105 241780
rect 10235 241720 10295 241780
rect 10415 241720 10475 241780
rect 10615 241720 10675 241780
rect 10805 241720 10865 241780
rect 10965 241720 11025 241780
rect 11155 241720 11215 241780
rect 11330 241720 11390 241780
rect 11470 241720 11530 241780
rect 9680 241520 9740 241580
rect 9845 241520 9905 241580
rect 10045 241520 10105 241580
rect 10235 241520 10295 241580
rect 10415 241520 10475 241580
rect 10615 241520 10675 241580
rect 10805 241520 10865 241580
rect 10965 241520 11025 241580
rect 11155 241520 11215 241580
rect 11330 241520 11390 241580
rect 11470 241520 11530 241580
rect 16100 241500 16300 241700
rect 9680 241330 9740 241390
rect 9845 241330 9905 241390
rect 10045 241330 10105 241390
rect 10235 241330 10295 241390
rect 10415 241330 10475 241390
rect 10615 241330 10675 241390
rect 10805 241330 10865 241390
rect 10965 241330 11025 241390
rect 11155 241330 11215 241390
rect 11330 241330 11390 241390
rect 11470 241330 11530 241390
rect 16100 241200 16300 241400
rect 9680 241130 9740 241190
rect 9845 241130 9905 241190
rect 10045 241130 10105 241190
rect 10235 241130 10295 241190
rect 10415 241130 10475 241190
rect 10615 241130 10675 241190
rect 10805 241130 10865 241190
rect 10965 241130 11025 241190
rect 11155 241130 11215 241190
rect 11330 241130 11390 241190
rect 11470 241130 11530 241190
rect 9680 240940 9740 241000
rect 9845 240930 9905 240990
rect 10045 240930 10105 240990
rect 10235 240930 10295 240990
rect 10415 240930 10475 240990
rect 10615 240930 10675 240990
rect 10805 240930 10865 240990
rect 10965 240930 11025 240990
rect 11155 240930 11215 240990
rect 11330 240930 11390 240990
rect 11470 240930 11530 240990
rect 16100 240900 16300 241100
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 703700 470394 704800
rect 510594 704000 515394 704800
rect 520594 704000 525394 704800
rect 566594 704000 571594 704800
rect 16200 702200 21200 702300
rect 16200 702000 16400 702200
rect 16600 702000 16800 702200
rect 17000 702000 17200 702200
rect 17400 702000 17600 702200
rect 17800 702000 18000 702200
rect 18200 702000 18400 702200
rect 18600 702000 18800 702200
rect 19000 702000 19200 702200
rect 19400 702000 19600 702200
rect 19800 702000 20000 702200
rect 20200 702000 20400 702200
rect 20600 702000 20800 702200
rect 21000 702000 21200 702200
rect 65050 702260 65250 702265
rect 23390 702180 23530 702185
rect 23390 702060 23400 702180
rect 23520 702060 23530 702180
rect 23390 702055 23530 702060
rect 23590 702180 23730 702185
rect 23590 702060 23600 702180
rect 23720 702060 23730 702180
rect 23590 702055 23730 702060
rect 23790 702180 23930 702185
rect 23790 702060 23800 702180
rect 23920 702060 23930 702180
rect 23790 702055 23930 702060
rect 23990 702180 24130 702185
rect 23990 702060 24000 702180
rect 24120 702060 24130 702180
rect 23990 702055 24130 702060
rect 24190 702180 24330 702185
rect 24190 702060 24200 702180
rect 24320 702060 24330 702180
rect 65050 702080 65060 702260
rect 65240 702080 65250 702260
rect 65050 702075 65250 702080
rect 65390 702260 65590 702265
rect 65390 702080 65400 702260
rect 65580 702080 65590 702260
rect 65390 702075 65590 702080
rect 65730 702260 65930 702265
rect 65730 702080 65740 702260
rect 65920 702080 65930 702260
rect 65730 702075 65930 702080
rect 68200 702200 73200 702300
rect 24190 702055 24330 702060
rect 16200 701800 21200 702000
rect 16200 701600 16400 701800
rect 16600 701600 16800 701800
rect 17000 701600 17200 701800
rect 17400 701600 17600 701800
rect 17800 701600 18000 701800
rect 18200 701600 18400 701800
rect 18600 701600 18800 701800
rect 19000 701600 19200 701800
rect 19400 701600 19600 701800
rect 19800 701600 20000 701800
rect 20200 701600 20400 701800
rect 20600 701600 20800 701800
rect 21000 701600 21200 701800
rect 16200 701400 21200 701600
rect 16200 701200 16400 701400
rect 16600 701200 16800 701400
rect 17000 701200 17200 701400
rect 17400 701200 17600 701400
rect 17800 701200 18000 701400
rect 18200 701200 18400 701400
rect 18600 701200 18800 701400
rect 19000 701200 19200 701400
rect 19400 701200 19600 701400
rect 19800 701200 20000 701400
rect 20200 701200 20400 701400
rect 20600 701200 20800 701400
rect 21000 701200 21200 701400
rect 16200 701000 21200 701200
rect 16200 700800 16400 701000
rect 16600 700800 16800 701000
rect 17000 700800 17200 701000
rect 17400 700800 17600 701000
rect 17800 700800 18000 701000
rect 18200 700800 18400 701000
rect 18600 700800 18800 701000
rect 19000 700800 19200 701000
rect 19400 700800 19600 701000
rect 19800 700800 20000 701000
rect 20200 700800 20400 701000
rect 20600 700800 20800 701000
rect 21000 700800 21200 701000
rect 16200 700600 21200 700800
rect 16200 700400 16400 700600
rect 16600 700400 16800 700600
rect 17000 700400 17200 700600
rect 17400 700400 17600 700600
rect 17800 700400 18000 700600
rect 18200 700400 18400 700600
rect 18600 700400 18800 700600
rect 19000 700400 19200 700600
rect 19400 700400 19600 700600
rect 19800 700400 20000 700600
rect 20200 700400 20400 700600
rect 20600 700400 20800 700600
rect 21000 700400 21200 700600
rect 16200 700200 21200 700400
rect 16200 700000 16400 700200
rect 16600 700000 16800 700200
rect 17000 700000 17200 700200
rect 17400 700000 17600 700200
rect 17800 700000 18000 700200
rect 18200 700000 18400 700200
rect 18600 700000 18800 700200
rect 19000 700000 19200 700200
rect 19400 700000 19600 700200
rect 19800 700000 20000 700200
rect 20200 700000 20400 700200
rect 20600 700000 20800 700200
rect 21000 700000 21200 700200
rect 16200 699800 21200 700000
rect 68200 702000 68400 702200
rect 68600 702000 68800 702200
rect 69000 702000 69200 702200
rect 69400 702000 69600 702200
rect 69800 702000 70000 702200
rect 70200 702000 70400 702200
rect 70600 702000 70800 702200
rect 71000 702000 71200 702200
rect 71400 702000 71600 702200
rect 71800 702000 72000 702200
rect 72200 702000 72400 702200
rect 72600 702000 72800 702200
rect 73000 702000 73200 702200
rect 68200 701800 73200 702000
rect 68200 701600 68400 701800
rect 68600 701600 68800 701800
rect 69000 701600 69200 701800
rect 69400 701600 69600 701800
rect 69800 701600 70000 701800
rect 70200 701600 70400 701800
rect 70600 701600 70800 701800
rect 71000 701600 71200 701800
rect 71400 701600 71600 701800
rect 71800 701600 72000 701800
rect 72200 701600 72400 701800
rect 72600 701600 72800 701800
rect 73000 701600 73200 701800
rect 68200 701400 73200 701600
rect 68200 701200 68400 701400
rect 68600 701200 68800 701400
rect 69000 701200 69200 701400
rect 69400 701200 69600 701400
rect 69800 701200 70000 701400
rect 70200 701200 70400 701400
rect 70600 701200 70800 701400
rect 71000 701200 71200 701400
rect 71400 701200 71600 701400
rect 71800 701200 72000 701400
rect 72200 701200 72400 701400
rect 72600 701200 72800 701400
rect 73000 701200 73200 701400
rect 68200 701000 73200 701200
rect 68200 700800 68400 701000
rect 68600 700800 68800 701000
rect 69000 700800 69200 701000
rect 69400 700800 69600 701000
rect 69800 700800 70000 701000
rect 70200 700800 70400 701000
rect 70600 700800 70800 701000
rect 71000 700800 71200 701000
rect 71400 700800 71600 701000
rect 71800 700800 72000 701000
rect 72200 700800 72400 701000
rect 72600 700800 72800 701000
rect 73000 700800 73200 701000
rect 68200 700600 73200 700800
rect 68200 700400 68400 700600
rect 68600 700400 68800 700600
rect 69000 700400 69200 700600
rect 69400 700400 69600 700600
rect 69800 700400 70000 700600
rect 70200 700400 70400 700600
rect 70600 700400 70800 700600
rect 71000 700400 71200 700600
rect 71400 700400 71600 700600
rect 71800 700400 72000 700600
rect 72200 700400 72400 700600
rect 72600 700400 72800 700600
rect 73000 700400 73200 700600
rect 68200 700200 73200 700400
rect 68200 700000 68400 700200
rect 68600 700000 68800 700200
rect 69000 700000 69200 700200
rect 69400 700000 69600 700200
rect 69800 700000 70000 700200
rect 70200 700000 70400 700200
rect 70600 700000 70800 700200
rect 71000 700000 71200 700200
rect 71400 700000 71600 700200
rect 71800 700000 72000 700200
rect 72200 700000 72400 700200
rect 72600 700000 72800 700200
rect 73000 700000 73200 700200
rect 68200 699800 73200 700000
rect 12990 698000 13000 698200
rect 13200 698000 13210 698200
rect 13590 698000 13600 698200
rect 13800 698000 13810 698200
rect 23390 698000 23400 698200
rect 23600 698000 23610 698200
rect 23790 698000 23800 698200
rect 24000 698000 24010 698200
rect 24190 698000 24200 698200
rect 24400 698000 24410 698200
rect 64990 698000 65000 698200
rect 65200 698000 65210 698200
rect 65590 698000 65600 698200
rect 65800 698000 65810 698200
rect 75390 698000 75400 698200
rect 75600 698000 75610 698200
rect 75990 698000 76000 698200
rect 76200 698000 76210 698200
rect 12990 697600 13000 697800
rect 13200 697600 13210 697800
rect 13590 697600 13600 697800
rect 13800 697600 13810 697800
rect 23390 697600 23400 697800
rect 23600 697600 23610 697800
rect 23790 697600 23800 697800
rect 24000 697600 24010 697800
rect 24190 697600 24200 697800
rect 24400 697600 24410 697800
rect 64990 697600 65000 697800
rect 65200 697600 65210 697800
rect 65590 697600 65600 697800
rect 65800 697600 65810 697800
rect 75390 697600 75400 697800
rect 75600 697600 75610 697800
rect 75990 697600 76000 697800
rect 76200 697600 76210 697800
rect 23390 697200 23400 697400
rect 23600 697200 23610 697400
rect 23790 697200 23800 697400
rect 24000 697200 24010 697400
rect 24190 697200 24200 697400
rect 24400 697200 24410 697400
rect 64990 697200 65000 697400
rect 65200 697200 65210 697400
rect 65590 697200 65600 697400
rect 65800 697200 65810 697400
rect 75390 697200 75400 697400
rect 75600 697200 75610 697400
rect 75990 697200 76000 697400
rect 76200 697200 76210 697400
rect 12990 697000 13000 697200
rect 13200 697000 13210 697200
rect 13590 697000 13600 697200
rect 13800 697000 13810 697200
rect 23390 696800 23400 697000
rect 23600 696800 23610 697000
rect 23790 696800 23800 697000
rect 24000 696800 24010 697000
rect 24190 696800 24200 697000
rect 24400 696800 24410 697000
rect 64990 696800 65000 697000
rect 65200 696800 65210 697000
rect 65590 696800 65600 697000
rect 65800 696800 65810 697000
rect 75390 696800 75400 697000
rect 75600 696800 75610 697000
rect 75990 696800 76000 697000
rect 76200 696800 76210 697000
rect 12990 696600 13000 696800
rect 13200 696600 13210 696800
rect 13590 696600 13600 696800
rect 13800 696600 13810 696800
rect 23300 696600 24400 696700
rect 23300 696400 23400 696600
rect 23600 696400 23800 696600
rect 24000 696400 24200 696600
rect 24400 696400 24410 696600
rect 64990 696400 65000 696600
rect 65200 696400 65210 696600
rect 65590 696400 65600 696600
rect 65800 696400 65810 696600
rect 75390 696400 75400 696600
rect 75600 696400 75610 696600
rect 75990 696400 76000 696600
rect 76200 696400 76210 696600
rect 24440 693020 39320 693060
rect 24440 692900 24460 693020
rect 24580 693000 39320 693020
rect 24580 692900 38700 693000
rect 24440 692840 38700 692900
rect 38860 692840 39120 693000
rect 39280 692840 39320 693000
rect 24440 692720 24460 692840
rect 24580 692780 39320 692840
rect 24580 692720 38700 692780
rect 24440 692660 38700 692720
rect 24440 692540 24460 692660
rect 24580 692620 38700 692660
rect 38860 692620 39120 692780
rect 39280 692620 39320 692780
rect 49920 693000 64880 693040
rect 49920 692860 49960 693000
rect 50100 692860 50180 693000
rect 50320 692860 50400 693000
rect 50540 692860 64720 693000
rect 64860 692860 64880 693000
rect 49920 692800 64880 692860
rect 49920 692660 49960 692800
rect 50100 692660 50180 692800
rect 50320 692660 50400 692800
rect 50540 692660 64720 692800
rect 64860 692660 64880 692800
rect 49920 692620 64880 692660
rect 66040 693000 75280 693040
rect 66040 692860 66060 693000
rect 66200 692860 75120 693000
rect 75260 692860 75280 693000
rect 66040 692800 75280 692860
rect 66040 692660 66060 692800
rect 66200 692660 75120 692800
rect 75260 692660 75280 692800
rect 66040 692620 75280 692660
rect 24580 692560 39320 692620
rect 24580 692540 38700 692560
rect 24440 692480 38700 692540
rect 24440 692360 24460 692480
rect 24580 692400 38700 692480
rect 38860 692400 39120 692560
rect 39280 692400 39320 692560
rect 24580 692360 39320 692400
rect 24440 692340 39320 692360
rect 24440 692300 38700 692340
rect 24440 692180 24460 692300
rect 24580 692180 38700 692300
rect 38860 692180 39120 692340
rect 39280 692180 39320 692340
rect 24440 692140 39320 692180
rect 12890 691900 13110 691905
rect 12890 691700 12900 691900
rect 13100 691700 13110 691900
rect 12890 691695 13110 691700
rect 13190 691900 13410 691905
rect 13190 691700 13200 691900
rect 13400 691700 13410 691900
rect 13190 691695 13410 691700
rect 13490 691900 13710 691905
rect 13490 691700 13500 691900
rect 13700 691700 13710 691900
rect 13490 691695 13710 691700
rect 13790 691900 14010 691905
rect 13790 691700 13800 691900
rect 14000 691700 14010 691900
rect 13790 691695 14010 691700
rect 46320 691900 62200 692040
rect 46320 691700 58000 691900
rect 58200 691700 58400 691900
rect 58600 691700 58800 691900
rect 59000 691700 59200 691900
rect 59400 691700 59600 691900
rect 59800 691700 60000 691900
rect 60200 691700 60400 691900
rect 60600 691700 60800 691900
rect 61000 691700 61200 691900
rect 61400 691700 61600 691900
rect 61800 691700 62200 691900
rect 46320 691560 62200 691700
rect 465100 690500 470600 703700
rect 510400 701600 525470 704000
rect 510400 701400 515700 701600
rect 515900 701400 516100 701600
rect 516300 701400 516500 701600
rect 516700 701400 516900 701600
rect 517100 701400 517300 701600
rect 517500 701400 517700 701600
rect 517900 701400 518100 701600
rect 518300 701400 518500 701600
rect 518700 701400 518900 701600
rect 519100 701400 519300 701600
rect 519500 701400 519700 701600
rect 519900 701400 520100 701600
rect 520300 701400 520500 701600
rect 520700 701400 525470 701600
rect 510400 701200 525470 701400
rect 510400 701000 515700 701200
rect 515900 701000 516100 701200
rect 516300 701000 516500 701200
rect 516700 701000 516900 701200
rect 517100 701000 517300 701200
rect 517500 701000 517700 701200
rect 517900 701000 518100 701200
rect 518300 701000 518500 701200
rect 518700 701000 518900 701200
rect 519100 701000 519300 701200
rect 519500 701000 519700 701200
rect 519900 701000 520100 701200
rect 520300 701000 520500 701200
rect 520700 701000 525470 701200
rect 510400 700800 525470 701000
rect 510400 700600 515700 700800
rect 515900 700600 516100 700800
rect 516300 700600 516500 700800
rect 516700 700600 516900 700800
rect 517100 700600 517300 700800
rect 517500 700600 517700 700800
rect 517900 700600 518100 700800
rect 518300 700600 518500 700800
rect 518700 700600 518900 700800
rect 519100 700600 519300 700800
rect 519500 700600 519700 700800
rect 519900 700600 520100 700800
rect 520300 700600 520500 700800
rect 520700 700600 525470 700800
rect 510400 700400 525470 700600
rect 510400 700200 515700 700400
rect 515900 700200 516100 700400
rect 516300 700200 516500 700400
rect 516700 700200 516900 700400
rect 517100 700200 517300 700400
rect 517500 700200 517700 700400
rect 517900 700200 518100 700400
rect 518300 700200 518500 700400
rect 518700 700200 518900 700400
rect 519100 700200 519300 700400
rect 519500 700200 519700 700400
rect 519900 700200 520100 700400
rect 520300 700200 520500 700400
rect 520700 700200 525470 700400
rect 510400 700000 525470 700200
rect 510400 699800 515700 700000
rect 515900 699800 516100 700000
rect 516300 699800 516500 700000
rect 516700 699800 516900 700000
rect 517100 699800 517300 700000
rect 517500 699800 517700 700000
rect 517900 699800 518100 700000
rect 518300 699800 518500 700000
rect 518700 699800 518900 700000
rect 519100 699800 519300 700000
rect 519500 699800 519700 700000
rect 519900 699800 520100 700000
rect 520300 699800 520500 700000
rect 520700 699800 525470 700000
rect 510400 699600 525470 699800
rect 510400 699400 515700 699600
rect 515900 699400 516100 699600
rect 516300 699400 516500 699600
rect 516700 699400 516900 699600
rect 517100 699400 517300 699600
rect 517500 699400 517700 699600
rect 517900 699400 518100 699600
rect 518300 699400 518500 699600
rect 518700 699400 518900 699600
rect 519100 699400 519300 699600
rect 519500 699400 519700 699600
rect 519900 699400 520100 699600
rect 520300 699400 520500 699600
rect 520700 699400 525470 699600
rect 510400 699200 525470 699400
rect 510400 699000 515700 699200
rect 515900 699000 516100 699200
rect 516300 699000 516500 699200
rect 516700 699000 516900 699200
rect 517100 699000 517300 699200
rect 517500 699000 517700 699200
rect 517900 699000 518100 699200
rect 518300 699000 518500 699200
rect 518700 699000 518900 699200
rect 519100 699000 519300 699200
rect 519500 699000 519700 699200
rect 519900 699000 520100 699200
rect 520300 699000 520500 699200
rect 520700 699000 525470 699200
rect 510400 698600 525470 699000
rect 560300 702120 565120 702400
rect 560300 702020 563840 702120
rect 563940 702020 563980 702120
rect 564080 702020 564120 702120
rect 564220 702020 564260 702120
rect 564360 702020 564400 702120
rect 564500 702020 564540 702120
rect 564640 702020 564680 702120
rect 564780 702020 564820 702120
rect 564920 702020 564960 702120
rect 565060 702020 565120 702120
rect 560300 701980 565120 702020
rect 560300 701880 563840 701980
rect 563940 701880 563980 701980
rect 564080 701880 564120 701980
rect 564220 701880 564260 701980
rect 564360 701880 564400 701980
rect 564500 701880 564540 701980
rect 564640 701880 564680 701980
rect 564780 701880 564820 701980
rect 564920 701880 564960 701980
rect 565060 701880 565120 701980
rect 560300 701800 565120 701880
rect 566200 702280 572000 704000
rect 566200 702240 574140 702280
rect 566200 702140 573280 702240
rect 573380 702140 573420 702240
rect 573520 702140 573560 702240
rect 573660 702140 573700 702240
rect 573800 702140 573840 702240
rect 573940 702140 573980 702240
rect 574080 702140 574140 702240
rect 566200 701980 574140 702140
rect 566200 701880 573280 701980
rect 573380 701880 573420 701980
rect 573520 701880 573560 701980
rect 573660 701880 573700 701980
rect 573800 701880 573840 701980
rect 573940 701880 573980 701980
rect 574080 701880 574140 701980
rect 566200 701840 574140 701880
rect 560300 697600 561600 701800
rect 566200 698160 572000 701840
rect 515500 697400 561600 697600
rect 515500 697200 515700 697400
rect 515900 697200 516100 697400
rect 516300 697200 516500 697400
rect 516700 697200 516900 697400
rect 517100 697200 517300 697400
rect 517500 697200 517700 697400
rect 517900 697200 518100 697400
rect 518300 697200 518500 697400
rect 518700 697200 518900 697400
rect 519100 697200 519300 697400
rect 519500 697200 519700 697400
rect 519900 697200 520100 697400
rect 520300 697200 520500 697400
rect 520700 697200 561600 697400
rect 515500 697000 561600 697200
rect 515500 696800 515700 697000
rect 515900 696800 516100 697000
rect 516300 696800 516500 697000
rect 516700 696800 516900 697000
rect 517100 696800 517300 697000
rect 517500 696800 517700 697000
rect 517900 696800 518100 697000
rect 518300 696800 518500 697000
rect 518700 696800 518900 697000
rect 519100 696800 519300 697000
rect 519500 696800 519700 697000
rect 519900 696800 520100 697000
rect 520300 696800 520500 697000
rect 520700 696800 561600 697000
rect 515500 696600 561600 696800
rect 515500 696400 515700 696600
rect 515900 696400 516100 696600
rect 516300 696400 516500 696600
rect 516700 696400 516900 696600
rect 517100 696400 517300 696600
rect 517500 696400 517700 696600
rect 517900 696400 518100 696600
rect 518300 696400 518500 696600
rect 518700 696400 518900 696600
rect 519100 696400 519300 696600
rect 519500 696400 519700 696600
rect 519900 696400 520100 696600
rect 520300 696400 520500 696600
rect 520700 696400 561600 696600
rect 515500 696000 561600 696400
rect 563800 696220 572000 698160
rect 566200 691100 572000 696220
rect 573100 698000 574220 698180
rect 573100 697800 573300 698000
rect 573500 697800 573800 698000
rect 574000 697800 574220 698000
rect 573100 697600 574220 697800
rect 573100 697400 573300 697600
rect 573500 697400 573800 697600
rect 574000 697400 574220 697600
rect 573100 697200 574220 697400
rect 573100 697000 573300 697200
rect 573500 697000 573800 697200
rect 574000 697000 574220 697200
rect 573100 696800 574220 697000
rect 573100 696600 573300 696800
rect 573500 696600 573800 696800
rect 574000 696600 574220 696800
rect 573100 696400 574220 696600
rect 573100 696200 573300 696400
rect 573500 696200 573800 696400
rect 574000 696200 574220 696400
rect 573100 696100 574220 696200
rect 566200 690900 566300 691100
rect 566500 690900 566700 691100
rect 566900 690900 567100 691100
rect 567300 690900 567500 691100
rect 567700 690900 567900 691100
rect 568100 690900 568300 691100
rect 568500 690900 568700 691100
rect 568900 690900 569100 691100
rect 569300 690900 569500 691100
rect 569700 690900 569900 691100
rect 570100 690900 570300 691100
rect 570500 690900 570700 691100
rect 570900 690900 571100 691100
rect 571300 690900 571500 691100
rect 571700 690900 572000 691100
rect 566200 690700 572000 690900
rect 566200 690500 566300 690700
rect 566500 690500 566700 690700
rect 566900 690500 567100 690700
rect 567300 690500 567500 690700
rect 567700 690500 567900 690700
rect 568100 690500 568300 690700
rect 568500 690500 568700 690700
rect 568900 690500 569100 690700
rect 569300 690500 569500 690700
rect 569700 690500 569900 690700
rect 570100 690500 570300 690700
rect 570500 690500 570700 690700
rect 570900 690500 571100 690700
rect 571300 690500 571500 690700
rect 571700 690500 572000 690700
rect 465100 690400 534200 690500
rect 47100 690300 73200 690400
rect 47100 690200 47200 690300
rect 47300 690200 73200 690300
rect 47100 690000 68400 690200
rect 68600 690000 68800 690200
rect 69000 690000 69200 690200
rect 69400 690000 69600 690200
rect 69800 690000 70000 690200
rect 70200 690000 70400 690200
rect 70600 690000 70800 690200
rect 71000 690000 71200 690200
rect 71400 690000 71600 690200
rect 71800 690000 72000 690200
rect 72200 690000 72400 690200
rect 72600 690000 72800 690200
rect 73000 690000 73200 690200
rect 47100 689800 47200 690000
rect 47300 689800 73200 690000
rect 47100 689600 68400 689800
rect 68600 689600 68800 689800
rect 69000 689600 69200 689800
rect 69400 689600 69600 689800
rect 69800 689600 70000 689800
rect 70200 689600 70400 689800
rect 70600 689600 70800 689800
rect 71000 689600 71200 689800
rect 71400 689600 71600 689800
rect 71800 689600 72000 689800
rect 72200 689600 72400 689800
rect 72600 689600 72800 689800
rect 73000 689600 73200 689800
rect 47100 689500 47200 689600
rect 47300 689500 73200 689600
rect 47100 689400 73200 689500
rect 465100 690200 532300 690400
rect 532500 690200 532700 690400
rect 532900 690200 533100 690400
rect 533300 690200 533500 690400
rect 533700 690200 533900 690400
rect 534100 690200 534200 690400
rect 465100 690100 534200 690200
rect 465100 689900 532300 690100
rect 532500 689900 532700 690100
rect 532900 689900 533100 690100
rect 533300 689900 533500 690100
rect 533700 689900 533900 690100
rect 534100 689900 534200 690100
rect 465100 689700 534200 689900
rect 465100 689500 532300 689700
rect 532500 689500 532700 689700
rect 532900 689500 533100 689700
rect 533300 689500 533500 689700
rect 533700 689500 533900 689700
rect 534100 689500 534200 689700
rect 465100 689300 534200 689500
rect 465100 689100 532300 689300
rect 532500 689100 532700 689300
rect 532900 689100 533100 689300
rect 533300 689100 533500 689300
rect 533700 689100 533900 689300
rect 534100 689100 534200 689300
rect 566200 690300 572000 690500
rect 566200 690100 566300 690300
rect 566500 690100 566700 690300
rect 566900 690100 567100 690300
rect 567300 690100 567500 690300
rect 567700 690100 567900 690300
rect 568100 690100 568300 690300
rect 568500 690100 568700 690300
rect 568900 690100 569100 690300
rect 569300 690100 569500 690300
rect 569700 690100 569900 690300
rect 570100 690100 570300 690300
rect 570500 690100 570700 690300
rect 570900 690100 571100 690300
rect 571300 690100 571500 690300
rect 571700 690100 572000 690300
rect 566200 689900 572000 690100
rect 566200 689700 566300 689900
rect 566500 689700 566700 689900
rect 566900 689700 567100 689900
rect 567300 689700 567500 689900
rect 567700 689700 567900 689900
rect 568100 689700 568300 689900
rect 568500 689700 568700 689900
rect 568900 689700 569100 689900
rect 569300 689700 569500 689900
rect 569700 689700 569900 689900
rect 570100 689700 570300 689900
rect 570500 689700 570700 689900
rect 570900 689700 571100 689900
rect 571300 689700 571500 689900
rect 571700 689700 572000 689900
rect 566200 689500 572000 689700
rect 566200 689300 566300 689500
rect 566500 689300 566700 689500
rect 566900 689300 567100 689500
rect 567300 689300 567500 689500
rect 567700 689300 567900 689500
rect 568100 689300 568300 689500
rect 568500 689300 568700 689500
rect 568900 689300 569100 689500
rect 569300 689300 569500 689500
rect 569700 689300 569900 689500
rect 570100 689300 570300 689500
rect 570500 689300 570700 689500
rect 570900 689300 571100 689500
rect 571300 689300 571500 689500
rect 571700 689300 572000 689500
rect 566200 689200 572000 689300
rect 465100 688900 534200 689100
rect 16200 688700 42200 688800
rect 16200 688500 16400 688700
rect 16600 688500 16800 688700
rect 17000 688500 17200 688700
rect 17400 688500 17600 688700
rect 17800 688500 18000 688700
rect 18200 688500 18400 688700
rect 18600 688500 18800 688700
rect 19000 688500 19200 688700
rect 19400 688500 19600 688700
rect 19800 688500 20000 688700
rect 20200 688500 20400 688700
rect 20600 688500 20800 688700
rect 21000 688600 42000 688700
rect 42100 688600 42200 688700
rect 465100 688700 532300 688900
rect 532500 688700 532700 688900
rect 532900 688700 533100 688900
rect 533300 688700 533500 688900
rect 533700 688700 533900 688900
rect 534100 688700 534200 688900
rect 465100 688600 534200 688700
rect 21000 688500 42200 688600
rect 16200 688300 42000 688500
rect 42100 688300 42200 688500
rect 16200 688100 16400 688300
rect 16600 688100 16800 688300
rect 17000 688100 17200 688300
rect 17400 688100 17600 688300
rect 17800 688100 18000 688300
rect 18200 688100 18400 688300
rect 18600 688100 18800 688300
rect 19000 688100 19200 688300
rect 19400 688100 19600 688300
rect 19800 688100 20000 688300
rect 20200 688100 20400 688300
rect 20600 688100 20800 688300
rect 21000 688200 42200 688300
rect 21000 688100 42000 688200
rect 42100 688100 42200 688200
rect 16200 688000 42200 688100
rect 36600 687300 47800 687400
rect 36600 687100 36800 687300
rect 37000 687100 37200 687300
rect 37400 687100 37600 687300
rect 37800 687100 38000 687300
rect 38200 687100 47800 687300
rect 36600 687000 47800 687100
rect 549890 687000 549900 687200
rect 550100 687000 550110 687200
rect 550190 687000 550200 687200
rect 550400 687000 550410 687200
rect 550490 687000 550500 687200
rect 550700 687000 550710 687200
rect 550790 687000 550800 687200
rect 551000 687000 551010 687200
rect 551190 687100 551200 687300
rect 551400 687100 551410 687300
rect 551190 686800 551200 687000
rect 551400 686800 551410 687000
rect 551190 686500 551200 686700
rect 551400 686500 551410 686700
rect 551190 686200 551200 686400
rect 551400 686200 551410 686400
rect 549790 685900 549800 686100
rect 550000 685900 550010 686100
rect 550090 685900 550100 686100
rect 550300 685900 550310 686100
rect 550390 685900 550400 686100
rect 550600 685900 550610 686100
rect 550790 685900 550800 686100
rect 551000 685900 551010 686100
rect 0 685300 38400 685400
rect 0 685242 36800 685300
rect -800 685100 36800 685242
rect 37000 685100 37200 685300
rect 37400 685100 37600 685300
rect 37800 685100 38000 685300
rect 38200 685100 38400 685300
rect -800 684900 38400 685100
rect -800 684700 36800 684900
rect 37000 684700 37200 684900
rect 37400 684700 37600 684900
rect 37800 684700 38000 684900
rect 38200 684700 38400 684900
rect -800 684500 38400 684700
rect -800 684300 36800 684500
rect 37000 684300 37200 684500
rect 37400 684300 37600 684500
rect 37800 684300 38000 684500
rect 38200 684300 38400 684500
rect -800 684100 38400 684300
rect -800 683900 36800 684100
rect 37000 683900 37200 684100
rect 37400 683900 37600 684100
rect 37800 683900 38000 684100
rect 38200 683900 38400 684100
rect -800 683700 38400 683900
rect -800 683500 36800 683700
rect 37000 683500 37200 683700
rect 37400 683500 37600 683700
rect 37800 683500 38000 683700
rect 38200 683500 38400 683700
rect -800 683300 38400 683500
rect -800 683100 36800 683300
rect 37000 683100 37200 683300
rect 37400 683100 37600 683300
rect 37800 683100 38000 683300
rect 38200 683100 38400 683300
rect 515500 684800 540560 684940
rect 515500 684600 515700 684800
rect 515900 684600 516100 684800
rect 516300 684600 516500 684800
rect 516700 684600 516900 684800
rect 517100 684600 517300 684800
rect 517500 684600 517700 684800
rect 517900 684600 518100 684800
rect 518300 684600 518500 684800
rect 518700 684600 518900 684800
rect 519100 684600 519300 684800
rect 519500 684600 519700 684800
rect 519900 684600 520100 684800
rect 520300 684600 520500 684800
rect 520700 684600 540560 684800
rect 515500 684400 540560 684600
rect 515500 684200 515700 684400
rect 515900 684200 516100 684400
rect 516300 684200 516500 684400
rect 516700 684200 516900 684400
rect 517100 684200 517300 684400
rect 517500 684200 517700 684400
rect 517900 684200 518100 684400
rect 518300 684200 518500 684400
rect 518700 684200 518900 684400
rect 519100 684200 519300 684400
rect 519500 684200 519700 684400
rect 519900 684200 520100 684400
rect 520300 684200 520500 684400
rect 520700 684200 540560 684400
rect 515500 684000 540560 684200
rect 515500 683800 515700 684000
rect 515900 683800 516100 684000
rect 516300 683800 516500 684000
rect 516700 683800 516900 684000
rect 517100 683800 517300 684000
rect 517500 683800 517700 684000
rect 517900 683800 518100 684000
rect 518300 683800 518500 684000
rect 518700 683800 518900 684000
rect 519100 683800 519300 684000
rect 519500 683800 519700 684000
rect 519900 683800 520100 684000
rect 520300 683800 520500 684000
rect 520700 683800 540560 684000
rect 515500 683600 540560 683800
rect 576600 684700 578700 684900
rect 576600 684400 576800 684700
rect 577100 684400 577300 684700
rect 577600 684400 577800 684700
rect 578100 684400 578300 684700
rect 578600 684400 578700 684700
rect 576600 684200 578700 684400
rect 576600 683900 576800 684200
rect 577100 683900 577300 684200
rect 577600 683900 577800 684200
rect 578100 683900 578300 684200
rect 578600 683900 578700 684200
rect 576600 683600 578700 683900
rect 582320 684600 582660 684660
rect 582320 684520 582360 684600
rect 582440 684520 582540 684600
rect 582620 684520 582660 684600
rect 582320 684440 582660 684520
rect 582320 684360 582360 684440
rect 582440 684360 582540 684440
rect 582620 684360 582660 684440
rect 582320 684280 582660 684360
rect 582320 684200 582360 684280
rect 582440 684200 582540 684280
rect 582620 684200 582660 684280
rect 582320 684100 582660 684200
rect 582320 684020 582360 684100
rect 582440 684020 582540 684100
rect 582620 684020 582660 684100
rect 582320 683940 582660 684020
rect 582320 683860 582360 683940
rect 582440 683860 582540 683940
rect 582620 683860 582660 683940
rect 515500 683400 515700 683600
rect 515900 683400 516100 683600
rect 516300 683400 516500 683600
rect 516700 683400 516900 683600
rect 517100 683400 517300 683600
rect 517500 683400 517700 683600
rect 517900 683400 518100 683600
rect 518300 683400 518500 683600
rect 518700 683400 518900 683600
rect 519100 683400 519300 683600
rect 519500 683400 519700 683600
rect 519900 683400 520100 683600
rect 520300 683400 520500 683600
rect 520700 683400 540560 683600
rect 515500 683200 540560 683400
rect 582320 683200 582660 683860
rect -800 682900 38400 683100
rect 42240 683120 43910 683140
rect 42240 683040 42260 683120
rect 42340 683040 42400 683120
rect 42480 683040 42540 683120
rect 42620 683040 43910 683120
rect 42240 683020 43910 683040
rect 45360 683120 47040 683140
rect 45360 683040 46660 683120
rect 46740 683040 46800 683120
rect 46880 683040 46940 683120
rect 47020 683040 47040 683120
rect 45360 683020 47040 683040
rect -800 682700 36800 682900
rect 37000 682700 37200 682900
rect 37400 682700 37600 682900
rect 37800 682700 38000 682900
rect 38200 682700 38400 682900
rect -800 682500 38400 682700
rect -800 682300 36800 682500
rect 37000 682300 37200 682500
rect 37400 682300 37600 682500
rect 37800 682300 38000 682500
rect 38200 682300 38400 682500
rect 515500 683000 515700 683200
rect 515900 683000 516100 683200
rect 516300 683000 516500 683200
rect 516700 683000 516900 683200
rect 517100 683000 517300 683200
rect 517500 683000 517700 683200
rect 517900 683000 518100 683200
rect 518300 683000 518500 683200
rect 518700 683000 518900 683200
rect 519100 683000 519300 683200
rect 519500 683000 519700 683200
rect 519900 683000 520100 683200
rect 520300 683000 520500 683200
rect 520700 683000 540560 683200
rect 515500 682800 540560 683000
rect 515500 682600 515700 682800
rect 515900 682600 516100 682800
rect 516300 682600 516500 682800
rect 516700 682600 516900 682800
rect 517100 682600 517300 682800
rect 517500 682600 517700 682800
rect 517900 682600 518100 682800
rect 518300 682600 518500 682800
rect 518700 682600 518900 682800
rect 519100 682600 519300 682800
rect 519500 682600 519700 682800
rect 519900 682600 520100 682800
rect 520300 682600 520500 682800
rect 520700 682600 540560 682800
rect 515500 682460 540560 682600
rect 561600 682984 584000 683200
rect 515500 682400 515600 682460
rect -800 682100 38400 682300
rect -800 681900 36800 682100
rect 37000 681900 37200 682100
rect 37400 681900 37600 682100
rect 37800 681900 38000 682100
rect 38200 681900 38400 682100
rect -800 681700 38400 681900
rect 45440 682200 62200 682320
rect 45440 682000 58000 682200
rect 58200 682000 58400 682200
rect 58600 682000 58800 682200
rect 59000 682000 59200 682200
rect 59400 682000 59600 682200
rect 59800 682000 60000 682200
rect 60200 682000 60400 682200
rect 60600 682000 60800 682200
rect 61000 682000 61200 682200
rect 61400 682000 61600 682200
rect 61800 682000 62200 682200
rect 45440 681860 62200 682000
rect 561600 682200 584800 682984
rect 561600 682000 561700 682200
rect 561900 682000 562100 682200
rect 562300 682000 562500 682200
rect 562700 682000 562900 682200
rect 563100 682000 563300 682200
rect 563500 682000 584800 682200
rect -800 681500 36800 681700
rect 37000 681500 37200 681700
rect 37400 681500 37600 681700
rect 37800 681500 38000 681700
rect 38200 681500 38400 681700
rect 561600 681800 584800 682000
rect 561600 681600 561700 681800
rect 561900 681600 562100 681800
rect 562300 681600 562500 681800
rect 562700 681600 562900 681800
rect 563100 681600 563300 681800
rect 563500 681600 584800 681800
rect -800 681300 38400 681500
rect -800 681100 36800 681300
rect 37000 681100 37200 681300
rect 37400 681100 37600 681300
rect 37800 681100 38000 681300
rect 38200 681100 38400 681300
rect -800 680900 38400 681100
rect -800 680700 36800 680900
rect 37000 680700 37200 680900
rect 37400 680700 37600 680900
rect 37800 680700 38000 680900
rect 38200 680700 38400 680900
rect 547600 681400 553100 681500
rect 547600 681200 549800 681400
rect 550000 681200 550200 681400
rect 550400 681200 550600 681400
rect 550800 681200 551000 681400
rect 551200 681200 551400 681400
rect 551600 681200 551800 681400
rect 552000 681200 552200 681400
rect 552400 681200 552600 681400
rect 552800 681200 553100 681400
rect 547600 681000 553100 681200
rect 547600 680800 549800 681000
rect 550000 680800 550200 681000
rect 550400 680800 550600 681000
rect 550800 680800 551000 681000
rect 551200 680800 551400 681000
rect 551600 680800 551800 681000
rect 552000 680800 552200 681000
rect 552400 680800 552600 681000
rect 552800 680800 553100 681000
rect 547600 680700 553100 680800
rect 561600 681400 584800 681600
rect 561600 681200 561700 681400
rect 561900 681200 562100 681400
rect 562300 681200 562500 681400
rect 562700 681200 562900 681400
rect 563100 681200 563300 681400
rect 563500 681200 584800 681400
rect 561600 681000 584800 681200
rect 561600 680800 561700 681000
rect 561900 680800 562100 681000
rect 562300 680800 562500 681000
rect 562700 680800 562900 681000
rect 563100 680800 563300 681000
rect 563500 680800 584800 681000
rect -800 680500 38400 680700
rect -800 680300 36800 680500
rect 37000 680300 37200 680500
rect 37400 680300 37600 680500
rect 37800 680300 38000 680500
rect 38200 680300 38400 680500
rect -800 680242 38400 680300
rect 0 680200 38400 680242
rect 561600 680600 584800 680800
rect 561600 680400 561700 680600
rect 561900 680400 562100 680600
rect 562300 680400 562500 680600
rect 562700 680400 562900 680600
rect 563100 680400 563300 680600
rect 563500 680400 584800 680600
rect 561600 680200 584800 680400
rect 561600 680000 561700 680200
rect 561900 680000 562100 680200
rect 562300 680000 562500 680200
rect 562700 680000 562900 680200
rect 563100 680000 563300 680200
rect 563500 680000 584800 680200
rect 561600 679800 584800 680000
rect 561600 679600 561700 679800
rect 561900 679600 562100 679800
rect 562300 679600 562500 679800
rect 562700 679600 562900 679800
rect 563100 679600 563300 679800
rect 563500 679600 584800 679800
rect 515500 679200 541760 679560
rect 515500 679000 515900 679200
rect 516100 679000 516300 679200
rect 516500 679000 516700 679200
rect 516900 679000 517100 679200
rect 517300 679000 517500 679200
rect 517700 679000 517900 679200
rect 518100 679000 518300 679200
rect 518500 679000 518700 679200
rect 518900 679000 519100 679200
rect 519300 679000 519500 679200
rect 519700 679000 519900 679200
rect 520100 679000 520300 679200
rect 520500 679000 520700 679200
rect 520900 679000 541760 679200
rect 515500 678800 541760 679000
rect 515500 678600 515900 678800
rect 516100 678600 516300 678800
rect 516500 678600 516700 678800
rect 516900 678600 517100 678800
rect 517300 678600 517500 678800
rect 517700 678600 517900 678800
rect 518100 678600 518300 678800
rect 518500 678600 518700 678800
rect 518900 678600 519100 678800
rect 519300 678600 519500 678800
rect 519700 678600 519900 678800
rect 520100 678600 520300 678800
rect 520500 678600 520700 678800
rect 520900 678600 541760 678800
rect 515500 678400 541760 678600
rect 515500 678200 515900 678400
rect 516100 678200 516300 678400
rect 516500 678200 516700 678400
rect 516900 678200 517100 678400
rect 517300 678200 517500 678400
rect 517700 678200 517900 678400
rect 518100 678200 518300 678400
rect 518500 678200 518700 678400
rect 518900 678200 519100 678400
rect 519300 678200 519500 678400
rect 519700 678200 519900 678400
rect 520100 678200 520300 678400
rect 520500 678200 520700 678400
rect 520900 678200 541760 678400
rect 515500 678000 541760 678200
rect 515500 677800 515900 678000
rect 516100 677800 516300 678000
rect 516500 677800 516700 678000
rect 516900 677800 517100 678000
rect 517300 677800 517500 678000
rect 517700 677800 517900 678000
rect 518100 677800 518300 678000
rect 518500 677800 518700 678000
rect 518900 677800 519100 678000
rect 519300 677800 519500 678000
rect 519700 677800 519900 678000
rect 520100 677800 520300 678000
rect 520500 677800 520700 678000
rect 520900 677800 541760 678000
rect 561600 679400 584800 679600
rect 561600 679200 561700 679400
rect 561900 679200 562100 679400
rect 562300 679200 562500 679400
rect 562700 679200 562900 679400
rect 563100 679200 563300 679400
rect 563500 679200 584800 679400
rect 561600 679000 584800 679200
rect 561600 678800 561700 679000
rect 561900 678800 562100 679000
rect 562300 678800 562500 679000
rect 562700 678800 562900 679000
rect 563100 678800 563300 679000
rect 563500 678800 584800 679000
rect 561600 678600 584800 678800
rect 561600 678400 561700 678600
rect 561900 678400 562100 678600
rect 562300 678400 562500 678600
rect 562700 678400 562900 678600
rect 563100 678400 563300 678600
rect 563500 678400 584800 678600
rect 561600 677984 584800 678400
rect 561600 677800 584000 677984
rect 515500 677600 541760 677800
rect 515500 677400 515900 677600
rect 516100 677400 516300 677600
rect 516500 677400 516700 677600
rect 516900 677400 517100 677600
rect 517300 677400 517500 677600
rect 517700 677400 517900 677600
rect 518100 677400 518300 677600
rect 518500 677400 518700 677600
rect 518900 677400 519100 677600
rect 519300 677400 519500 677600
rect 519700 677400 519900 677600
rect 520100 677400 520300 677600
rect 520500 677400 520700 677600
rect 520900 677400 541760 677600
rect 515500 677200 541760 677400
rect 515500 677000 515900 677200
rect 516100 677000 516300 677200
rect 516500 677000 516700 677200
rect 516900 677000 517100 677200
rect 517300 677000 517500 677200
rect 517700 677000 517900 677200
rect 518100 677000 518300 677200
rect 518500 677000 518700 677200
rect 518900 677000 519100 677200
rect 519300 677000 519500 677200
rect 519700 677000 519900 677200
rect 520100 677000 520300 677200
rect 520500 677000 520700 677200
rect 520900 677000 541760 677200
rect 515500 676800 541760 677000
rect 515500 676600 515900 676800
rect 516100 676600 516300 676800
rect 516500 676600 516700 676800
rect 516900 676600 517100 676800
rect 517300 676600 517500 676800
rect 517700 676600 517900 676800
rect 518100 676600 518300 676800
rect 518500 676600 518700 676800
rect 518900 676600 519100 676800
rect 519300 676600 519500 676800
rect 519700 676600 519900 676800
rect 520100 676600 520300 676800
rect 520500 676600 520700 676800
rect 520900 676600 541760 676800
rect 515500 676460 541760 676600
rect 547600 677300 572280 677400
rect 547600 677100 571900 677300
rect 572100 677100 572280 677300
rect 547600 677000 572280 677100
rect 547600 676800 571900 677000
rect 572100 676800 572280 677000
rect 547600 676700 572280 676800
rect 547600 676500 571900 676700
rect 572100 676500 572280 676700
rect 547600 676400 572280 676500
rect 547600 676200 571900 676400
rect 572100 676200 572280 676400
rect 547600 676100 572280 676200
rect 576700 676100 578700 677800
rect 32790 663300 33110 663305
rect 32790 663000 32800 663300
rect 33100 663000 33110 663300
rect 32790 662995 33110 663000
rect 33290 663300 33610 663305
rect 33290 663000 33300 663300
rect 33600 663000 33610 663300
rect 33290 662995 33610 663000
rect 33790 663300 34110 663305
rect 33790 663000 33800 663300
rect 34100 663000 34110 663300
rect 33790 662995 34110 663000
rect 34290 663300 34610 663305
rect 34290 663000 34300 663300
rect 34600 663000 34610 663300
rect 34290 662995 34610 663000
rect 34790 663300 35110 663305
rect 34790 663000 34800 663300
rect 35100 663000 35110 663300
rect 34790 662995 35110 663000
rect 35290 663300 35610 663305
rect 35290 663000 35300 663300
rect 35600 663000 35610 663300
rect 35290 662995 35610 663000
rect 35790 663300 36110 663305
rect 35790 663000 35800 663300
rect 36100 663000 36110 663300
rect 35790 662995 36110 663000
rect 36290 663300 36610 663305
rect 36290 663000 36300 663300
rect 36600 663000 36610 663300
rect 36290 662995 36610 663000
rect 36790 663300 37110 663305
rect 36790 663000 36800 663300
rect 37100 663000 37110 663300
rect 36790 662995 37110 663000
rect 37290 663300 37610 663305
rect 37290 663000 37300 663300
rect 37600 663000 37610 663300
rect 37290 662995 37610 663000
rect 37790 663300 38110 663305
rect 37790 663000 37800 663300
rect 38100 663000 38110 663300
rect 37790 662995 38110 663000
rect 38290 663300 38610 663305
rect 38290 663000 38300 663300
rect 38600 663000 38610 663300
rect 38290 662995 38610 663000
rect 38790 663300 39110 663305
rect 38790 663000 38800 663300
rect 39100 663000 39110 663300
rect 38790 662995 39110 663000
rect 39290 663300 39610 663305
rect 39290 663000 39300 663300
rect 39600 663000 39610 663300
rect 39290 662995 39610 663000
rect 39790 663300 40110 663305
rect 39790 663000 39800 663300
rect 40100 663000 40110 663300
rect 39790 662995 40110 663000
rect 40290 663300 40610 663305
rect 40290 663000 40300 663300
rect 40600 663000 40610 663300
rect 40290 662995 40610 663000
rect 0 648642 4000 648800
rect -800 648600 4000 648642
rect -800 648300 2500 648600
rect 2800 648300 3000 648600
rect 3300 648300 3500 648600
rect 3800 648300 4000 648600
rect -800 648100 4000 648300
rect -800 647800 2500 648100
rect 2800 647800 3000 648100
rect 3300 647800 3500 648100
rect 3800 647800 4000 648100
rect -800 647600 4000 647800
rect -800 647300 2500 647600
rect 2800 647300 3000 647600
rect 3300 647300 3500 647600
rect 3800 647300 4000 647600
rect -800 647100 4000 647300
rect -800 646800 2500 647100
rect 2800 646800 3000 647100
rect 3300 646800 3500 647100
rect 3800 646800 4000 647100
rect -800 646600 4000 646800
rect -800 646300 2500 646600
rect 2800 646300 3000 646600
rect 3300 646300 3500 646600
rect 3800 646300 4000 646600
rect -800 646100 4000 646300
rect -800 645800 2500 646100
rect 2800 645800 3000 646100
rect 3300 645800 3500 646100
rect 3800 645800 4000 646100
rect -800 645600 4000 645800
rect -800 645300 2500 645600
rect 2800 645300 3000 645600
rect 3300 645300 3500 645600
rect 3800 645300 4000 645600
rect -800 645100 4000 645300
rect -800 644800 2500 645100
rect 2800 644800 3000 645100
rect 3300 644800 3500 645100
rect 3800 644800 4000 645100
rect -800 644600 4000 644800
rect -800 644300 2500 644600
rect 2800 644300 3000 644600
rect 3300 644300 3500 644600
rect 3800 644300 4000 644600
rect -800 644100 4000 644300
rect -800 643842 2500 644100
rect 0 643800 2500 643842
rect 2800 643800 3000 644100
rect 3300 643800 3500 644100
rect 3800 643800 4000 644100
rect 0 643600 4000 643800
rect 0 643300 2500 643600
rect 2800 643300 3000 643600
rect 3300 643300 3500 643600
rect 3800 643300 4000 643600
rect 0 643100 4000 643300
rect 0 642800 2500 643100
rect 2800 642800 3000 643100
rect 3300 642800 3500 643100
rect 3800 642800 4000 643100
rect 0 642600 4000 642800
rect 0 642300 2500 642600
rect 2800 642300 3000 642600
rect 3300 642300 3500 642600
rect 3800 642300 4000 642600
rect 0 642100 4000 642300
rect 0 641800 2500 642100
rect 2800 641800 3000 642100
rect 3300 641800 3500 642100
rect 3800 641800 4000 642100
rect 0 641600 4000 641800
rect 0 641300 2500 641600
rect 2800 641300 3000 641600
rect 3300 641300 3500 641600
rect 3800 641300 4000 641600
rect 0 641100 4000 641300
rect 0 640800 2500 641100
rect 2800 640800 3000 641100
rect 3300 640800 3500 641100
rect 3800 640800 4000 641100
rect 0 640600 4000 640800
rect 0 640300 2500 640600
rect 2800 640300 3000 640600
rect 3300 640300 3500 640600
rect 3800 640300 4000 640600
rect 0 640100 4000 640300
rect 0 639800 2500 640100
rect 2800 639800 3000 640100
rect 3300 639800 3500 640100
rect 3800 639800 4000 640100
rect 0 639600 4000 639800
rect 0 639300 2500 639600
rect 2800 639300 3000 639600
rect 3300 639300 3500 639600
rect 3800 639300 4000 639600
rect 0 639100 4000 639300
rect 0 638800 2500 639100
rect 2800 638800 3000 639100
rect 3300 638800 3500 639100
rect 3800 638800 4000 639100
rect 0 638642 4000 638800
rect -800 638600 4000 638642
rect -800 638300 2500 638600
rect 2800 638300 3000 638600
rect 3300 638300 3500 638600
rect 3800 638300 4000 638600
rect -800 638100 4000 638300
rect -800 637800 2500 638100
rect 2800 637800 3000 638100
rect 3300 637800 3500 638100
rect 3800 637800 4000 638100
rect -800 637600 4000 637800
rect -800 637300 2500 637600
rect 2800 637300 3000 637600
rect 3300 637300 3500 637600
rect 3800 637300 4000 637600
rect -800 637100 4000 637300
rect -800 636800 2500 637100
rect 2800 636800 3000 637100
rect 3300 636800 3500 637100
rect 3800 636800 4000 637100
rect -800 636600 4000 636800
rect -800 636300 2500 636600
rect 2800 636300 3000 636600
rect 3300 636300 3500 636600
rect 3800 636300 4000 636600
rect -800 636100 4000 636300
rect -800 635800 2500 636100
rect 2800 635800 3000 636100
rect 3300 635800 3500 636100
rect 3800 635800 4000 636100
rect -800 635600 4000 635800
rect -800 635300 2500 635600
rect 2800 635300 3000 635600
rect 3300 635300 3500 635600
rect 3800 635300 4000 635600
rect -800 635100 4000 635300
rect -800 634800 2500 635100
rect 2800 634800 3000 635100
rect 3300 634800 3500 635100
rect 3800 634800 4000 635100
rect -800 634600 4000 634800
rect -800 634300 2500 634600
rect 2800 634300 3000 634600
rect 3300 634300 3500 634600
rect 3800 634300 4000 634600
rect -800 633842 4000 634300
rect 0 633800 4000 633842
rect 549600 644600 584000 644800
rect 549600 644400 550000 644600
rect 550200 644400 550400 644600
rect 550600 644400 550800 644600
rect 551000 644400 551200 644600
rect 551400 644400 551600 644600
rect 551800 644400 552000 644600
rect 552200 644400 552400 644600
rect 552600 644400 552800 644600
rect 553000 644584 584000 644600
rect 553000 644400 584800 644584
rect 549600 644200 584800 644400
rect 549600 644000 550000 644200
rect 550200 644000 550400 644200
rect 550600 644000 550800 644200
rect 551000 644000 551200 644200
rect 551400 644000 551600 644200
rect 551800 644000 552000 644200
rect 552200 644000 552400 644200
rect 552600 644000 552800 644200
rect 553000 644000 584800 644200
rect 549600 643800 584800 644000
rect 549600 643600 550000 643800
rect 550200 643600 550400 643800
rect 550600 643600 550800 643800
rect 551000 643600 551200 643800
rect 551400 643600 551600 643800
rect 551800 643600 552000 643800
rect 552200 643600 552400 643800
rect 552600 643600 552800 643800
rect 553000 643600 584800 643800
rect 549600 643400 584800 643600
rect 549600 643200 550000 643400
rect 550200 643200 550400 643400
rect 550600 643200 550800 643400
rect 551000 643200 551200 643400
rect 551400 643200 551600 643400
rect 551800 643200 552000 643400
rect 552200 643200 552400 643400
rect 552600 643200 552800 643400
rect 553000 643200 584800 643400
rect 549600 643000 584800 643200
rect 549600 642800 550000 643000
rect 550200 642800 550400 643000
rect 550600 642800 550800 643000
rect 551000 642800 551200 643000
rect 551400 642800 551600 643000
rect 551800 642800 552000 643000
rect 552200 642800 552400 643000
rect 552600 642800 552800 643000
rect 553000 642800 584800 643000
rect 549600 642600 584800 642800
rect 549600 642400 550000 642600
rect 550200 642400 550400 642600
rect 550600 642400 550800 642600
rect 551000 642400 551200 642600
rect 551400 642400 551600 642600
rect 551800 642400 552000 642600
rect 552200 642400 552400 642600
rect 552600 642400 552800 642600
rect 553000 642400 584800 642600
rect 549600 642200 584800 642400
rect 549600 642000 550000 642200
rect 550200 642000 550400 642200
rect 550600 642000 550800 642200
rect 551000 642000 551200 642200
rect 551400 642000 551600 642200
rect 551800 642000 552000 642200
rect 552200 642000 552400 642200
rect 552600 642000 552800 642200
rect 553000 642000 584800 642200
rect 549600 641800 584800 642000
rect 549600 641600 550000 641800
rect 550200 641600 550400 641800
rect 550600 641600 550800 641800
rect 551000 641600 551200 641800
rect 551400 641600 551600 641800
rect 551800 641600 552000 641800
rect 552200 641600 552400 641800
rect 552600 641600 552800 641800
rect 553000 641600 584800 641800
rect 549600 641400 584800 641600
rect 549600 641200 550000 641400
rect 550200 641200 550400 641400
rect 550600 641200 550800 641400
rect 551000 641200 551200 641400
rect 551400 641200 551600 641400
rect 551800 641200 552000 641400
rect 552200 641200 552400 641400
rect 552600 641200 552800 641400
rect 553000 641200 584800 641400
rect 549600 641000 584800 641200
rect 549600 640800 550000 641000
rect 550200 640800 550400 641000
rect 550600 640800 550800 641000
rect 551000 640800 551200 641000
rect 551400 640800 551600 641000
rect 551800 640800 552000 641000
rect 552200 640800 552400 641000
rect 552600 640800 552800 641000
rect 553000 640800 584800 641000
rect 549600 640600 584800 640800
rect 549600 640400 550000 640600
rect 550200 640400 550400 640600
rect 550600 640400 550800 640600
rect 551000 640400 551200 640600
rect 551400 640400 551600 640600
rect 551800 640400 552000 640600
rect 552200 640400 552400 640600
rect 552600 640400 552800 640600
rect 553000 640400 584800 640600
rect 549600 640200 584800 640400
rect 549600 640000 550000 640200
rect 550200 640000 550400 640200
rect 550600 640000 550800 640200
rect 551000 640000 551200 640200
rect 551400 640000 551600 640200
rect 551800 640000 552000 640200
rect 552200 640000 552400 640200
rect 552600 640000 552800 640200
rect 553000 640000 584800 640200
rect 549600 639800 584800 640000
rect 549600 639600 550000 639800
rect 550200 639600 550400 639800
rect 550600 639600 550800 639800
rect 551000 639600 551200 639800
rect 551400 639600 551600 639800
rect 551800 639600 552000 639800
rect 552200 639600 552400 639800
rect 552600 639600 552800 639800
rect 553000 639784 584800 639800
rect 553000 639600 584000 639784
rect 549600 639400 584000 639600
rect 549600 639200 550000 639400
rect 550200 639200 550400 639400
rect 550600 639200 550800 639400
rect 551000 639200 551200 639400
rect 551400 639200 551600 639400
rect 551800 639200 552000 639400
rect 552200 639200 552400 639400
rect 552600 639200 552800 639400
rect 553000 639200 584000 639400
rect 549600 639000 584000 639200
rect 549600 638800 550000 639000
rect 550200 638800 550400 639000
rect 550600 638800 550800 639000
rect 551000 638800 551200 639000
rect 551400 638800 551600 639000
rect 551800 638800 552000 639000
rect 552200 638800 552400 639000
rect 552600 638800 552800 639000
rect 553000 638800 584000 639000
rect 549600 638600 584000 638800
rect 549600 638400 550000 638600
rect 550200 638400 550400 638600
rect 550600 638400 550800 638600
rect 551000 638400 551200 638600
rect 551400 638400 551600 638600
rect 551800 638400 552000 638600
rect 552200 638400 552400 638600
rect 552600 638400 552800 638600
rect 553000 638400 584000 638600
rect 549600 638200 584000 638400
rect 549600 638000 550000 638200
rect 550200 638000 550400 638200
rect 550600 638000 550800 638200
rect 551000 638000 551200 638200
rect 551400 638000 551600 638200
rect 551800 638000 552000 638200
rect 552200 638000 552400 638200
rect 552600 638000 552800 638200
rect 553000 638000 584000 638200
rect 549600 637800 584000 638000
rect 549600 637600 550000 637800
rect 550200 637600 550400 637800
rect 550600 637600 550800 637800
rect 551000 637600 551200 637800
rect 551400 637600 551600 637800
rect 551800 637600 552000 637800
rect 552200 637600 552400 637800
rect 552600 637600 552800 637800
rect 553000 637600 584000 637800
rect 549600 637400 584000 637600
rect 549600 637200 550000 637400
rect 550200 637200 550400 637400
rect 550600 637200 550800 637400
rect 551000 637200 551200 637400
rect 551400 637200 551600 637400
rect 551800 637200 552000 637400
rect 552200 637200 552400 637400
rect 552600 637200 552800 637400
rect 553000 637200 584000 637400
rect 549600 637000 584000 637200
rect 549600 636800 550000 637000
rect 550200 636800 550400 637000
rect 550600 636800 550800 637000
rect 551000 636800 551200 637000
rect 551400 636800 551600 637000
rect 551800 636800 552000 637000
rect 552200 636800 552400 637000
rect 552600 636800 552800 637000
rect 553000 636800 584000 637000
rect 549600 636600 584000 636800
rect 549600 636400 550000 636600
rect 550200 636400 550400 636600
rect 550600 636400 550800 636600
rect 551000 636400 551200 636600
rect 551400 636400 551600 636600
rect 551800 636400 552000 636600
rect 552200 636400 552400 636600
rect 552600 636400 552800 636600
rect 553000 636400 584000 636600
rect 549600 636200 584000 636400
rect 549600 636000 550000 636200
rect 550200 636000 550400 636200
rect 550600 636000 550800 636200
rect 551000 636000 551200 636200
rect 551400 636000 551600 636200
rect 551800 636000 552000 636200
rect 552200 636000 552400 636200
rect 552600 636000 552800 636200
rect 553000 636000 584000 636200
rect 549600 635800 584000 636000
rect 549600 635600 550000 635800
rect 550200 635600 550400 635800
rect 550600 635600 550800 635800
rect 551000 635600 551200 635800
rect 551400 635600 551600 635800
rect 551800 635600 552000 635800
rect 552200 635600 552400 635800
rect 552600 635600 552800 635800
rect 553000 635600 584000 635800
rect 549600 635400 584000 635600
rect 549600 635200 550000 635400
rect 550200 635200 550400 635400
rect 550600 635200 550800 635400
rect 551000 635200 551200 635400
rect 551400 635200 551600 635400
rect 551800 635200 552000 635400
rect 552200 635200 552400 635400
rect 552600 635200 552800 635400
rect 553000 635200 584000 635400
rect 549600 635000 584000 635200
rect 549600 634800 550000 635000
rect 550200 634800 550400 635000
rect 550600 634800 550800 635000
rect 551000 634800 551200 635000
rect 551400 634800 551600 635000
rect 551800 634800 552000 635000
rect 552200 634800 552400 635000
rect 552600 634800 552800 635000
rect 553000 634800 584000 635000
rect 549600 634600 584000 634800
rect 549600 634400 550000 634600
rect 550200 634400 550400 634600
rect 550600 634400 550800 634600
rect 551000 634400 551200 634600
rect 551400 634400 551600 634600
rect 551800 634400 552000 634600
rect 552200 634400 552400 634600
rect 552600 634400 552800 634600
rect 553000 634584 584000 634600
rect 553000 634400 584800 634584
rect 549600 634200 584800 634400
rect 549600 634000 550000 634200
rect 550200 634000 550400 634200
rect 550600 634000 550800 634200
rect 551000 634000 551200 634200
rect 551400 634000 551600 634200
rect 551800 634000 552000 634200
rect 552200 634000 552400 634200
rect 552600 634000 552800 634200
rect 553000 634000 584800 634200
rect 549600 633800 584800 634000
rect 549600 633600 550000 633800
rect 550200 633600 550400 633800
rect 550600 633600 550800 633800
rect 551000 633600 551200 633800
rect 551400 633600 551600 633800
rect 551800 633600 552000 633800
rect 552200 633600 552400 633800
rect 552600 633600 552800 633800
rect 553000 633600 584800 633800
rect 549600 633400 584800 633600
rect 549600 633200 550000 633400
rect 550200 633200 550400 633400
rect 550600 633200 550800 633400
rect 551000 633200 551200 633400
rect 551400 633200 551600 633400
rect 551800 633200 552000 633400
rect 552200 633200 552400 633400
rect 552600 633200 552800 633400
rect 553000 633200 584800 633400
rect 549600 633000 584800 633200
rect 549600 632800 550000 633000
rect 550200 632800 550400 633000
rect 550600 632800 550800 633000
rect 551000 632800 551200 633000
rect 551400 632800 551600 633000
rect 551800 632800 552000 633000
rect 552200 632800 552400 633000
rect 552600 632800 552800 633000
rect 553000 632800 584800 633000
rect 549600 632600 584800 632800
rect 549600 632400 550000 632600
rect 550200 632400 550400 632600
rect 550600 632400 550800 632600
rect 551000 632400 551200 632600
rect 551400 632400 551600 632600
rect 551800 632400 552000 632600
rect 552200 632400 552400 632600
rect 552600 632400 552800 632600
rect 553000 632400 584800 632600
rect 549600 632200 584800 632400
rect 549600 632000 550000 632200
rect 550200 632000 550400 632200
rect 550600 632000 550800 632200
rect 551000 632000 551200 632200
rect 551400 632000 551600 632200
rect 551800 632000 552000 632200
rect 552200 632000 552400 632200
rect 552600 632000 552800 632200
rect 553000 632000 584800 632200
rect 549600 631800 584800 632000
rect 549600 631600 550000 631800
rect 550200 631600 550400 631800
rect 550600 631600 550800 631800
rect 551000 631600 551200 631800
rect 551400 631600 551600 631800
rect 551800 631600 552000 631800
rect 552200 631600 552400 631800
rect 552600 631600 552800 631800
rect 553000 631600 584800 631800
rect 549600 631400 584800 631600
rect 549600 631200 550000 631400
rect 550200 631200 550400 631400
rect 550600 631200 550800 631400
rect 551000 631200 551200 631400
rect 551400 631200 551600 631400
rect 551800 631200 552000 631400
rect 552200 631200 552400 631400
rect 552600 631200 552800 631400
rect 553000 631200 584800 631400
rect 549600 631000 584800 631200
rect 549600 630800 550000 631000
rect 550200 630800 550400 631000
rect 550600 630800 550800 631000
rect 551000 630800 551200 631000
rect 551400 630800 551600 631000
rect 551800 630800 552000 631000
rect 552200 630800 552400 631000
rect 552600 630800 552800 631000
rect 553000 630800 584800 631000
rect 549600 630700 584800 630800
rect 549600 630500 550000 630700
rect 550200 630500 550400 630700
rect 550600 630500 550800 630700
rect 551000 630500 551200 630700
rect 551400 630500 551600 630700
rect 551800 630500 552000 630700
rect 552200 630500 552400 630700
rect 552600 630500 552800 630700
rect 553000 630500 584800 630700
rect 549600 630400 584800 630500
rect 549600 630200 550000 630400
rect 550200 630200 550400 630400
rect 550600 630200 550800 630400
rect 551000 630200 551200 630400
rect 551400 630200 551600 630400
rect 551800 630200 552000 630400
rect 552200 630200 552400 630400
rect 552600 630200 552800 630400
rect 553000 630200 584800 630400
rect 549600 630000 584800 630200
rect 549600 629800 550000 630000
rect 550200 629800 550400 630000
rect 550600 629800 550800 630000
rect 551000 629800 551200 630000
rect 551400 629800 551600 630000
rect 551800 629800 552000 630000
rect 552200 629800 552400 630000
rect 552600 629800 552800 630000
rect 553000 629800 584800 630000
rect 549600 629784 584800 629800
rect 549600 629400 584000 629784
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 282000 583800 584000 584200
rect 282000 583400 282400 583800
rect 282800 583400 283200 583800
rect 283600 583674 584000 583800
rect 283600 583562 584800 583674
rect 283600 583400 584000 583562
rect 282000 583000 584000 583400
rect 282000 582600 282400 583000
rect 282800 582600 283200 583000
rect 283600 582600 584000 583000
rect 282000 582200 584000 582600
rect 282000 581800 282400 582200
rect 282800 581800 283200 582200
rect 283600 581800 584000 582200
rect 282000 581400 584000 581800
rect 282000 581000 282400 581400
rect 282800 581000 283200 581400
rect 283600 581000 584000 581400
rect 282000 580600 584000 581000
rect 282000 580200 282400 580600
rect 282800 580200 283200 580600
rect 283600 580200 584000 580600
rect 282000 579800 584000 580200
rect 282000 579400 282400 579800
rect 282800 579400 283200 579800
rect 283600 579400 584000 579800
rect 282000 579000 584000 579400
rect 0 564242 12020 564300
rect -800 559442 12020 564242
rect 0 554242 12020 559442
rect -800 549442 12020 554242
rect 0 549400 12020 549442
rect 12540 564100 40800 564300
rect 12540 563900 32800 564100
rect 33000 563900 33200 564100
rect 33400 563900 33600 564100
rect 33800 563900 34000 564100
rect 34200 563900 34400 564100
rect 34600 563900 34800 564100
rect 35000 563900 35200 564100
rect 35400 563900 35600 564100
rect 35800 563900 36000 564100
rect 36200 563900 36400 564100
rect 36600 563900 36800 564100
rect 37000 563900 37200 564100
rect 37400 563900 37600 564100
rect 37800 563900 38000 564100
rect 38200 563900 38400 564100
rect 38600 563900 38800 564100
rect 39000 563900 39200 564100
rect 39400 563900 39600 564100
rect 39800 563900 40000 564100
rect 40200 563900 40400 564100
rect 40600 563900 40800 564100
rect 12540 563700 40800 563900
rect 12540 563500 32800 563700
rect 33000 563500 33200 563700
rect 33400 563500 33600 563700
rect 33800 563500 34000 563700
rect 34200 563500 34400 563700
rect 34600 563500 34800 563700
rect 35000 563500 35200 563700
rect 35400 563500 35600 563700
rect 35800 563500 36000 563700
rect 36200 563500 36400 563700
rect 36600 563500 36800 563700
rect 37000 563500 37200 563700
rect 37400 563500 37600 563700
rect 37800 563500 38000 563700
rect 38200 563500 38400 563700
rect 38600 563500 38800 563700
rect 39000 563500 39200 563700
rect 39400 563500 39600 563700
rect 39800 563500 40000 563700
rect 40200 563500 40400 563700
rect 40600 563500 40800 563700
rect 12540 563300 40800 563500
rect 12540 563100 32800 563300
rect 33000 563100 33200 563300
rect 33400 563100 33600 563300
rect 33800 563100 34000 563300
rect 34200 563100 34400 563300
rect 34600 563100 34800 563300
rect 35000 563100 35200 563300
rect 35400 563100 35600 563300
rect 35800 563100 36000 563300
rect 36200 563100 36400 563300
rect 36600 563100 36800 563300
rect 37000 563100 37200 563300
rect 37400 563100 37600 563300
rect 37800 563100 38000 563300
rect 38200 563100 38400 563300
rect 38600 563100 38800 563300
rect 39000 563100 39200 563300
rect 39400 563100 39600 563300
rect 39800 563100 40000 563300
rect 40200 563100 40400 563300
rect 40600 563220 40800 563300
rect 40600 563100 40760 563220
rect 12540 563060 40760 563100
rect 12540 562900 40800 563060
rect 12540 562700 32800 562900
rect 33000 562700 33200 562900
rect 33400 562700 33600 562900
rect 33800 562700 34000 562900
rect 34200 562700 34400 562900
rect 34600 562700 34800 562900
rect 35000 562700 35200 562900
rect 35400 562700 35600 562900
rect 35800 562700 36000 562900
rect 36200 562700 36400 562900
rect 36600 562700 36800 562900
rect 37000 562700 37200 562900
rect 37400 562700 37600 562900
rect 37800 562700 38000 562900
rect 38200 562700 38400 562900
rect 38600 562700 38800 562900
rect 39000 562700 39200 562900
rect 39400 562700 39600 562900
rect 39800 562700 40000 562900
rect 40200 562700 40400 562900
rect 40600 562700 40800 562900
rect 12540 562500 40800 562700
rect 12540 562300 32800 562500
rect 33000 562300 33200 562500
rect 33400 562300 33600 562500
rect 33800 562300 34000 562500
rect 34200 562300 34400 562500
rect 34600 562300 34800 562500
rect 35000 562300 35200 562500
rect 35400 562300 35600 562500
rect 35800 562300 36000 562500
rect 36200 562300 36400 562500
rect 36600 562300 36800 562500
rect 37000 562300 37200 562500
rect 37400 562300 37600 562500
rect 37800 562300 38000 562500
rect 38200 562300 38400 562500
rect 38600 562300 38800 562500
rect 39000 562300 39200 562500
rect 39400 562300 39600 562500
rect 39800 562300 40000 562500
rect 40200 562300 40400 562500
rect 40600 562300 40800 562500
rect 12540 562100 40800 562300
rect 12540 561900 32800 562100
rect 33000 561900 33200 562100
rect 33400 561900 33600 562100
rect 33800 561900 34000 562100
rect 34200 561900 34400 562100
rect 34600 561900 34800 562100
rect 35000 561900 35200 562100
rect 35400 561900 35600 562100
rect 35800 561900 36000 562100
rect 36200 561900 36400 562100
rect 36600 561900 36800 562100
rect 37000 561900 37200 562100
rect 37400 561900 37600 562100
rect 37800 561900 38000 562100
rect 38200 561900 38400 562100
rect 38600 561900 38800 562100
rect 39000 561900 39200 562100
rect 39400 561900 39600 562100
rect 39800 561900 40000 562100
rect 40200 561900 40400 562100
rect 40600 561900 40800 562100
rect 12540 561700 40800 561900
rect 12540 561500 32800 561700
rect 33000 561500 33200 561700
rect 33400 561500 33600 561700
rect 33800 561500 34000 561700
rect 34200 561500 34400 561700
rect 34600 561500 34800 561700
rect 35000 561500 35200 561700
rect 35400 561500 35600 561700
rect 35800 561500 36000 561700
rect 36200 561500 36400 561700
rect 36600 561500 36800 561700
rect 37000 561500 37200 561700
rect 37400 561500 37600 561700
rect 37800 561500 38000 561700
rect 38200 561500 38400 561700
rect 38600 561500 38800 561700
rect 39000 561500 39200 561700
rect 39400 561500 39600 561700
rect 39800 561500 40000 561700
rect 40200 561500 40400 561700
rect 40600 561500 40800 561700
rect 12540 561300 40800 561500
rect 12540 561100 32800 561300
rect 33000 561100 33200 561300
rect 33400 561100 33600 561300
rect 33800 561100 34000 561300
rect 34200 561100 34400 561300
rect 34600 561100 34800 561300
rect 35000 561100 35200 561300
rect 35400 561100 35600 561300
rect 35800 561100 36000 561300
rect 36200 561100 36400 561300
rect 36600 561100 36800 561300
rect 37000 561100 37200 561300
rect 37400 561100 37600 561300
rect 37800 561100 38000 561300
rect 38200 561100 38400 561300
rect 38600 561100 38800 561300
rect 39000 561100 39200 561300
rect 39400 561100 39600 561300
rect 39800 561100 40000 561300
rect 40200 561100 40400 561300
rect 40600 561100 40800 561300
rect 12540 560900 40800 561100
rect 12540 560700 32800 560900
rect 33000 560700 33200 560900
rect 33400 560700 33600 560900
rect 33800 560700 34000 560900
rect 34200 560700 34400 560900
rect 34600 560700 34800 560900
rect 35000 560700 35200 560900
rect 35400 560700 35600 560900
rect 35800 560700 36000 560900
rect 36200 560700 36400 560900
rect 36600 560700 36800 560900
rect 37000 560700 37200 560900
rect 37400 560700 37600 560900
rect 37800 560700 38000 560900
rect 38200 560700 38400 560900
rect 38600 560700 38800 560900
rect 39000 560700 39200 560900
rect 39400 560700 39600 560900
rect 39800 560700 40000 560900
rect 40200 560700 40400 560900
rect 40600 560700 40800 560900
rect 12540 560500 40800 560700
rect 12540 560300 32800 560500
rect 33000 560300 33200 560500
rect 33400 560300 33600 560500
rect 33800 560300 34000 560500
rect 34200 560300 34400 560500
rect 34600 560300 34800 560500
rect 35000 560300 35200 560500
rect 35400 560300 35600 560500
rect 35800 560300 36000 560500
rect 36200 560300 36400 560500
rect 36600 560300 36800 560500
rect 37000 560300 37200 560500
rect 37400 560300 37600 560500
rect 37800 560300 38000 560500
rect 38200 560300 38400 560500
rect 38600 560300 38800 560500
rect 39000 560300 39200 560500
rect 39400 560300 39600 560500
rect 39800 560300 40000 560500
rect 40200 560300 40400 560500
rect 40600 560300 40800 560500
rect 12540 560100 40800 560300
rect 12540 559900 32800 560100
rect 33000 559900 33200 560100
rect 33400 559900 33600 560100
rect 33800 559900 34000 560100
rect 34200 559900 34400 560100
rect 34600 559900 34800 560100
rect 35000 559900 35200 560100
rect 35400 559900 35600 560100
rect 35800 559900 36000 560100
rect 36200 559900 36400 560100
rect 36600 559900 36800 560100
rect 37000 559900 37200 560100
rect 37400 559900 37600 560100
rect 37800 559900 38000 560100
rect 38200 559900 38400 560100
rect 38600 559900 38800 560100
rect 39000 559900 39200 560100
rect 39400 559900 39600 560100
rect 39800 559900 40000 560100
rect 40200 559900 40400 560100
rect 40600 559900 40800 560100
rect 12540 559700 40800 559900
rect 12540 559500 32800 559700
rect 33000 559500 33200 559700
rect 33400 559500 33600 559700
rect 33800 559500 34000 559700
rect 34200 559500 34400 559700
rect 34600 559500 34800 559700
rect 35000 559500 35200 559700
rect 35400 559500 35600 559700
rect 35800 559500 36000 559700
rect 36200 559500 36400 559700
rect 36600 559500 36800 559700
rect 37000 559500 37200 559700
rect 37400 559500 37600 559700
rect 37800 559500 38000 559700
rect 38200 559500 38400 559700
rect 38600 559500 38800 559700
rect 39000 559500 39200 559700
rect 39400 559500 39600 559700
rect 39800 559500 40000 559700
rect 40200 559500 40400 559700
rect 40600 559500 40800 559700
rect 12540 559300 40800 559500
rect 12540 559100 32800 559300
rect 33000 559100 33200 559300
rect 33400 559100 33600 559300
rect 33800 559100 34000 559300
rect 34200 559100 34400 559300
rect 34600 559100 34800 559300
rect 35000 559100 35200 559300
rect 35400 559100 35600 559300
rect 35800 559100 36000 559300
rect 36200 559100 36400 559300
rect 36600 559100 36800 559300
rect 37000 559100 37200 559300
rect 37400 559100 37600 559300
rect 37800 559100 38000 559300
rect 38200 559100 38400 559300
rect 38600 559100 38800 559300
rect 39000 559100 39200 559300
rect 39400 559100 39600 559300
rect 39800 559100 40000 559300
rect 40200 559100 40400 559300
rect 40600 559100 40800 559300
rect 12540 558900 40800 559100
rect 12540 558700 32800 558900
rect 33000 558700 33200 558900
rect 33400 558700 33600 558900
rect 33800 558700 34000 558900
rect 34200 558700 34400 558900
rect 34600 558700 34800 558900
rect 35000 558700 35200 558900
rect 35400 558700 35600 558900
rect 35800 558700 36000 558900
rect 36200 558700 36400 558900
rect 36600 558700 36800 558900
rect 37000 558700 37200 558900
rect 37400 558700 37600 558900
rect 37800 558700 38000 558900
rect 38200 558700 38400 558900
rect 38600 558700 38800 558900
rect 39000 558700 39200 558900
rect 39400 558700 39600 558900
rect 39800 558700 40000 558900
rect 40200 558700 40400 558900
rect 40600 558700 40800 558900
rect 12540 558500 40800 558700
rect 12540 558300 32800 558500
rect 33000 558300 33200 558500
rect 33400 558300 33600 558500
rect 33800 558300 34000 558500
rect 34200 558300 34400 558500
rect 34600 558300 34800 558500
rect 35000 558300 35200 558500
rect 35400 558300 35600 558500
rect 35800 558300 36000 558500
rect 36200 558300 36400 558500
rect 36600 558300 36800 558500
rect 37000 558300 37200 558500
rect 37400 558300 37600 558500
rect 37800 558300 38000 558500
rect 38200 558300 38400 558500
rect 38600 558300 38800 558500
rect 39000 558300 39200 558500
rect 39400 558300 39600 558500
rect 39800 558300 40000 558500
rect 40200 558300 40400 558500
rect 40600 558300 40800 558500
rect 12540 558100 40800 558300
rect 12540 557900 32800 558100
rect 33000 557900 33200 558100
rect 33400 557900 33600 558100
rect 33800 557900 34000 558100
rect 34200 557900 34400 558100
rect 34600 557900 34800 558100
rect 35000 557900 35200 558100
rect 35400 557900 35600 558100
rect 35800 557900 36000 558100
rect 36200 557900 36400 558100
rect 36600 557900 36800 558100
rect 37000 557900 37200 558100
rect 37400 557900 37600 558100
rect 37800 557900 38000 558100
rect 38200 557900 38400 558100
rect 38600 557900 38800 558100
rect 39000 557900 39200 558100
rect 39400 557900 39600 558100
rect 39800 557900 40000 558100
rect 40200 557900 40400 558100
rect 40600 557900 40800 558100
rect 12540 557700 40800 557900
rect 12540 557500 32800 557700
rect 33000 557500 33200 557700
rect 33400 557500 33600 557700
rect 33800 557500 34000 557700
rect 34200 557500 34400 557700
rect 34600 557500 34800 557700
rect 35000 557500 35200 557700
rect 35400 557500 35600 557700
rect 35800 557500 36000 557700
rect 36200 557500 36400 557700
rect 36600 557500 36800 557700
rect 37000 557500 37200 557700
rect 37400 557500 37600 557700
rect 37800 557500 38000 557700
rect 38200 557500 38400 557700
rect 38600 557500 38800 557700
rect 39000 557500 39200 557700
rect 39400 557500 39600 557700
rect 39800 557500 40000 557700
rect 40200 557500 40400 557700
rect 40600 557500 40800 557700
rect 12540 557300 40800 557500
rect 12540 557100 32800 557300
rect 33000 557100 33200 557300
rect 33400 557100 33600 557300
rect 33800 557100 34000 557300
rect 34200 557100 34400 557300
rect 34600 557100 34800 557300
rect 35000 557100 35200 557300
rect 35400 557100 35600 557300
rect 35800 557100 36000 557300
rect 36200 557100 36400 557300
rect 36600 557100 36800 557300
rect 37000 557100 37200 557300
rect 37400 557100 37600 557300
rect 37800 557100 38000 557300
rect 38200 557100 38400 557300
rect 38600 557100 38800 557300
rect 39000 557100 39200 557300
rect 39400 557100 39600 557300
rect 39800 557100 40000 557300
rect 40200 557100 40400 557300
rect 40600 557100 40800 557300
rect 12540 556900 40800 557100
rect 12540 556700 32800 556900
rect 33000 556700 33200 556900
rect 33400 556700 33600 556900
rect 33800 556700 34000 556900
rect 34200 556700 34400 556900
rect 34600 556700 34800 556900
rect 35000 556700 35200 556900
rect 35400 556700 35600 556900
rect 35800 556700 36000 556900
rect 36200 556700 36400 556900
rect 36600 556700 36800 556900
rect 37000 556700 37200 556900
rect 37400 556700 37600 556900
rect 37800 556700 38000 556900
rect 38200 556700 38400 556900
rect 38600 556700 38800 556900
rect 39000 556700 39200 556900
rect 39400 556700 39600 556900
rect 39800 556700 40000 556900
rect 40200 556700 40400 556900
rect 40600 556700 40800 556900
rect 12540 556500 40800 556700
rect 12540 556300 32800 556500
rect 33000 556300 33200 556500
rect 33400 556300 33600 556500
rect 33800 556300 34000 556500
rect 34200 556300 34400 556500
rect 34600 556300 34800 556500
rect 35000 556300 35200 556500
rect 35400 556300 35600 556500
rect 35800 556300 36000 556500
rect 36200 556300 36400 556500
rect 36600 556300 36800 556500
rect 37000 556300 37200 556500
rect 37400 556300 37600 556500
rect 37800 556300 38000 556500
rect 38200 556300 38400 556500
rect 38600 556300 38800 556500
rect 39000 556300 39200 556500
rect 39400 556300 39600 556500
rect 39800 556300 40000 556500
rect 40200 556300 40400 556500
rect 40600 556300 40800 556500
rect 12540 556100 40800 556300
rect 12540 555900 32800 556100
rect 33000 555900 33200 556100
rect 33400 555900 33600 556100
rect 33800 555900 34000 556100
rect 34200 555900 34400 556100
rect 34600 555900 34800 556100
rect 35000 555900 35200 556100
rect 35400 555900 35600 556100
rect 35800 555900 36000 556100
rect 36200 555900 36400 556100
rect 36600 555900 36800 556100
rect 37000 555900 37200 556100
rect 37400 555900 37600 556100
rect 37800 555900 38000 556100
rect 38200 555900 38400 556100
rect 38600 555900 38800 556100
rect 39000 555900 39200 556100
rect 39400 555900 39600 556100
rect 39800 555900 40000 556100
rect 40200 555900 40400 556100
rect 40600 555900 40800 556100
rect 12540 555700 40800 555900
rect 12540 555500 32800 555700
rect 33000 555500 33200 555700
rect 33400 555500 33600 555700
rect 33800 555500 34000 555700
rect 34200 555500 34400 555700
rect 34600 555500 34800 555700
rect 35000 555500 35200 555700
rect 35400 555500 35600 555700
rect 35800 555500 36000 555700
rect 36200 555500 36400 555700
rect 36600 555500 36800 555700
rect 37000 555500 37200 555700
rect 37400 555500 37600 555700
rect 37800 555500 38000 555700
rect 38200 555500 38400 555700
rect 38600 555500 38800 555700
rect 39000 555500 39200 555700
rect 39400 555500 39600 555700
rect 39800 555500 40000 555700
rect 40200 555500 40400 555700
rect 40600 555500 40800 555700
rect 12540 555300 40800 555500
rect 12540 555100 32800 555300
rect 33000 555100 33200 555300
rect 33400 555100 33600 555300
rect 33800 555100 34000 555300
rect 34200 555100 34400 555300
rect 34600 555100 34800 555300
rect 35000 555100 35200 555300
rect 35400 555100 35600 555300
rect 35800 555100 36000 555300
rect 36200 555100 36400 555300
rect 36600 555100 36800 555300
rect 37000 555100 37200 555300
rect 37400 555100 37600 555300
rect 37800 555100 38000 555300
rect 38200 555100 38400 555300
rect 38600 555100 38800 555300
rect 39000 555100 39200 555300
rect 39400 555100 39600 555300
rect 39800 555100 40000 555300
rect 40200 555100 40400 555300
rect 40600 555100 40800 555300
rect 12540 554900 40800 555100
rect 12540 554700 32800 554900
rect 33000 554700 33200 554900
rect 33400 554700 33600 554900
rect 33800 554700 34000 554900
rect 34200 554700 34400 554900
rect 34600 554700 34800 554900
rect 35000 554700 35200 554900
rect 35400 554700 35600 554900
rect 35800 554700 36000 554900
rect 36200 554700 36400 554900
rect 36600 554700 36800 554900
rect 37000 554700 37200 554900
rect 37400 554700 37600 554900
rect 37800 554700 38000 554900
rect 38200 554700 38400 554900
rect 38600 554700 38800 554900
rect 39000 554700 39200 554900
rect 39400 554700 39600 554900
rect 39800 554700 40000 554900
rect 40200 554700 40400 554900
rect 40600 554700 40800 554900
rect 12540 554500 40800 554700
rect 12540 554300 32800 554500
rect 33000 554300 33200 554500
rect 33400 554300 33600 554500
rect 33800 554300 34000 554500
rect 34200 554300 34400 554500
rect 34600 554300 34800 554500
rect 35000 554300 35200 554500
rect 35400 554300 35600 554500
rect 35800 554300 36000 554500
rect 36200 554300 36400 554500
rect 36600 554300 36800 554500
rect 37000 554300 37200 554500
rect 37400 554300 37600 554500
rect 37800 554300 38000 554500
rect 38200 554300 38400 554500
rect 38600 554300 38800 554500
rect 39000 554300 39200 554500
rect 39400 554300 39600 554500
rect 39800 554300 40000 554500
rect 40200 554300 40400 554500
rect 40600 554300 40800 554500
rect 12540 554100 40800 554300
rect 12540 553900 32800 554100
rect 33000 553900 33200 554100
rect 33400 553900 33600 554100
rect 33800 553900 34000 554100
rect 34200 553900 34400 554100
rect 34600 553900 34800 554100
rect 35000 553900 35200 554100
rect 35400 553900 35600 554100
rect 35800 553900 36000 554100
rect 36200 553900 36400 554100
rect 36600 553900 36800 554100
rect 37000 553900 37200 554100
rect 37400 553900 37600 554100
rect 37800 553900 38000 554100
rect 38200 553900 38400 554100
rect 38600 553900 38800 554100
rect 39000 553900 39200 554100
rect 39400 553900 39600 554100
rect 39800 553900 40000 554100
rect 40200 553900 40400 554100
rect 40600 553900 40800 554100
rect 12540 553700 40800 553900
rect 12540 553500 32800 553700
rect 33000 553500 33200 553700
rect 33400 553500 33600 553700
rect 33800 553500 34000 553700
rect 34200 553500 34400 553700
rect 34600 553500 34800 553700
rect 35000 553500 35200 553700
rect 35400 553500 35600 553700
rect 35800 553500 36000 553700
rect 36200 553500 36400 553700
rect 36600 553500 36800 553700
rect 37000 553500 37200 553700
rect 37400 553500 37600 553700
rect 37800 553500 38000 553700
rect 38200 553500 38400 553700
rect 38600 553500 38800 553700
rect 39000 553500 39200 553700
rect 39400 553500 39600 553700
rect 39800 553500 40000 553700
rect 40200 553500 40400 553700
rect 40600 553500 40800 553700
rect 12540 553300 40800 553500
rect 12540 553100 32800 553300
rect 33000 553100 33200 553300
rect 33400 553100 33600 553300
rect 33800 553100 34000 553300
rect 34200 553100 34400 553300
rect 34600 553100 34800 553300
rect 35000 553100 35200 553300
rect 35400 553100 35600 553300
rect 35800 553100 36000 553300
rect 36200 553100 36400 553300
rect 36600 553100 36800 553300
rect 37000 553100 37200 553300
rect 37400 553100 37600 553300
rect 37800 553100 38000 553300
rect 38200 553100 38400 553300
rect 38600 553100 38800 553300
rect 39000 553100 39200 553300
rect 39400 553100 39600 553300
rect 39800 553100 40000 553300
rect 40200 553100 40400 553300
rect 40600 553100 40800 553300
rect 12540 552900 40800 553100
rect 12540 552700 32800 552900
rect 33000 552700 33200 552900
rect 33400 552700 33600 552900
rect 33800 552700 34000 552900
rect 34200 552700 34400 552900
rect 34600 552700 34800 552900
rect 35000 552700 35200 552900
rect 35400 552700 35600 552900
rect 35800 552700 36000 552900
rect 36200 552700 36400 552900
rect 36600 552700 36800 552900
rect 37000 552700 37200 552900
rect 37400 552700 37600 552900
rect 37800 552700 38000 552900
rect 38200 552700 38400 552900
rect 38600 552700 38800 552900
rect 39000 552700 39200 552900
rect 39400 552700 39600 552900
rect 39800 552700 40000 552900
rect 40200 552700 40400 552900
rect 40600 552700 40800 552900
rect 12540 552500 40800 552700
rect 12540 552300 32800 552500
rect 33000 552300 33200 552500
rect 33400 552300 33600 552500
rect 33800 552300 34000 552500
rect 34200 552300 34400 552500
rect 34600 552300 34800 552500
rect 35000 552300 35200 552500
rect 35400 552300 35600 552500
rect 35800 552300 36000 552500
rect 36200 552300 36400 552500
rect 36600 552300 36800 552500
rect 37000 552300 37200 552500
rect 37400 552300 37600 552500
rect 37800 552300 38000 552500
rect 38200 552300 38400 552500
rect 38600 552300 38800 552500
rect 39000 552300 39200 552500
rect 39400 552300 39600 552500
rect 39800 552300 40000 552500
rect 40200 552300 40400 552500
rect 40600 552300 40800 552500
rect 12540 552100 40800 552300
rect 12540 551900 32800 552100
rect 33000 551900 33200 552100
rect 33400 551900 33600 552100
rect 33800 551900 34000 552100
rect 34200 551900 34400 552100
rect 34600 551900 34800 552100
rect 35000 551900 35200 552100
rect 35400 551900 35600 552100
rect 35800 551900 36000 552100
rect 36200 551900 36400 552100
rect 36600 551900 36800 552100
rect 37000 551900 37200 552100
rect 37400 551900 37600 552100
rect 37800 551900 38000 552100
rect 38200 551900 38400 552100
rect 38600 551900 38800 552100
rect 39000 551900 39200 552100
rect 39400 551900 39600 552100
rect 39800 551900 40000 552100
rect 40200 551900 40400 552100
rect 40600 551900 40800 552100
rect 12540 551700 40800 551900
rect 12540 551500 32800 551700
rect 33000 551500 33200 551700
rect 33400 551500 33600 551700
rect 33800 551500 34000 551700
rect 34200 551500 34400 551700
rect 34600 551500 34800 551700
rect 35000 551500 35200 551700
rect 35400 551500 35600 551700
rect 35800 551500 36000 551700
rect 36200 551500 36400 551700
rect 36600 551500 36800 551700
rect 37000 551500 37200 551700
rect 37400 551500 37600 551700
rect 37800 551500 38000 551700
rect 38200 551500 38400 551700
rect 38600 551500 38800 551700
rect 39000 551500 39200 551700
rect 39400 551500 39600 551700
rect 39800 551500 40000 551700
rect 40200 551500 40400 551700
rect 40600 551500 40800 551700
rect 12540 551300 40800 551500
rect 12540 551100 32800 551300
rect 33000 551100 33200 551300
rect 33400 551100 33600 551300
rect 33800 551100 34000 551300
rect 34200 551100 34400 551300
rect 34600 551100 34800 551300
rect 35000 551100 35200 551300
rect 35400 551100 35600 551300
rect 35800 551100 36000 551300
rect 36200 551100 36400 551300
rect 36600 551100 36800 551300
rect 37000 551100 37200 551300
rect 37400 551100 37600 551300
rect 37800 551100 38000 551300
rect 38200 551100 38400 551300
rect 38600 551100 38800 551300
rect 39000 551100 39200 551300
rect 39400 551100 39600 551300
rect 39800 551100 40000 551300
rect 40200 551100 40400 551300
rect 40600 551100 40800 551300
rect 12540 550900 40800 551100
rect 12540 550700 32800 550900
rect 33000 550700 33200 550900
rect 33400 550700 33600 550900
rect 33800 550700 34000 550900
rect 34200 550700 34400 550900
rect 34600 550700 34800 550900
rect 35000 550700 35200 550900
rect 35400 550700 35600 550900
rect 35800 550700 36000 550900
rect 36200 550700 36400 550900
rect 36600 550700 36800 550900
rect 37000 550700 37200 550900
rect 37400 550700 37600 550900
rect 37800 550700 38000 550900
rect 38200 550700 38400 550900
rect 38600 550700 38800 550900
rect 39000 550700 39200 550900
rect 39400 550700 39600 550900
rect 39800 550700 40000 550900
rect 40200 550700 40400 550900
rect 40600 550700 40800 550900
rect 12540 550500 40800 550700
rect 582340 550562 584800 555362
rect 12540 550300 32800 550500
rect 33000 550300 33200 550500
rect 33400 550300 33600 550500
rect 33800 550300 34000 550500
rect 34200 550300 34400 550500
rect 34600 550300 34800 550500
rect 35000 550300 35200 550500
rect 35400 550300 35600 550500
rect 35800 550300 36000 550500
rect 36200 550300 36400 550500
rect 36600 550300 36800 550500
rect 37000 550300 37200 550500
rect 37400 550300 37600 550500
rect 37800 550300 38000 550500
rect 38200 550300 38400 550500
rect 38600 550300 38800 550500
rect 39000 550300 39200 550500
rect 39400 550300 39600 550500
rect 39800 550300 40000 550500
rect 40200 550300 40400 550500
rect 40600 550300 40800 550500
rect 12540 550100 40800 550300
rect 12540 549900 32800 550100
rect 33000 549900 33200 550100
rect 33400 549900 33600 550100
rect 33800 549900 34000 550100
rect 34200 549900 34400 550100
rect 34600 549900 34800 550100
rect 35000 549900 35200 550100
rect 35400 549900 35600 550100
rect 35800 549900 36000 550100
rect 36200 549900 36400 550100
rect 36600 549900 36800 550100
rect 37000 549900 37200 550100
rect 37400 549900 37600 550100
rect 37800 549900 38000 550100
rect 38200 549900 38400 550100
rect 38600 549900 38800 550100
rect 39000 549900 39200 550100
rect 39400 549900 39600 550100
rect 39800 549900 40000 550100
rect 40200 549900 40400 550100
rect 40600 549900 40800 550100
rect 12540 549700 40800 549900
rect 12540 549500 32800 549700
rect 33000 549500 33200 549700
rect 33400 549500 33600 549700
rect 33800 549500 34000 549700
rect 34200 549500 34400 549700
rect 34600 549500 34800 549700
rect 35000 549500 35200 549700
rect 35400 549500 35600 549700
rect 35800 549500 36000 549700
rect 36200 549500 36400 549700
rect 36600 549500 36800 549700
rect 37000 549500 37200 549700
rect 37400 549500 37600 549700
rect 37800 549500 38000 549700
rect 38200 549500 38400 549700
rect 38600 549500 38800 549700
rect 39000 549500 39200 549700
rect 39400 549500 39600 549700
rect 39800 549500 40000 549700
rect 40200 549500 40400 549700
rect 40600 549500 40800 549700
rect 12540 549400 40800 549500
rect 582340 540562 584800 545362
rect 0 511642 277400 516200
rect -800 511530 277400 511642
rect 0 511000 277400 511530
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 0 468420 271200 473000
rect -800 468308 271200 468420
rect 0 467800 271200 468308
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 0 425198 265000 429600
rect -800 425086 265000 425198
rect 0 424400 265000 425086
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 0 381976 258800 386600
rect -800 381864 258800 381976
rect 0 381400 258800 381864
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 253600 347800 258800 381400
rect 259800 349500 265000 424400
rect 266000 351200 271200 467800
rect 272200 352700 277400 511000
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 285000 494252 584000 494600
rect 285000 494200 584800 494252
rect 285000 493800 285400 494200
rect 285800 493800 286200 494200
rect 286600 494140 584800 494200
rect 286600 493800 584000 494140
rect 285000 493400 584000 493800
rect 285000 493000 285400 493400
rect 285800 493000 286200 493400
rect 286600 493000 584000 493400
rect 285000 492600 584000 493000
rect 285000 492200 285400 492600
rect 285800 492200 286200 492600
rect 286600 492200 584000 492600
rect 285000 491800 584000 492200
rect 285000 491400 285400 491800
rect 285800 491400 286200 491800
rect 286600 491400 584000 491800
rect 285000 491000 584000 491400
rect 285000 490600 285400 491000
rect 285800 490600 286200 491000
rect 286600 490600 584000 491000
rect 285000 490200 584000 490600
rect 285000 489800 285400 490200
rect 285800 489800 286200 490200
rect 286600 489800 584000 490200
rect 285000 489400 584000 489800
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 288000 449830 584000 450100
rect 288000 449800 584800 449830
rect 288000 449400 288400 449800
rect 288800 449400 289200 449800
rect 289600 449718 584800 449800
rect 289600 449400 584000 449718
rect 288000 449000 584000 449400
rect 288000 448600 288400 449000
rect 288800 448600 289200 449000
rect 289600 448600 584000 449000
rect 288000 448200 584000 448600
rect 288000 447800 288400 448200
rect 288800 447800 289200 448200
rect 289600 447800 584000 448200
rect 288000 447400 584000 447800
rect 288000 447000 288400 447400
rect 288800 447000 289200 447400
rect 289600 447000 584000 447400
rect 288000 446600 584000 447000
rect 288000 446200 288400 446600
rect 288800 446200 289200 446600
rect 289600 446200 584000 446600
rect 288000 445800 584000 446200
rect 288000 445400 288400 445800
rect 288800 445400 289200 445800
rect 289600 445400 584000 445800
rect 288000 444900 584000 445400
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 291100 405408 584000 405700
rect 291100 405400 584800 405408
rect 291100 405000 291400 405400
rect 291800 405000 292200 405400
rect 292600 405296 584800 405400
rect 292600 405000 584000 405296
rect 291100 404600 584000 405000
rect 291100 404200 291400 404600
rect 291800 404200 292200 404600
rect 292600 404200 584000 404600
rect 291100 403800 584000 404200
rect 291100 403400 291400 403800
rect 291800 403400 292200 403800
rect 292600 403400 584000 403800
rect 291100 403000 584000 403400
rect 291100 402600 291400 403000
rect 291800 402600 292200 403000
rect 292600 402600 584000 403000
rect 291100 402200 584000 402600
rect 291100 401800 291400 402200
rect 291800 401800 292200 402200
rect 292600 401800 584000 402200
rect 291100 401400 584000 401800
rect 291100 401000 291400 401400
rect 291800 401000 292200 401400
rect 292600 401000 584000 401400
rect 291100 400500 584000 401000
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583524 360056 584800 360168
rect 294000 359000 584000 359400
rect 294000 358600 294400 359000
rect 294800 358600 295200 359000
rect 295600 358986 584000 359000
rect 295600 358874 584800 358986
rect 295600 358600 584000 358874
rect 294000 358200 584000 358600
rect 294000 357800 294400 358200
rect 294800 357800 295200 358200
rect 295600 357800 584000 358200
rect 294000 357400 584000 357800
rect 294000 357000 294400 357400
rect 294800 357000 295200 357400
rect 295600 357000 584000 357400
rect 294000 356600 584000 357000
rect 294000 356200 294400 356600
rect 294800 356200 295200 356600
rect 295600 356200 584000 356600
rect 294000 355800 584000 356200
rect 294000 355400 294400 355800
rect 294800 355400 295200 355800
rect 295600 355400 584000 355800
rect 294000 355000 584000 355400
rect 294000 354600 294400 355000
rect 294800 354600 295200 355000
rect 295600 354600 584000 355000
rect 294000 354200 584000 354600
rect 272200 352640 281300 352700
rect 272200 352580 281080 352640
rect 281140 352580 281180 352640
rect 281240 352580 281300 352640
rect 272200 352540 281300 352580
rect 272200 352480 281080 352540
rect 281140 352480 281180 352540
rect 281240 352480 281300 352540
rect 272200 352300 281300 352480
rect 294700 352660 348000 352800
rect 294700 352600 294760 352660
rect 294820 352600 294860 352660
rect 294920 352600 348000 352660
rect 294700 352560 348000 352600
rect 294700 352500 294760 352560
rect 294820 352500 294860 352560
rect 294920 352500 348000 352560
rect 294700 352400 348000 352500
rect 266000 351080 281300 351200
rect 266000 351020 281060 351080
rect 281120 351020 281160 351080
rect 281220 351020 281300 351080
rect 266000 350980 281300 351020
rect 266000 350920 281060 350980
rect 281120 350920 281160 350980
rect 281220 350920 281300 350980
rect 266000 350800 281300 350920
rect 294700 350920 341800 351000
rect 294700 350860 294760 350920
rect 294820 350860 294860 350920
rect 294920 350860 341800 350920
rect 294700 350820 341800 350860
rect 294700 350760 294760 350820
rect 294820 350760 294860 350820
rect 294920 350760 341800 350820
rect 294700 350600 341800 350760
rect 259800 349380 281300 349500
rect 259800 349320 281060 349380
rect 281120 349320 281160 349380
rect 281220 349320 281300 349380
rect 259800 349280 281300 349320
rect 259800 349220 281060 349280
rect 281120 349220 281160 349280
rect 281220 349220 281300 349280
rect 259800 349100 281300 349220
rect 294700 349220 335600 349300
rect 294700 349160 294760 349220
rect 294820 349160 294860 349220
rect 294920 349160 335600 349220
rect 294700 349120 335600 349160
rect 294700 349060 294760 349120
rect 294820 349060 294860 349120
rect 294920 349060 335600 349120
rect 294700 348900 335600 349060
rect 253600 347680 281300 347800
rect 253600 347620 281040 347680
rect 281100 347620 281140 347680
rect 281200 347620 281300 347680
rect 253600 347580 281300 347620
rect 253600 347520 281040 347580
rect 281100 347520 281140 347580
rect 281200 347520 281300 347580
rect 253600 347400 281300 347520
rect 294700 347520 329400 347600
rect 294700 347460 294760 347520
rect 294820 347460 294860 347520
rect 294920 347460 329400 347520
rect 294700 347420 329400 347460
rect 294700 347360 294760 347420
rect 294820 347360 294860 347420
rect 294920 347360 329400 347420
rect 294700 347200 329400 347360
rect 253600 345980 281300 346100
rect 253600 345920 281060 345980
rect 281120 345920 281160 345980
rect 281220 345920 281300 345980
rect 253600 345880 281300 345920
rect 253600 345820 281060 345880
rect 281120 345820 281160 345880
rect 281220 345820 281300 345880
rect 253600 345700 281300 345820
rect 294700 345820 323200 345900
rect 294700 345760 294760 345820
rect 294820 345760 294860 345820
rect 294920 345760 323200 345820
rect 294700 345720 323200 345760
rect 253600 343100 258800 345700
rect 294700 345660 294760 345720
rect 294820 345660 294860 345720
rect 294920 345660 323200 345720
rect 294700 345500 323200 345660
rect 0 338754 258800 343100
rect -800 338642 258800 338754
rect 0 337900 258800 338642
rect 259800 344260 281300 344400
rect 259800 344200 281060 344260
rect 281120 344200 281160 344260
rect 281220 344200 281300 344260
rect 259800 344160 281300 344200
rect 259800 344100 281060 344160
rect 281120 344100 281160 344160
rect 281220 344100 281300 344160
rect 259800 344000 281300 344100
rect 294790 344200 295110 344205
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 9650 304380 11580 304410
rect 9650 304320 9680 304380
rect 9740 304320 9845 304380
rect 9905 304320 10045 304380
rect 10105 304320 10235 304380
rect 10295 304320 10415 304380
rect 10475 304320 10615 304380
rect 10675 304320 10805 304380
rect 10865 304320 10965 304380
rect 11025 304320 11155 304380
rect 11215 304320 11330 304380
rect 11390 304320 11470 304380
rect 11530 304320 11580 304380
rect 9650 304210 11580 304320
rect 9650 304200 11600 304210
rect 9650 304180 9800 304200
rect 10000 304180 10200 304200
rect 10400 304180 10600 304200
rect 10800 304180 11000 304200
rect 11200 304180 11400 304200
rect 9650 304120 9680 304180
rect 9740 304120 9800 304180
rect 10000 304120 10045 304180
rect 10105 304120 10200 304180
rect 10400 304120 10415 304180
rect 10475 304120 10600 304180
rect 10800 304120 10805 304180
rect 10865 304120 10965 304180
rect 11215 304120 11330 304180
rect 11390 304120 11400 304180
rect 9650 304000 9800 304120
rect 10000 304000 10200 304120
rect 10400 304000 10600 304120
rect 10800 304000 11000 304120
rect 11200 304000 11400 304120
rect 9650 303990 11600 304000
rect 9650 303980 11580 303990
rect 9650 303920 9680 303980
rect 9740 303920 9845 303980
rect 9905 303920 10045 303980
rect 10105 303920 10235 303980
rect 10295 303920 10415 303980
rect 10475 303920 10615 303980
rect 10675 303920 10805 303980
rect 10865 303920 10965 303980
rect 11025 303920 11155 303980
rect 11215 303920 11330 303980
rect 11390 303920 11470 303980
rect 11530 303920 11580 303980
rect 9650 303790 11580 303920
rect 9650 303730 9680 303790
rect 9740 303730 9845 303790
rect 9905 303730 10045 303790
rect 10105 303730 10235 303790
rect 10295 303730 10415 303790
rect 10475 303730 10615 303790
rect 10675 303730 10805 303790
rect 10865 303730 10965 303790
rect 11025 303730 11155 303790
rect 11215 303730 11330 303790
rect 11390 303730 11470 303790
rect 11530 303730 11580 303790
rect 9650 303610 11580 303730
rect 9650 303600 11600 303610
rect 9650 303590 9800 303600
rect 10000 303590 10200 303600
rect 10400 303590 10600 303600
rect 10800 303590 11000 303600
rect 11200 303590 11400 303600
rect 9650 303530 9680 303590
rect 9740 303530 9800 303590
rect 10000 303530 10045 303590
rect 10105 303530 10200 303590
rect 10400 303530 10415 303590
rect 10475 303530 10600 303590
rect 10800 303530 10805 303590
rect 10865 303530 10965 303590
rect 11215 303530 11330 303590
rect 11390 303530 11400 303590
rect 9650 303400 9800 303530
rect 10000 303400 10200 303530
rect 10400 303400 10600 303530
rect 10800 303400 11000 303530
rect 11200 303400 11400 303530
rect 9650 303340 9680 303400
rect 9740 303390 11600 303400
rect 9740 303340 9845 303390
rect 9650 303330 9845 303340
rect 9905 303330 10045 303390
rect 10105 303330 10235 303390
rect 10295 303330 10415 303390
rect 10475 303330 10615 303390
rect 10675 303330 10805 303390
rect 10865 303330 10965 303390
rect 11025 303330 11155 303390
rect 11215 303330 11330 303390
rect 11390 303330 11470 303390
rect 11530 303330 11580 303390
rect 9650 303300 11580 303330
rect 14960 303260 15380 303280
rect 14960 303120 15000 303260
rect 15140 303120 15200 303260
rect 15340 303120 15380 303260
rect 5700 301194 8200 301200
rect 4000 301000 8200 301194
rect 4000 300800 5800 301000
rect 6000 300800 6200 301000
rect 6400 300800 6600 301000
rect 6800 300800 7000 301000
rect 7200 300800 7400 301000
rect 7600 300800 7800 301000
rect 8000 300800 8200 301000
rect 4000 300600 8200 300800
rect 4000 300400 5800 300600
rect 6000 300400 6200 300600
rect 6400 300400 6600 300600
rect 6800 300400 7000 300600
rect 7200 300400 7400 300600
rect 7600 300400 7800 300600
rect 8000 300400 8200 300600
rect 4000 300200 8200 300400
rect 4000 300000 5800 300200
rect 6000 300000 6200 300200
rect 6400 300000 6600 300200
rect 6800 300000 7000 300200
rect 7200 300000 7400 300200
rect 7600 300000 7800 300200
rect 8000 300000 8200 300200
rect 4000 299800 8200 300000
rect 4000 299600 5800 299800
rect 6000 299600 6200 299800
rect 6400 299600 6600 299800
rect 6800 299600 7000 299800
rect 7200 299600 7400 299800
rect 7600 299600 7800 299800
rect 8000 299600 8200 299800
rect 4000 299400 8200 299600
rect 4000 299200 5800 299400
rect 6000 299200 6200 299400
rect 6400 299200 6600 299400
rect 6800 299200 7000 299400
rect 7200 299200 7400 299400
rect 7600 299200 7800 299400
rect 8000 299200 8200 299400
rect 4000 299000 8200 299200
rect 4000 298800 5800 299000
rect 6000 298800 6200 299000
rect 6400 298800 6600 299000
rect 6800 298800 7000 299000
rect 7200 298800 7400 299000
rect 7600 298800 7800 299000
rect 8000 298800 8200 299000
rect 4000 298600 8200 298800
rect 4000 298400 5800 298600
rect 6000 298400 6200 298600
rect 6400 298400 6600 298600
rect 6800 298400 7000 298600
rect 7200 298400 7400 298600
rect 7600 298400 7800 298600
rect 8000 298400 8200 298600
rect 4000 298200 8200 298400
rect 4000 298000 5800 298200
rect 6000 298000 6200 298200
rect 6400 298000 6600 298200
rect 6800 298000 7000 298200
rect 7200 298000 7400 298200
rect 7600 298000 7800 298200
rect 8000 298000 8200 298200
rect 4000 297800 8200 298000
rect 4000 297600 5800 297800
rect 6000 297600 6200 297800
rect 6400 297600 6600 297800
rect 6800 297600 7000 297800
rect 7200 297600 7400 297800
rect 7600 297600 7800 297800
rect 8000 297600 8200 297800
rect 4000 297400 8200 297600
rect 4000 297200 5800 297400
rect 6000 297200 6200 297400
rect 6400 297200 6600 297400
rect 6800 297200 7000 297400
rect 7200 297200 7400 297400
rect 7600 297200 7800 297400
rect 8000 297200 8200 297400
rect 4000 297000 8200 297200
rect 4000 296800 5800 297000
rect 6000 296800 6200 297000
rect 6400 296800 6600 297000
rect 6800 296800 7000 297000
rect 7200 296800 7400 297000
rect 7600 296800 7800 297000
rect 8000 296800 8200 297000
rect 4000 296600 8200 296800
rect 4000 296400 5800 296600
rect 6000 296400 6200 296600
rect 6400 296400 6600 296600
rect 6800 296400 7000 296600
rect 7200 296400 7400 296600
rect 7600 296400 7800 296600
rect 8000 296400 8200 296600
rect 4000 296200 8200 296400
rect 0 295532 5700 296200
rect -800 295420 5700 295532
rect 0 295200 5700 295420
rect -800 294238 480 294350
rect 14960 294200 15380 303120
rect 14960 294060 15000 294200
rect 15140 294060 15200 294200
rect 15340 294060 15380 294200
rect 14960 294040 15380 294060
rect 17600 301000 18600 301200
rect 17600 300800 17800 301000
rect 18000 300800 18200 301000
rect 18400 300800 18600 301000
rect 17600 300600 18600 300800
rect 17600 300400 17800 300600
rect 18000 300400 18200 300600
rect 18400 300400 18600 300600
rect 17600 300200 18600 300400
rect 17600 300000 17800 300200
rect 18000 300000 18200 300200
rect 18400 300000 18600 300200
rect 17600 299800 18600 300000
rect 17600 299600 17800 299800
rect 18000 299600 18200 299800
rect 18400 299600 18600 299800
rect 17600 299400 18600 299600
rect 17600 299200 17800 299400
rect 18000 299200 18200 299400
rect 18400 299200 18600 299400
rect 17600 299000 18600 299200
rect 259800 299000 265000 344000
rect 294790 343900 294800 344200
rect 295100 343900 295110 344200
rect 294790 343895 295110 343900
rect 17600 298800 17800 299000
rect 18000 298800 18200 299000
rect 18400 298800 18600 299000
rect 17600 298600 18600 298800
rect 17600 298400 17800 298600
rect 18000 298400 18200 298600
rect 18400 298400 18600 298600
rect 17600 298200 18600 298400
rect 17600 298000 17800 298200
rect 18000 298000 18200 298200
rect 18400 298000 18600 298200
rect 17600 297800 18600 298000
rect 17600 297600 17800 297800
rect 18000 297600 18200 297800
rect 18400 297600 18600 297800
rect 17600 297400 18600 297600
rect 17600 297200 17800 297400
rect 18000 297200 18200 297400
rect 18400 297200 18600 297400
rect 17600 297000 18600 297200
rect 17600 296800 17800 297000
rect 18000 296800 18200 297000
rect 18400 296800 18600 297000
rect 17600 296600 18600 296800
rect 17600 296400 17800 296600
rect 18000 296400 18200 296600
rect 18400 296400 18600 296600
rect 9650 293980 11580 294010
rect 5735 293920 5925 293930
rect 5735 293740 5740 293920
rect 5920 293740 5925 293920
rect 5735 293730 5925 293740
rect 9650 293920 9680 293980
rect 9740 293920 9845 293980
rect 9905 293920 10045 293980
rect 10105 293920 10235 293980
rect 10295 293920 10415 293980
rect 10475 293920 10615 293980
rect 10675 293920 10805 293980
rect 10865 293920 10965 293980
rect 11025 293920 11155 293980
rect 11215 293920 11330 293980
rect 11390 293920 11470 293980
rect 11530 293920 11580 293980
rect 9650 293810 11580 293920
rect 9650 293800 11600 293810
rect 9650 293780 9800 293800
rect 10000 293780 10200 293800
rect 10400 293780 10600 293800
rect 10800 293780 11000 293800
rect 11200 293780 11400 293800
rect 9650 293720 9680 293780
rect 9740 293720 9800 293780
rect 10000 293720 10045 293780
rect 10105 293720 10200 293780
rect 10400 293720 10415 293780
rect 10475 293720 10600 293780
rect 10800 293720 10805 293780
rect 10865 293720 10965 293780
rect 11215 293720 11330 293780
rect 11390 293720 11400 293780
rect 9650 293600 9800 293720
rect 10000 293600 10200 293720
rect 10400 293600 10600 293720
rect 10800 293600 11000 293720
rect 11200 293600 11400 293720
rect 9650 293590 11600 293600
rect 5735 293580 5925 293590
rect 5735 293400 5740 293580
rect 5920 293400 5925 293580
rect 5735 293390 5925 293400
rect 9650 293580 11580 293590
rect 9650 293520 9680 293580
rect 9740 293520 9845 293580
rect 9905 293520 10045 293580
rect 10105 293520 10235 293580
rect 10295 293520 10415 293580
rect 10475 293520 10615 293580
rect 10675 293520 10805 293580
rect 10865 293520 10965 293580
rect 11025 293520 11155 293580
rect 11215 293520 11330 293580
rect 11390 293520 11470 293580
rect 11530 293520 11580 293580
rect 9650 293390 11580 293520
rect 9650 293330 9680 293390
rect 9740 293330 9845 293390
rect 9905 293330 10045 293390
rect 10105 293330 10235 293390
rect 10295 293330 10415 293390
rect 10475 293330 10615 293390
rect 10675 293330 10805 293390
rect 10865 293330 10965 293390
rect 11025 293330 11155 293390
rect 11215 293330 11330 293390
rect 11390 293330 11470 293390
rect 11530 293330 11580 293390
rect 5735 293240 5925 293250
rect -800 293056 480 293168
rect 5735 293060 5740 293240
rect 5920 293060 5925 293240
rect 5735 293050 5925 293060
rect 9650 293210 11580 293330
rect 9650 293200 11600 293210
rect 9650 293190 9800 293200
rect 10000 293190 10200 293200
rect 10400 293190 10600 293200
rect 10800 293190 11000 293200
rect 11200 293190 11400 293200
rect 9650 293130 9680 293190
rect 9740 293130 9800 293190
rect 10000 293130 10045 293190
rect 10105 293130 10200 293190
rect 10400 293130 10415 293190
rect 10475 293130 10600 293190
rect 10800 293130 10805 293190
rect 10865 293130 10965 293190
rect 11215 293130 11330 293190
rect 11390 293130 11400 293190
rect 9650 293000 9800 293130
rect 10000 293000 10200 293130
rect 10400 293000 10600 293130
rect 10800 293000 11000 293130
rect 11200 293000 11400 293130
rect 9650 292940 9680 293000
rect 9740 292990 11600 293000
rect 9740 292940 9845 292990
rect 9650 292930 9845 292940
rect 9905 292930 10045 292990
rect 10105 292930 10235 292990
rect 10295 292930 10415 292990
rect 10475 292930 10615 292990
rect 10675 292930 10805 292990
rect 10865 292930 10965 292990
rect 11025 292930 11155 292990
rect 11215 292930 11330 292990
rect 11390 292930 11470 292990
rect 11530 292930 11580 292990
rect 9650 292900 11580 292930
rect 14960 292860 15380 292880
rect 14960 292720 15000 292860
rect 15140 292720 15200 292860
rect 15340 292720 15380 292860
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 13060 280500 13280 280520
rect 13060 280430 13190 280500
rect 13260 280430 13280 280500
rect 13060 280390 13280 280430
rect 13060 280320 13080 280390
rect 13150 280320 13280 280390
rect 13060 280300 13280 280320
rect 6871 280022 10370 280050
rect 6871 276678 6891 280022
rect 6955 276678 10370 280022
rect 14535 278550 14645 278560
rect 14535 278370 14540 278550
rect 14640 278370 14645 278550
rect 14535 278360 14645 278370
rect 14960 278540 15380 292720
rect 14960 278400 15000 278540
rect 15140 278400 15200 278540
rect 15340 278400 15380 278540
rect 14960 278320 15380 278400
rect 14960 278180 15000 278320
rect 15140 278180 15200 278320
rect 15340 278180 15380 278320
rect 14535 278130 14645 278140
rect 14535 277950 14540 278130
rect 14640 277950 14645 278130
rect 14535 277940 14645 277950
rect 14960 278100 15380 278180
rect 14960 277960 15000 278100
rect 15140 277960 15200 278100
rect 15340 277960 15380 278100
rect 14960 277920 15380 277960
rect 15960 289800 16440 290200
rect 15960 289600 16100 289800
rect 16300 289600 16440 289800
rect 15960 289400 16440 289600
rect 15960 289200 16100 289400
rect 16300 289200 16440 289400
rect 15960 289000 16440 289200
rect 15960 288800 16100 289000
rect 16300 288800 16440 289000
rect 15960 288600 16440 288800
rect 15960 288400 16100 288600
rect 16300 288400 16440 288600
rect 15960 288200 16440 288400
rect 15960 288000 16100 288200
rect 16300 288000 16440 288200
rect 15960 287800 16440 288000
rect 15960 287600 16100 287800
rect 16300 287600 16440 287800
rect 15960 287400 16440 287600
rect 15960 287200 16100 287400
rect 16300 287200 16440 287400
rect 15960 287000 16440 287200
rect 15960 286800 16100 287000
rect 16300 286800 16440 287000
rect 15960 286600 16440 286800
rect 15960 286400 16100 286600
rect 16300 286400 16440 286600
rect 15960 286200 16440 286400
rect 15960 286000 16100 286200
rect 16300 286000 16440 286200
rect 6871 276650 10370 276678
rect 14020 276600 14160 276620
rect 14020 276510 14040 276600
rect 14140 276510 14160 276600
rect 14020 276410 14160 276510
rect 14020 276320 14040 276410
rect 14140 276320 14160 276410
rect 6871 276222 10370 276250
rect 6871 272878 6891 276222
rect 6955 272878 10370 276222
rect 12835 275850 12915 275860
rect 13075 275850 13155 275860
rect 12830 275780 12840 275850
rect 12910 275780 13080 275850
rect 13150 275780 13160 275850
rect 12830 275540 13160 275780
rect 12830 275470 12840 275540
rect 12910 275470 13080 275540
rect 13150 275470 13160 275540
rect 12830 275220 12870 275470
rect 13120 275220 13160 275470
rect 12830 275150 12840 275220
rect 12910 275150 13080 275220
rect 13150 275150 13160 275220
rect 12830 274900 13160 275150
rect 12830 274830 12840 274900
rect 12910 274830 13080 274900
rect 13150 274830 13160 274900
rect 12830 274590 13160 274830
rect 12830 274520 12840 274590
rect 12910 274520 13080 274590
rect 13150 274520 13160 274590
rect 12830 274270 13160 274520
rect 12830 274200 12840 274270
rect 12910 274200 13080 274270
rect 13150 274200 13160 274270
rect 12830 273960 13160 274200
rect 12830 273890 12840 273960
rect 12910 273890 13080 273960
rect 13150 273890 13160 273960
rect 12830 273640 13160 273890
rect 12830 273570 12840 273640
rect 12910 273570 13080 273640
rect 13150 273570 13160 273640
rect 12355 273330 12635 273340
rect 12355 273060 12360 273330
rect 12630 273060 12635 273330
rect 12355 273050 12635 273060
rect 12830 273320 12870 273570
rect 13120 273320 13160 273570
rect 12830 273250 12840 273320
rect 12910 273250 13080 273320
rect 13150 273250 13160 273320
rect 6871 272850 10370 272878
rect 12830 273010 13160 273250
rect 12830 272940 12840 273010
rect 12910 272940 13080 273010
rect 13150 272940 13160 273010
rect 12830 272690 13160 272940
rect 12830 272620 12840 272690
rect 12910 272620 13080 272690
rect 13150 272620 13160 272690
rect 6871 272422 10370 272450
rect 6871 269078 6891 272422
rect 6955 269078 10370 272422
rect 12830 272380 13160 272620
rect 12830 272310 12840 272380
rect 12910 272310 13080 272380
rect 13150 272310 13160 272380
rect 12355 272280 12635 272290
rect 12355 272010 12360 272280
rect 12630 272010 12635 272280
rect 12355 272000 12635 272010
rect 12830 272060 13160 272310
rect 12830 271990 12840 272060
rect 12910 271990 13080 272060
rect 13150 271990 13160 272060
rect 12830 271740 12870 271990
rect 13120 271740 13160 271990
rect 12830 271670 12840 271740
rect 12910 271670 13080 271740
rect 13150 271670 13160 271740
rect 12830 271430 13160 271670
rect 12830 271360 12840 271430
rect 12910 271360 13080 271430
rect 13150 271360 13160 271430
rect 12830 271110 13160 271360
rect 12830 271040 12840 271110
rect 12910 271040 13080 271110
rect 13150 271040 13160 271110
rect 12830 270790 13160 271040
rect 12830 270720 12840 270790
rect 12910 270720 13080 270790
rect 13150 270720 13160 270790
rect 12830 270480 13160 270720
rect 12830 270410 12840 270480
rect 12910 270410 13080 270480
rect 13150 270410 13160 270480
rect 12830 270160 13160 270410
rect 12830 270090 12840 270160
rect 12910 270090 13080 270160
rect 13150 270090 13160 270160
rect 12830 269850 12860 270090
rect 13110 269850 13160 270090
rect 12830 269780 12840 269850
rect 12910 269780 13080 269840
rect 13150 269780 13160 269850
rect 12830 269530 13160 269780
rect 12830 269460 12840 269530
rect 12910 269460 13080 269530
rect 13150 269460 13160 269530
rect 13440 275700 13770 275850
rect 13440 275630 13450 275700
rect 13520 275630 13690 275700
rect 13760 275630 13770 275700
rect 13440 275380 13770 275630
rect 14020 275700 14160 276320
rect 14020 275630 14060 275700
rect 14130 275630 14160 275700
rect 14020 275600 14160 275630
rect 13440 275310 13450 275380
rect 13520 275310 13690 275380
rect 13760 275310 13770 275380
rect 13440 275060 13770 275310
rect 13440 274990 13450 275060
rect 13520 274990 13690 275060
rect 13760 274990 13770 275060
rect 13440 274750 13770 274990
rect 13440 274680 13450 274750
rect 13520 274680 13690 274750
rect 13760 274680 13770 274750
rect 13440 274430 13770 274680
rect 13440 274360 13450 274430
rect 13520 274360 13690 274430
rect 13760 274360 13770 274430
rect 13440 274110 13770 274360
rect 15140 274720 15440 274760
rect 15140 274640 15160 274720
rect 15240 274640 15340 274720
rect 15420 274640 15440 274720
rect 15140 274350 15440 274640
rect 13440 274040 13450 274110
rect 13520 274040 13690 274110
rect 13760 274040 13770 274110
rect 13440 273800 13770 274040
rect 13440 273730 13450 273800
rect 13520 273730 13690 273800
rect 13760 273730 13770 273800
rect 13440 273480 13770 273730
rect 13440 273410 13450 273480
rect 13520 273410 13690 273480
rect 13760 273410 13770 273480
rect 13440 273170 13770 273410
rect 14500 274190 14800 274350
rect 14500 274120 14510 274190
rect 14580 274130 14720 274190
rect 14790 274120 14800 274190
rect 14500 273880 14520 274120
rect 14780 273880 14800 274120
rect 14500 273810 14510 273880
rect 14580 273810 14720 273870
rect 14790 273810 14800 273880
rect 14500 273560 14800 273810
rect 14500 273490 14510 273560
rect 14580 273490 14720 273560
rect 14790 273490 14800 273560
rect 13440 273100 13450 273170
rect 13520 273100 13690 273170
rect 13760 273100 13770 273170
rect 13440 272850 13770 273100
rect 13995 273330 14275 273340
rect 13995 273060 14000 273330
rect 14270 273060 14275 273330
rect 13995 273050 14275 273060
rect 14500 273250 14800 273490
rect 14500 273180 14510 273250
rect 14580 273180 14720 273250
rect 14790 273180 14800 273250
rect 13440 272780 13450 272850
rect 13520 272780 13690 272850
rect 13760 272780 13770 272850
rect 13440 272530 13770 272780
rect 13440 272460 13450 272530
rect 13520 272460 13690 272530
rect 13760 272460 13770 272530
rect 13440 272220 13770 272460
rect 14500 272930 14800 273180
rect 14500 272860 14510 272930
rect 14580 272870 14720 272930
rect 14790 272860 14800 272930
rect 14500 272610 14520 272860
rect 14780 272610 14800 272860
rect 14500 272540 14510 272610
rect 14580 272540 14720 272610
rect 14790 272540 14800 272610
rect 14500 272300 14800 272540
rect 13440 272150 13450 272220
rect 13520 272150 13690 272220
rect 13760 272150 13770 272220
rect 13440 271900 13770 272150
rect 13995 272280 14275 272290
rect 13995 272010 14000 272280
rect 14270 272010 14275 272280
rect 13995 272000 14275 272010
rect 14500 272230 14510 272300
rect 14580 272230 14720 272300
rect 14790 272230 14800 272300
rect 13440 271830 13450 271900
rect 13520 271830 13690 271900
rect 13760 271830 13770 271900
rect 13440 271580 13770 271830
rect 13440 271510 13450 271580
rect 13520 271510 13690 271580
rect 13760 271510 13770 271580
rect 13440 271270 13770 271510
rect 13440 271200 13450 271270
rect 13520 271200 13690 271270
rect 13760 271200 13770 271270
rect 13440 270950 13770 271200
rect 14500 271980 14800 272230
rect 14500 271910 14510 271980
rect 14580 271910 14720 271980
rect 14790 271910 14800 271980
rect 14500 271660 14800 271910
rect 14500 271590 14510 271660
rect 14580 271600 14720 271660
rect 14790 271590 14800 271660
rect 14500 271350 14520 271590
rect 14780 271350 14800 271590
rect 14500 271280 14510 271350
rect 14580 271280 14720 271340
rect 14790 271280 14800 271350
rect 14500 271030 14800 271280
rect 14500 270960 14510 271030
rect 14580 270960 14720 271030
rect 14790 270960 14800 271030
rect 15140 274280 15150 274350
rect 15220 274280 15360 274350
rect 15430 274280 15440 274350
rect 15960 274320 16440 286000
rect 17600 275300 18600 296400
rect 17600 275200 17700 275300
rect 17800 275200 18000 275300
rect 18200 275200 18400 275300
rect 18500 275200 18600 275300
rect 17600 275100 18600 275200
rect 19000 293800 265000 299000
rect 266000 342560 281300 342700
rect 266000 342500 281040 342560
rect 281100 342500 281140 342560
rect 281200 342500 281300 342560
rect 266000 342460 281300 342500
rect 266000 342400 281040 342460
rect 281100 342400 281140 342460
rect 281200 342400 281300 342460
rect 266000 342300 281300 342400
rect 294700 342420 317000 342500
rect 294700 342360 294760 342420
rect 294820 342360 294860 342420
rect 294920 342360 317000 342420
rect 294700 342320 317000 342360
rect 19000 275000 19600 293800
rect 25680 289800 26140 290200
rect 25680 289600 25800 289800
rect 26000 289600 26140 289800
rect 25680 289400 26140 289600
rect 25680 289200 25800 289400
rect 26000 289200 26140 289400
rect 25680 289000 26140 289200
rect 25680 288800 25800 289000
rect 26000 288800 26140 289000
rect 25680 288600 26140 288800
rect 25680 288400 25800 288600
rect 26000 288400 26140 288600
rect 25680 288200 26140 288400
rect 25680 288000 25800 288200
rect 26000 288000 26140 288200
rect 25680 287800 26140 288000
rect 25680 287600 25800 287800
rect 26000 287600 26140 287800
rect 25680 287400 26140 287600
rect 25680 287200 25800 287400
rect 26000 287200 26140 287400
rect 25680 287000 26140 287200
rect 25680 286800 25800 287000
rect 26000 286800 26140 287000
rect 25680 286600 26140 286800
rect 25680 286400 25800 286600
rect 26000 286400 26140 286600
rect 25680 286200 26140 286400
rect 25680 286000 25800 286200
rect 26000 286000 26140 286200
rect 17600 274740 19600 275000
rect 17600 274620 17630 274740
rect 17750 274620 17850 274740
rect 17970 274620 19600 274740
rect 17600 274600 19600 274620
rect 20600 275700 21000 275800
rect 20600 275630 20670 275700
rect 20740 275630 20830 275700
rect 20900 275630 21000 275700
rect 16685 274350 16765 274360
rect 16895 274350 16975 274360
rect 15140 274040 15440 274280
rect 15140 273970 15150 274040
rect 15220 273970 15360 274040
rect 15430 273970 15440 274040
rect 15140 273720 15440 273970
rect 15140 273650 15150 273720
rect 15220 273650 15360 273720
rect 15430 273650 15440 273720
rect 15140 273400 15440 273650
rect 16050 274190 16350 274320
rect 16050 274120 16060 274190
rect 16130 274130 16270 274190
rect 16340 274120 16350 274190
rect 16050 273880 16070 274120
rect 16330 273880 16350 274120
rect 16050 273810 16060 273880
rect 16130 273810 16270 273870
rect 16340 273810 16350 273880
rect 16050 273560 16350 273810
rect 15140 273330 15150 273400
rect 15220 273330 15360 273400
rect 15430 273330 15440 273400
rect 15140 273090 15440 273330
rect 15605 273540 15875 273550
rect 15605 273280 15610 273540
rect 15870 273280 15875 273540
rect 15605 273270 15875 273280
rect 16050 273490 16060 273560
rect 16130 273490 16270 273560
rect 16340 273490 16350 273560
rect 15140 273020 15150 273090
rect 15220 273020 15360 273090
rect 15430 273020 15440 273090
rect 15140 272770 15440 273020
rect 15140 272700 15150 272770
rect 15220 272700 15360 272770
rect 15430 272700 15440 272770
rect 15140 272460 15440 272700
rect 15140 272390 15150 272460
rect 15220 272390 15360 272460
rect 15430 272390 15440 272460
rect 15140 272140 15440 272390
rect 15140 272070 15150 272140
rect 15220 272070 15360 272140
rect 15430 272070 15440 272140
rect 15140 271820 15440 272070
rect 16050 273240 16350 273490
rect 16050 273170 16060 273240
rect 16130 273170 16270 273240
rect 16340 273170 16350 273240
rect 16050 272930 16350 273170
rect 16050 272860 16060 272930
rect 16130 272870 16270 272930
rect 16340 272860 16350 272930
rect 16050 272610 16070 272860
rect 16330 272610 16350 272860
rect 16050 272540 16060 272610
rect 16130 272540 16270 272610
rect 16340 272540 16350 272610
rect 16050 272300 16350 272540
rect 16050 272230 16060 272300
rect 16130 272230 16270 272300
rect 16340 272230 16350 272300
rect 15140 271750 15150 271820
rect 15220 271750 15360 271820
rect 15430 271750 15440 271820
rect 15605 272040 15875 272050
rect 15605 271780 15610 272040
rect 15870 271780 15875 272040
rect 15605 271770 15875 271780
rect 16050 271980 16350 272230
rect 16050 271910 16060 271980
rect 16130 271910 16270 271980
rect 16340 271910 16350 271980
rect 15140 271510 15440 271750
rect 15140 271440 15150 271510
rect 15220 271440 15360 271510
rect 15430 271440 15440 271510
rect 15140 271190 15440 271440
rect 15140 271120 15150 271190
rect 15220 271120 15360 271190
rect 15430 271120 15440 271190
rect 14505 270950 14585 270960
rect 14715 270950 14795 270960
rect 13440 270880 13450 270950
rect 13520 270880 13690 270950
rect 13760 270880 13770 270950
rect 13440 270640 13770 270880
rect 13440 270570 13450 270640
rect 13520 270570 13690 270640
rect 13760 270570 13770 270640
rect 13440 270320 13770 270570
rect 15140 270660 15440 271120
rect 16050 271660 16350 271910
rect 16050 271590 16060 271660
rect 16130 271600 16270 271660
rect 16340 271590 16350 271660
rect 16050 271350 16070 271590
rect 16330 271350 16350 271590
rect 16050 271280 16060 271350
rect 16130 271280 16270 271340
rect 16340 271280 16350 271350
rect 16050 271030 16350 271280
rect 16050 270960 16060 271030
rect 16130 270960 16270 271030
rect 16340 270960 16350 271030
rect 16680 274280 16690 274350
rect 16760 274280 16900 274350
rect 16970 274280 16980 274350
rect 16680 274030 16980 274280
rect 16680 273960 16690 274030
rect 16760 273960 16900 274030
rect 16970 273960 16980 274030
rect 16680 273720 16980 273960
rect 16680 273650 16690 273720
rect 16760 273650 16900 273720
rect 16970 273650 16980 273720
rect 16680 273400 16980 273650
rect 16680 273330 16690 273400
rect 16760 273330 16900 273400
rect 16970 273330 16980 273400
rect 16680 273090 16980 273330
rect 16680 273020 16690 273090
rect 16760 273020 16900 273090
rect 16970 273020 16980 273090
rect 16680 272770 16980 273020
rect 16680 272700 16690 272770
rect 16760 272700 16900 272770
rect 16970 272700 16980 272770
rect 16680 272450 16980 272700
rect 16680 272380 16690 272450
rect 16760 272380 16900 272450
rect 16970 272380 16980 272450
rect 16680 272140 16980 272380
rect 16680 272070 16690 272140
rect 16760 272070 16900 272140
rect 16970 272070 16980 272140
rect 16680 271820 16980 272070
rect 16680 271750 16690 271820
rect 16760 271750 16900 271820
rect 16970 271750 16980 271820
rect 16680 271510 16980 271750
rect 16680 271440 16690 271510
rect 16760 271440 16900 271510
rect 16970 271440 16980 271510
rect 16680 271190 16980 271440
rect 16680 271120 16690 271190
rect 16760 271120 16900 271190
rect 16970 271120 16980 271190
rect 16680 270960 16980 271120
rect 17610 273080 17990 274600
rect 17610 273010 17620 273080
rect 17690 273010 17910 273080
rect 17980 273010 17990 273080
rect 17610 272760 17990 273010
rect 17610 272690 17620 272760
rect 17690 272690 17910 272760
rect 17980 272690 17990 272760
rect 17610 272450 17990 272690
rect 17610 272380 17620 272450
rect 17690 272380 17910 272450
rect 17980 272380 17990 272450
rect 17610 272130 17990 272380
rect 17610 272060 17620 272130
rect 17690 272060 17910 272130
rect 17980 272060 17990 272130
rect 16055 270950 16135 270960
rect 16265 270950 16345 270960
rect 15140 270580 15160 270660
rect 15240 270580 15340 270660
rect 15420 270580 15440 270660
rect 15140 270540 15440 270580
rect 17610 270680 17990 272060
rect 18170 274500 18550 274520
rect 18170 274380 18190 274500
rect 18310 274380 18410 274500
rect 18530 274380 18550 274500
rect 18170 273240 18550 274380
rect 18170 273170 18180 273240
rect 18250 273170 18470 273240
rect 18540 273170 18550 273240
rect 18170 272920 18550 273170
rect 18170 272850 18180 272920
rect 18250 272850 18470 272920
rect 18540 272850 18550 272920
rect 18170 272600 18550 272850
rect 19130 274500 19510 274520
rect 19130 274380 19150 274500
rect 19270 274380 19370 274500
rect 19490 274380 19510 274500
rect 19130 273080 19510 274380
rect 20600 274240 21000 275630
rect 24860 275020 24980 275040
rect 24860 274940 24880 275020
rect 24960 274940 24980 275020
rect 24860 274880 24980 274940
rect 24860 274800 24880 274880
rect 24960 274800 24980 274880
rect 24860 274740 24980 274800
rect 24860 274660 24880 274740
rect 24960 274660 24980 274740
rect 22175 274490 22255 274500
rect 22355 274490 22435 274500
rect 22170 274420 22180 274490
rect 22250 274420 22360 274490
rect 22430 274420 22440 274490
rect 20600 274170 20660 274240
rect 20730 274170 20840 274240
rect 20910 274170 21000 274240
rect 19130 273010 19140 273080
rect 19210 273010 19430 273080
rect 19500 273010 19510 273080
rect 18170 272530 18180 272600
rect 18250 272530 18470 272600
rect 18540 272530 18550 272600
rect 18170 272290 18550 272530
rect 18705 272780 18975 272790
rect 18705 272520 18710 272780
rect 18970 272520 18975 272780
rect 18705 272510 18975 272520
rect 19130 272760 19510 273010
rect 19130 272690 19140 272760
rect 19210 272690 19430 272760
rect 19500 272690 19510 272760
rect 18170 272220 18180 272290
rect 18250 272220 18470 272290
rect 18540 272220 18550 272290
rect 18170 270920 18550 272220
rect 18170 270800 18190 270920
rect 18310 270800 18410 270920
rect 18530 270800 18550 270920
rect 18170 270780 18550 270800
rect 19130 272450 19510 272690
rect 19130 272380 19140 272450
rect 19210 272380 19430 272450
rect 19500 272380 19510 272450
rect 19130 272130 19510 272380
rect 19130 272060 19140 272130
rect 19210 272060 19430 272130
rect 19500 272060 19510 272130
rect 19130 270920 19510 272060
rect 19690 274030 20070 274060
rect 19690 273960 19720 274030
rect 19790 273960 19970 274030
rect 20040 273960 20070 274030
rect 19690 273240 20070 273960
rect 19690 273170 19700 273240
rect 19770 273170 19990 273240
rect 20060 273170 20070 273240
rect 19690 272920 20070 273170
rect 19690 272850 19700 272920
rect 19770 272850 19990 272920
rect 20060 272850 20070 272920
rect 19690 272600 20070 272850
rect 20600 273720 21000 274170
rect 20600 273650 20660 273720
rect 20730 273650 20840 273720
rect 20910 273650 21000 273720
rect 20600 273200 21000 273650
rect 20600 273130 20660 273200
rect 20730 273130 20840 273200
rect 20910 273130 21000 273200
rect 19690 272530 19700 272600
rect 19770 272530 19990 272600
rect 20060 272530 20070 272600
rect 19690 272290 20070 272530
rect 20225 272780 20495 272790
rect 20225 272520 20230 272780
rect 20490 272520 20495 272780
rect 20225 272510 20495 272520
rect 20600 272690 21000 273130
rect 20600 272620 20660 272690
rect 20730 272620 20840 272690
rect 20910 272620 21000 272690
rect 19690 272220 19700 272290
rect 19770 272220 19990 272290
rect 20060 272220 20070 272290
rect 19690 271510 20070 272220
rect 19690 271440 19720 271510
rect 19790 271440 19970 271510
rect 20040 271440 20070 271510
rect 19690 271410 20070 271440
rect 20600 272170 21000 272620
rect 20600 272100 20660 272170
rect 20730 272100 20840 272170
rect 20910 272100 21000 272170
rect 20600 271660 21000 272100
rect 20600 271590 20660 271660
rect 20730 271590 20840 271660
rect 20910 271590 21000 271660
rect 19130 270800 19150 270920
rect 19270 270800 19370 270920
rect 19490 270800 19510 270920
rect 19130 270780 19510 270800
rect 20600 271140 21000 271590
rect 20600 271070 20660 271140
rect 20730 271070 20840 271140
rect 20910 271070 21000 271140
rect 21320 273980 21590 274240
rect 21320 273910 21330 273980
rect 21400 273910 21510 273980
rect 21580 273910 21590 273980
rect 21320 273810 21590 273910
rect 21320 273560 21330 273810
rect 21580 273560 21590 273810
rect 21320 273460 21590 273560
rect 21320 273390 21330 273460
rect 21400 273390 21510 273460
rect 21580 273390 21590 273460
rect 21320 272950 21590 273390
rect 21320 272880 21330 272950
rect 21400 272880 21510 272950
rect 21580 272880 21590 272950
rect 21320 272430 21590 272880
rect 22170 273980 22440 274420
rect 22170 273910 22180 273980
rect 22250 273910 22360 273980
rect 22430 273910 22440 273980
rect 22170 273460 22440 273910
rect 22170 273390 22180 273460
rect 22250 273390 22360 273460
rect 22430 273390 22440 273460
rect 22170 272940 22440 273390
rect 22170 272870 22180 272940
rect 22250 272870 22360 272940
rect 22430 272870 22440 272940
rect 21745 272780 22005 272790
rect 21745 272530 21750 272780
rect 22000 272530 22005 272780
rect 21745 272520 22005 272530
rect 21320 272360 21330 272430
rect 21400 272360 21510 272430
rect 21580 272360 21590 272430
rect 21320 271910 21590 272360
rect 21320 271840 21330 271910
rect 21400 271840 21510 271910
rect 21580 271840 21590 271910
rect 21320 271750 21590 271840
rect 21320 271500 21330 271750
rect 21580 271500 21590 271750
rect 21320 271400 21590 271500
rect 21320 271330 21330 271400
rect 21400 271330 21510 271400
rect 21580 271330 21590 271400
rect 21320 271070 21590 271330
rect 22170 272430 22440 272870
rect 22170 272360 22180 272430
rect 22250 272360 22360 272430
rect 22430 272360 22440 272430
rect 22170 271910 22440 272360
rect 22170 271840 22180 271910
rect 22250 271840 22360 271910
rect 22430 271840 22440 271910
rect 22170 271400 22440 271840
rect 22170 271330 22180 271400
rect 22250 271330 22360 271400
rect 22430 271330 22440 271400
rect 17610 270560 17630 270680
rect 17750 270560 17850 270680
rect 17970 270560 17990 270680
rect 17610 270540 17990 270560
rect 13440 270250 13450 270320
rect 13520 270250 13690 270320
rect 13760 270250 13770 270320
rect 13440 270000 13770 270250
rect 13440 269930 13450 270000
rect 13520 269930 13690 270000
rect 13760 269930 13770 270000
rect 13440 269690 13770 269930
rect 19200 270100 20000 270200
rect 19200 270000 19300 270100
rect 19400 270000 19500 270100
rect 19700 270000 19800 270100
rect 19900 270000 20000 270100
rect 13440 269620 13450 269690
rect 13520 269620 13690 269690
rect 13760 269620 13770 269690
rect 13440 269460 13770 269620
rect 14020 269690 14160 269720
rect 14020 269620 14060 269690
rect 14130 269620 14160 269690
rect 12835 269450 12915 269460
rect 13075 269450 13155 269460
rect 6871 269050 10370 269078
rect 14020 268990 14160 269620
rect 14020 268900 14040 268990
rect 14140 268900 14160 268990
rect 14020 268800 14160 268900
rect 14020 268710 14040 268800
rect 14140 268710 14160 268800
rect 14020 268690 14160 268710
rect 6871 268622 10370 268650
rect 6871 265278 6891 268622
rect 6955 265278 10370 268622
rect 14535 267300 14645 267310
rect 14535 267120 14540 267300
rect 14640 267120 14645 267300
rect 14535 267110 14645 267120
rect 14940 267280 15860 267320
rect 14940 267120 15000 267280
rect 15160 267120 15220 267280
rect 15380 267120 15440 267280
rect 15600 267120 15660 267280
rect 15820 267120 15860 267280
rect 14535 266880 14645 266890
rect 14535 266700 14540 266880
rect 14640 266700 14645 266880
rect 14535 266690 14645 266700
rect 14940 266860 15860 267120
rect 14940 266700 15000 266860
rect 15160 266700 15220 266860
rect 15380 266700 15440 266860
rect 15600 266700 15660 266860
rect 15820 266700 15860 266860
rect 6871 265250 10370 265278
rect 13060 265000 13280 265020
rect 13060 264930 13080 265000
rect 13150 264930 13280 265000
rect 13060 264890 13280 264930
rect 13060 264820 13190 264890
rect 13260 264820 13280 264890
rect 13060 264800 13280 264820
rect 0 252510 5050 253200
rect -800 252398 5050 252510
rect 14940 252580 15860 266700
rect 14940 252460 14980 252580
rect 15100 252460 15160 252580
rect 15280 252460 15340 252580
rect 15460 252460 15520 252580
rect 15640 252460 15700 252580
rect 15820 252460 15860 252580
rect 14940 252440 15860 252460
rect 0 252100 5050 252398
rect 9650 252400 11600 252410
rect 9650 252380 9800 252400
rect 10000 252380 10200 252400
rect 10400 252380 10600 252400
rect 10800 252380 11000 252400
rect 11200 252380 11400 252400
rect 5815 252320 5945 252330
rect 5815 252200 5820 252320
rect 5940 252200 5945 252320
rect 5815 252190 5945 252200
rect 9650 252320 9680 252380
rect 9740 252320 9800 252380
rect 10000 252320 10045 252380
rect 10105 252320 10200 252380
rect 10400 252320 10415 252380
rect 10475 252320 10600 252380
rect 10800 252320 10805 252380
rect 10865 252320 10965 252380
rect 11215 252320 11330 252380
rect 11390 252320 11400 252380
rect 9650 252200 9800 252320
rect 10000 252200 10200 252320
rect 10400 252200 10600 252320
rect 10800 252200 11000 252320
rect 11200 252200 11400 252320
rect 9650 252180 11600 252200
rect -800 251216 480 251328
rect -800 250034 480 250146
rect 3950 249194 5050 252100
rect 5815 252120 5945 252130
rect 5815 252000 5820 252120
rect 5940 252000 5945 252120
rect 5815 251990 5945 252000
rect 9650 252120 9680 252180
rect 9740 252120 9845 252180
rect 9905 252120 10045 252180
rect 10105 252120 10235 252180
rect 10295 252120 10415 252180
rect 10475 252120 10615 252180
rect 10675 252120 10805 252180
rect 10865 252120 10965 252180
rect 11025 252120 11155 252180
rect 11215 252120 11330 252180
rect 11390 252120 11470 252180
rect 11530 252120 11600 252180
rect 9650 252000 11600 252120
rect 9650 251980 9800 252000
rect 10000 251980 10200 252000
rect 10400 251980 10600 252000
rect 10800 251980 11000 252000
rect 11200 251980 11400 252000
rect 5815 251920 5945 251930
rect 5815 251800 5820 251920
rect 5940 251800 5945 251920
rect 5815 251790 5945 251800
rect 9650 251920 9680 251980
rect 9740 251920 9800 251980
rect 10000 251920 10045 251980
rect 10105 251920 10200 251980
rect 10400 251920 10415 251980
rect 10475 251920 10600 251980
rect 10800 251920 10805 251980
rect 10865 251920 10965 251980
rect 11215 251920 11330 251980
rect 11390 251920 11400 251980
rect 9650 251800 9800 251920
rect 10000 251800 10200 251920
rect 10400 251800 10600 251920
rect 10800 251800 11000 251920
rect 11200 251800 11400 251920
rect 9650 251790 11600 251800
rect 9650 251730 9680 251790
rect 9740 251730 9845 251790
rect 9905 251730 10045 251790
rect 10105 251730 10235 251790
rect 10295 251730 10415 251790
rect 10475 251730 10615 251790
rect 10675 251730 10805 251790
rect 10865 251730 10965 251790
rect 11025 251730 11155 251790
rect 11215 251730 11330 251790
rect 11390 251730 11470 251790
rect 11530 251730 11600 251790
rect 5815 251720 5945 251730
rect 5815 251600 5820 251720
rect 5940 251600 5945 251720
rect 5815 251590 5945 251600
rect 9650 251600 11600 251730
rect 9650 251590 9800 251600
rect 10000 251590 10200 251600
rect 10400 251590 10600 251600
rect 10800 251590 11000 251600
rect 11200 251590 11400 251600
rect 9650 251530 9680 251590
rect 9740 251530 9800 251590
rect 10000 251530 10045 251590
rect 10105 251530 10200 251590
rect 10400 251530 10415 251590
rect 10475 251530 10600 251590
rect 10800 251530 10805 251590
rect 10865 251530 10965 251590
rect 11215 251530 11330 251590
rect 11390 251530 11400 251590
rect 5815 251520 5945 251530
rect 5815 251400 5820 251520
rect 5940 251400 5945 251520
rect 5815 251390 5945 251400
rect 9650 251400 9800 251530
rect 10000 251400 10200 251530
rect 10400 251400 10600 251530
rect 10800 251400 11000 251530
rect 11200 251400 11400 251530
rect 9650 251340 9680 251400
rect 9740 251390 11600 251400
rect 9740 251340 9845 251390
rect 9650 251330 9845 251340
rect 9905 251330 10045 251390
rect 10105 251330 10235 251390
rect 10295 251330 10415 251390
rect 10475 251330 10615 251390
rect 10675 251330 10805 251390
rect 10865 251330 10965 251390
rect 11025 251330 11155 251390
rect 11215 251330 11330 251390
rect 11390 251330 11470 251390
rect 11530 251330 11600 251390
rect 9650 251300 11600 251330
rect 5700 249194 8200 249200
rect 3950 249000 8200 249194
rect -800 248852 480 248964
rect 3950 248800 5800 249000
rect 6000 248800 6200 249000
rect 6400 248800 6600 249000
rect 6800 248800 7000 249000
rect 7200 248800 7400 249000
rect 7600 248800 7800 249000
rect 8000 248800 8200 249000
rect 3950 248600 8200 248800
rect 3950 248400 5800 248600
rect 6000 248400 6200 248600
rect 6400 248400 6600 248600
rect 6800 248400 7000 248600
rect 7200 248400 7400 248600
rect 7600 248400 7800 248600
rect 8000 248400 8200 248600
rect 3950 248200 8200 248400
rect 3950 248000 5800 248200
rect 6000 248000 6200 248200
rect 6400 248000 6600 248200
rect 6800 248000 7000 248200
rect 7200 248000 7400 248200
rect 7600 248000 7800 248200
rect 8000 248000 8200 248200
rect 3950 247800 8200 248000
rect -800 247670 480 247782
rect 3950 247600 5800 247800
rect 6000 247600 6200 247800
rect 6400 247600 6600 247800
rect 6800 247600 7000 247800
rect 7200 247600 7400 247800
rect 7600 247600 7800 247800
rect 8000 247600 8200 247800
rect 3950 247400 8200 247600
rect 3950 247200 5800 247400
rect 6000 247200 6200 247400
rect 6400 247200 6600 247400
rect 6800 247200 7000 247400
rect 7200 247200 7400 247400
rect 7600 247200 7800 247400
rect 8000 247200 8200 247400
rect 3950 247000 8200 247200
rect 3950 246800 5800 247000
rect 6000 246800 6200 247000
rect 6400 246800 6600 247000
rect 6800 246800 7000 247000
rect 7200 246800 7400 247000
rect 7600 246800 7800 247000
rect 8000 246800 8200 247000
rect 3950 246600 8200 246800
rect -800 246488 480 246600
rect 3950 246400 5800 246600
rect 6000 246400 6200 246600
rect 6400 246400 6600 246600
rect 6800 246400 7000 246600
rect 7200 246400 7400 246600
rect 7600 246400 7800 246600
rect 8000 246400 8200 246600
rect 3950 246200 8200 246400
rect 3950 246025 5800 246200
rect 6000 246000 6200 246200
rect 6400 246000 6600 246200
rect 6800 246000 7000 246200
rect 7200 246000 7400 246200
rect 7600 246000 7800 246200
rect 8000 246000 8200 246200
rect 5800 245800 8200 246000
rect 6000 245600 6200 245800
rect 6400 245600 6600 245800
rect 6800 245600 7000 245800
rect 7200 245600 7400 245800
rect 7600 245600 7800 245800
rect 8000 245600 8200 245800
rect 5800 245400 8200 245600
rect 6000 245200 6200 245400
rect 6400 245200 6600 245400
rect 6800 245200 7000 245400
rect 7200 245200 7400 245400
rect 7600 245200 7800 245400
rect 8000 245200 8200 245400
rect 5800 245000 8200 245200
rect 6000 244800 6200 245000
rect 6400 244800 6600 245000
rect 6800 244800 7000 245000
rect 7200 244800 7400 245000
rect 7600 244800 7800 245000
rect 8000 244800 8200 245000
rect 5800 244600 8200 244800
rect 6000 244400 6200 244600
rect 6400 244400 6600 244600
rect 6800 244400 7000 244600
rect 7200 244400 7400 244600
rect 7600 244400 7800 244600
rect 8000 244400 8200 244600
rect 5800 244200 8200 244400
rect 19200 249000 20000 270000
rect 20600 269690 21000 271070
rect 22170 270880 22440 271330
rect 22170 270810 22180 270880
rect 22250 270810 22360 270880
rect 22430 270810 22440 270880
rect 22840 274230 23110 274490
rect 22840 274160 22850 274230
rect 22920 274160 23030 274230
rect 23100 274160 23110 274230
rect 22840 274070 23110 274160
rect 22840 273820 22850 274070
rect 23100 273820 23110 274070
rect 22840 273720 23110 273820
rect 22840 273650 22850 273720
rect 22920 273650 23030 273720
rect 23100 273650 23110 273720
rect 22840 273200 23110 273650
rect 22840 273130 22850 273200
rect 22920 273130 23030 273200
rect 23100 273130 23110 273200
rect 22840 272690 23110 273130
rect 24380 273470 24500 273480
rect 24380 273390 24400 273470
rect 24480 273390 24500 273470
rect 24380 272950 24500 273390
rect 24380 272870 24400 272950
rect 24480 272870 24500 272950
rect 22840 272620 22850 272690
rect 22920 272620 23030 272690
rect 23100 272620 23110 272690
rect 22840 272170 23110 272620
rect 23275 272780 23535 272790
rect 23275 272530 23280 272780
rect 23530 272530 23535 272780
rect 23275 272520 23535 272530
rect 22840 272100 22850 272170
rect 22920 272100 23030 272170
rect 23100 272100 23110 272170
rect 22840 271650 23110 272100
rect 24380 272430 24500 272870
rect 24380 272350 24400 272430
rect 24480 272350 24500 272430
rect 24380 271930 24500 272350
rect 24380 271800 24500 271810
rect 24860 273210 24980 274660
rect 25680 273690 26140 286000
rect 266000 277654 271200 342300
rect 294700 342260 294760 342320
rect 294820 342260 294860 342320
rect 294920 342260 317000 342320
rect 294700 342100 317000 342260
rect 288290 340800 288610 340805
rect 31015 276140 31265 276150
rect 31015 275900 31020 276140
rect 31260 275900 31265 276140
rect 31015 275890 31265 275900
rect 32735 276140 32985 276150
rect 32735 275900 32740 276140
rect 32980 275900 32985 276140
rect 32735 275890 32985 275900
rect 34455 276140 34705 276150
rect 34455 275900 34460 276140
rect 34700 275900 34705 276140
rect 34455 275890 34705 275900
rect 35935 276140 36185 276150
rect 35935 275900 35940 276140
rect 36180 275900 36185 276140
rect 35935 275890 36185 275900
rect 37655 276140 37905 276150
rect 37655 275900 37660 276140
rect 37900 275900 37905 276140
rect 37655 275890 37905 275900
rect 39255 276140 39505 276150
rect 39255 275900 39260 276140
rect 39500 275900 39505 276140
rect 39255 275890 39505 275900
rect 40975 276140 41225 276150
rect 40975 275900 40980 276140
rect 41220 275900 41225 276140
rect 40975 275890 41225 275900
rect 42575 276140 42825 276150
rect 42575 275900 42580 276140
rect 42820 275900 42825 276140
rect 42575 275890 42825 275900
rect 44295 276140 44545 276150
rect 44295 275900 44300 276140
rect 44540 275900 44545 276140
rect 44295 275890 44545 275900
rect 46010 275040 271200 277654
rect 26900 274980 271200 275040
rect 26900 274900 26960 274980
rect 27040 274900 271200 274980
rect 26900 274860 271200 274900
rect 26900 274780 26960 274860
rect 27040 274780 271200 274860
rect 26900 274740 271200 274780
rect 26900 274660 26960 274740
rect 27040 274660 271200 274740
rect 26900 274640 271200 274660
rect 25680 273670 26320 273690
rect 25680 273590 25860 273670
rect 25940 273590 26080 273670
rect 26160 273590 26220 273670
rect 26300 273590 26320 273670
rect 25680 273570 26320 273590
rect 25680 273470 26140 273570
rect 25680 273440 25860 273470
rect 24860 273130 24880 273210
rect 24960 273130 24980 273210
rect 24860 272690 24980 273130
rect 24860 272610 24880 272690
rect 24960 272610 24980 272690
rect 24860 272170 24980 272610
rect 24860 272090 24880 272170
rect 24960 272090 24980 272170
rect 22840 271580 22850 271650
rect 22920 271580 23030 271650
rect 23100 271580 23110 271650
rect 22840 271490 23110 271580
rect 22840 271240 22850 271490
rect 23100 271240 23110 271490
rect 22840 271140 23110 271240
rect 22840 271070 22850 271140
rect 22920 271070 23030 271140
rect 23100 271070 23110 271140
rect 22840 270810 23110 271070
rect 22175 270800 22255 270810
rect 22355 270800 22435 270810
rect 24860 270620 24980 272090
rect 25840 273390 25860 273440
rect 25940 273440 26140 273470
rect 29300 273440 29380 273450
rect 25940 273390 25960 273440
rect 25840 272950 25960 273390
rect 29300 273380 29310 273440
rect 29370 273380 29380 273440
rect 28350 273190 28480 273210
rect 28350 273100 28370 273190
rect 28460 273100 28480 273190
rect 25840 272870 25860 272950
rect 25940 272870 25960 272950
rect 27465 273010 27595 273020
rect 27465 272890 27470 273010
rect 27590 272890 27595 273010
rect 27465 272880 27595 272890
rect 25840 272430 25960 272870
rect 25840 272350 25860 272430
rect 25940 272350 25960 272430
rect 28350 272680 28480 273100
rect 29300 272920 29380 273380
rect 29300 272860 29310 272920
rect 29370 272860 29380 272920
rect 28350 272590 28370 272680
rect 28460 272590 28480 272680
rect 25840 271920 25960 272350
rect 27475 272390 27605 272400
rect 27475 272270 27480 272390
rect 27600 272270 27605 272390
rect 27475 272260 27605 272270
rect 28350 272160 28480 272590
rect 28745 272670 28845 272680
rect 28745 272580 28750 272670
rect 28840 272580 28845 272670
rect 28745 272570 28845 272580
rect 28350 272070 28370 272160
rect 28460 272070 28480 272160
rect 28350 272050 28480 272070
rect 29300 272410 29380 272860
rect 29300 272350 29310 272410
rect 29370 272350 29380 272410
rect 25840 271840 25860 271920
rect 25940 271840 25960 271920
rect 25840 271710 25960 271840
rect 29300 271890 29380 272350
rect 29300 271830 29310 271890
rect 29370 271830 29380 271890
rect 29710 273180 29790 273430
rect 29710 273120 29720 273180
rect 29780 273120 29790 273180
rect 29710 272670 29790 273120
rect 29710 272610 29720 272670
rect 29780 272610 29790 272670
rect 29710 272150 29790 272610
rect 30185 272670 30285 272680
rect 30185 272580 30190 272670
rect 30280 272580 30285 272670
rect 30185 272570 30285 272580
rect 46010 272454 271200 274640
rect 272200 340720 281300 340800
rect 272200 340660 281060 340720
rect 281120 340660 281160 340720
rect 281220 340660 281300 340720
rect 272200 340620 281300 340660
rect 272200 340560 281060 340620
rect 281120 340560 281160 340620
rect 281220 340560 281300 340620
rect 272200 340400 281300 340560
rect 288290 340500 288300 340800
rect 288600 340500 288610 340800
rect 288290 340495 288610 340500
rect 29710 272090 29720 272150
rect 29780 272090 29790 272150
rect 29710 271840 29790 272090
rect 29300 271820 29380 271830
rect 25840 271630 25860 271710
rect 25940 271630 25960 271710
rect 25840 271570 25960 271630
rect 26060 271710 26320 271730
rect 26060 271630 26080 271710
rect 26160 271630 26220 271710
rect 26300 271630 26320 271710
rect 26060 271610 26320 271630
rect 24860 270540 24880 270620
rect 24960 270540 24980 270620
rect 24860 270480 24980 270540
rect 24860 270400 24880 270480
rect 24960 270400 24980 270480
rect 24860 270340 24980 270400
rect 24860 270260 24880 270340
rect 24960 270260 24980 270340
rect 24860 270240 24980 270260
rect 20600 269620 20670 269690
rect 20740 269620 20830 269690
rect 20900 269620 21000 269690
rect 20600 266200 21000 269620
rect 31015 269440 31265 269450
rect 31015 269200 31020 269440
rect 31260 269200 31265 269440
rect 31015 269190 31265 269200
rect 32735 269440 32985 269450
rect 32735 269200 32740 269440
rect 32980 269200 32985 269440
rect 32735 269190 32985 269200
rect 34455 269440 34705 269450
rect 34455 269200 34460 269440
rect 34700 269200 34705 269440
rect 34455 269190 34705 269200
rect 35935 269440 36185 269450
rect 35935 269200 35940 269440
rect 36180 269200 36185 269440
rect 35935 269190 36185 269200
rect 37655 269440 37905 269450
rect 37655 269200 37660 269440
rect 37900 269200 37905 269440
rect 37655 269190 37905 269200
rect 39255 269440 39505 269450
rect 39255 269200 39260 269440
rect 39500 269200 39505 269440
rect 39255 269190 39505 269200
rect 40975 269440 41225 269450
rect 40975 269200 40980 269440
rect 41220 269200 41225 269440
rect 40975 269190 41225 269200
rect 42575 269440 42825 269450
rect 42575 269200 42580 269440
rect 42820 269200 42825 269440
rect 42575 269190 42825 269200
rect 44295 269440 44545 269450
rect 44295 269200 44300 269440
rect 44540 269200 44545 269440
rect 44295 269190 44545 269200
rect 44695 268600 45005 268610
rect 44695 268300 44700 268600
rect 45000 268300 45005 268600
rect 44695 268290 45005 268300
rect 44695 268100 45005 268110
rect 44695 267800 44700 268100
rect 45000 267800 45005 268100
rect 44695 267790 45005 267800
rect 44695 267600 45005 267610
rect 44695 267300 44700 267600
rect 45000 267300 45005 267600
rect 44695 267290 45005 267300
rect 44695 267100 45005 267110
rect 44695 266800 44700 267100
rect 45000 266800 45005 267100
rect 44695 266790 45005 266800
rect 44695 266600 45005 266610
rect 20600 266000 20700 266200
rect 20900 266000 21000 266200
rect 20600 265800 21000 266000
rect 20600 265600 20700 265800
rect 20900 265600 21000 265800
rect 20600 265400 21000 265600
rect 20600 265200 20700 265400
rect 20900 265200 21000 265400
rect 20600 265000 21000 265200
rect 20600 264800 20700 265000
rect 20900 264800 21000 265000
rect 20600 264600 21000 264800
rect 22600 266200 27800 266400
rect 44695 266300 44700 266600
rect 45000 266300 45005 266600
rect 44695 266290 45005 266300
rect 22600 266000 22700 266200
rect 22900 266000 23100 266200
rect 23300 266000 23500 266200
rect 23700 266000 23900 266200
rect 24100 266000 24300 266200
rect 24500 266000 24700 266200
rect 24900 266000 25100 266200
rect 25300 266000 25500 266200
rect 25700 266000 25900 266200
rect 26100 266000 26300 266200
rect 26500 266000 26700 266200
rect 26900 266000 27100 266200
rect 27300 266000 27500 266200
rect 27700 266000 27800 266200
rect 22600 265800 27800 266000
rect 22600 265600 22700 265800
rect 22900 265600 23100 265800
rect 23300 265600 23500 265800
rect 23700 265600 23900 265800
rect 24100 265600 24300 265800
rect 24500 265600 24700 265800
rect 24900 265600 25100 265800
rect 25300 265600 25500 265800
rect 25700 265600 25900 265800
rect 26100 265600 26300 265800
rect 26500 265600 26700 265800
rect 26900 265600 27100 265800
rect 27300 265600 27500 265800
rect 27700 265600 27800 265800
rect 44695 266100 45005 266110
rect 44695 265800 44700 266100
rect 45000 265800 45005 266100
rect 44695 265790 45005 265800
rect 22600 265400 27800 265600
rect 22600 265200 22700 265400
rect 22900 265200 23100 265400
rect 23300 265200 23500 265400
rect 23700 265200 23900 265400
rect 24100 265200 24300 265400
rect 24500 265200 24700 265400
rect 24900 265200 25100 265400
rect 25300 265200 25500 265400
rect 25700 265200 25900 265400
rect 26100 265200 26300 265400
rect 26500 265200 26700 265400
rect 26900 265200 27100 265400
rect 27300 265200 27500 265400
rect 27700 265200 27800 265400
rect 44695 265600 45005 265610
rect 44695 265300 44700 265600
rect 45000 265300 45005 265600
rect 44695 265290 45005 265300
rect 22600 265000 27800 265200
rect 22600 264800 22700 265000
rect 22900 264800 23100 265000
rect 23300 264800 23500 265000
rect 23700 264800 23900 265000
rect 24100 264800 24300 265000
rect 24500 264800 24700 265000
rect 24900 264800 25100 265000
rect 25300 264800 25500 265000
rect 25700 264800 25900 265000
rect 26100 264800 26300 265000
rect 26500 264800 26700 265000
rect 26900 264800 27100 265000
rect 27300 264800 27500 265000
rect 27700 264800 27800 265000
rect 19200 248800 19300 249000
rect 19500 248800 19700 249000
rect 19900 248800 20000 249000
rect 19200 248600 20000 248800
rect 19200 248400 19300 248600
rect 19500 248400 19700 248600
rect 19900 248400 20000 248600
rect 19200 248200 20000 248400
rect 19200 248000 19300 248200
rect 19500 248000 19700 248200
rect 19900 248000 20000 248200
rect 19200 247800 20000 248000
rect 19200 247600 19300 247800
rect 19500 247600 19700 247800
rect 19900 247600 20000 247800
rect 19200 247400 20000 247600
rect 19200 247200 19300 247400
rect 19500 247200 19700 247400
rect 19900 247200 20000 247400
rect 19200 247000 20000 247200
rect 19200 246800 19300 247000
rect 19500 246800 19700 247000
rect 19900 246800 20000 247000
rect 19200 246600 20000 246800
rect 19200 246400 19300 246600
rect 19500 246400 19700 246600
rect 19900 246400 20000 246600
rect 19200 246200 20000 246400
rect 19200 246000 19300 246200
rect 19500 246000 19700 246200
rect 19900 246000 20000 246200
rect 19200 245800 20000 246000
rect 19200 245600 19300 245800
rect 19500 245600 19700 245800
rect 19900 245600 20000 245800
rect 19200 245400 20000 245600
rect 19200 245200 19300 245400
rect 19500 245200 19700 245400
rect 19900 245200 20000 245400
rect 19200 245000 20000 245200
rect 19200 244800 19300 245000
rect 19500 244800 19700 245000
rect 19900 244800 20000 245000
rect 19200 244600 20000 244800
rect 19200 244400 19300 244600
rect 19500 244400 19700 244600
rect 19900 244400 20000 244600
rect 22600 249600 27800 264800
rect 44695 265100 45005 265110
rect 44695 264800 44700 265100
rect 45000 264800 45005 265100
rect 44695 264790 45005 264800
rect 44695 264600 45005 264610
rect 44695 264300 44700 264600
rect 45000 264300 45005 264600
rect 44695 264290 45005 264300
rect 44695 264100 45005 264110
rect 44695 263800 44700 264100
rect 45000 263800 45005 264100
rect 44695 263790 45005 263800
rect 44695 263600 45005 263610
rect 44695 263300 44700 263600
rect 45000 263300 45005 263600
rect 44695 263290 45005 263300
rect 44695 263100 45005 263110
rect 44695 262800 44700 263100
rect 45000 262800 45005 263100
rect 44695 262790 45005 262800
rect 44695 262600 45005 262610
rect 44695 262300 44700 262600
rect 45000 262300 45005 262600
rect 44695 262290 45005 262300
rect 44695 262100 45005 262110
rect 44695 261800 44700 262100
rect 45000 261800 45005 262100
rect 44695 261790 45005 261800
rect 44695 261600 45005 261610
rect 44695 261300 44700 261600
rect 45000 261300 45005 261600
rect 44695 261290 45005 261300
rect 44695 261100 45005 261110
rect 44695 260800 44700 261100
rect 45000 260800 45005 261100
rect 44695 260790 45005 260800
rect 272200 249600 277400 340400
rect 22600 244400 277400 249600
rect 19200 244200 20000 244400
rect 9650 241980 11580 242010
rect 9650 241920 9680 241980
rect 9740 241920 9845 241980
rect 9905 241920 10045 241980
rect 10105 241920 10235 241980
rect 10295 241920 10415 241980
rect 10475 241920 10615 241980
rect 10675 241920 10805 241980
rect 10865 241920 10965 241980
rect 11025 241920 11155 241980
rect 11215 241920 11330 241980
rect 11390 241920 11470 241980
rect 11530 241920 11580 241980
rect 9650 241800 11580 241920
rect 9650 241780 9800 241800
rect 10000 241780 10200 241800
rect 10400 241780 10800 241800
rect 11000 241780 11200 241800
rect 11400 241780 11580 241800
rect 16095 242000 16305 242010
rect 16095 241800 16100 242000
rect 16300 241800 16305 242000
rect 16095 241790 16305 241800
rect 9650 241720 9680 241780
rect 9740 241720 9800 241780
rect 10000 241720 10045 241780
rect 10105 241720 10200 241780
rect 10400 241720 10415 241780
rect 10475 241720 10615 241780
rect 10675 241720 10800 241780
rect 11025 241720 11155 241780
rect 11400 241720 11470 241780
rect 11530 241720 11580 241780
rect 9650 241600 9800 241720
rect 10000 241600 10200 241720
rect 10400 241600 10800 241720
rect 11000 241600 11200 241720
rect 11400 241600 11580 241720
rect 9650 241580 11580 241600
rect 9650 241520 9680 241580
rect 9740 241520 9845 241580
rect 9905 241520 10045 241580
rect 10105 241520 10235 241580
rect 10295 241520 10415 241580
rect 10475 241520 10615 241580
rect 10675 241520 10805 241580
rect 10865 241520 10965 241580
rect 11025 241520 11155 241580
rect 11215 241520 11330 241580
rect 11390 241520 11470 241580
rect 11530 241520 11580 241580
rect 9650 241390 11580 241520
rect 16095 241700 16305 241710
rect 16095 241500 16100 241700
rect 16300 241500 16305 241700
rect 16095 241490 16305 241500
rect 9650 241330 9680 241390
rect 9740 241330 9845 241390
rect 9905 241330 10045 241390
rect 10105 241330 10235 241390
rect 10295 241330 10415 241390
rect 10475 241330 10615 241390
rect 10675 241330 10805 241390
rect 10865 241330 10965 241390
rect 11025 241330 11155 241390
rect 11215 241330 11330 241390
rect 11390 241330 11470 241390
rect 11530 241330 11580 241390
rect 9650 241200 11580 241330
rect 9650 241190 9800 241200
rect 10000 241190 10200 241200
rect 10400 241190 10800 241200
rect 11000 241190 11200 241200
rect 11400 241190 11580 241200
rect 16095 241400 16305 241410
rect 16095 241200 16100 241400
rect 16300 241200 16305 241400
rect 16095 241190 16305 241200
rect 9650 241130 9680 241190
rect 9740 241130 9800 241190
rect 10000 241130 10045 241190
rect 10105 241130 10200 241190
rect 10400 241130 10415 241190
rect 10475 241130 10615 241190
rect 10675 241130 10800 241190
rect 11025 241130 11155 241190
rect 11400 241130 11470 241190
rect 11530 241130 11580 241190
rect 9650 241000 9800 241130
rect 10000 241000 10200 241130
rect 10400 241000 10800 241130
rect 11000 241000 11200 241130
rect 11400 241000 11580 241130
rect 9650 240940 9680 241000
rect 9740 240990 11580 241000
rect 9740 240940 9845 240990
rect 9650 240930 9845 240940
rect 9905 240930 10045 240990
rect 10105 240930 10235 240990
rect 10295 240930 10415 240990
rect 10475 240930 10615 240990
rect 10675 240930 10805 240990
rect 10865 240930 10965 240990
rect 11025 240930 11155 240990
rect 11215 240930 11330 240990
rect 11390 240930 11470 240990
rect 11530 240930 11580 240990
rect 9650 240900 11580 240930
rect 16095 241100 16305 241110
rect 16095 240900 16100 241100
rect 16300 240900 16305 241100
rect 16095 240890 16305 240900
rect 0 219688 292200 219800
rect -800 219400 292200 219688
rect -800 219000 285400 219400
rect 285800 219000 286200 219400
rect 286600 219000 287000 219400
rect 287400 219000 287800 219400
rect 288200 219000 288600 219400
rect 289000 219000 289400 219400
rect 289800 219000 292200 219400
rect -800 218800 292200 219000
rect -800 218400 60000 218800
rect 60400 218400 60800 218800
rect 61200 218400 61600 218800
rect 62000 218400 62400 218800
rect 62800 218400 63200 218800
rect 63600 218400 64000 218800
rect 64400 218400 69000 218800
rect 69400 218400 69800 218800
rect 70200 218400 70600 218800
rect 71000 218400 71400 218800
rect 71800 218400 72200 218800
rect 72600 218400 73000 218800
rect 73400 218600 292200 218800
rect 73400 218400 285400 218600
rect -800 218200 285400 218400
rect 285800 218200 286200 218600
rect 286600 218200 287000 218600
rect 287400 218200 287800 218600
rect 288200 218200 288600 218600
rect 289000 218200 289400 218600
rect 289800 218200 292200 218600
rect -800 218000 292200 218200
rect -800 217600 60000 218000
rect 60400 217600 60800 218000
rect 61200 217600 61600 218000
rect 62000 217600 62400 218000
rect 62800 217600 63200 218000
rect 63600 217600 64000 218000
rect 64400 217600 69000 218000
rect 69400 217600 69800 218000
rect 70200 217600 70600 218000
rect 71000 217600 71400 218000
rect 71800 217600 72200 218000
rect 72600 217600 73000 218000
rect 73400 217800 292200 218000
rect 73400 217600 285400 217800
rect -800 217400 285400 217600
rect 285800 217400 286200 217800
rect 286600 217400 287000 217800
rect 287400 217400 287800 217800
rect 288200 217400 288600 217800
rect 289000 217400 289400 217800
rect 289800 217400 292200 217800
rect -800 217200 292200 217400
rect -800 216800 60000 217200
rect 60400 216800 60800 217200
rect 61200 216800 61600 217200
rect 62000 216800 62400 217200
rect 62800 216800 63200 217200
rect 63600 216800 64000 217200
rect 64400 216800 69000 217200
rect 69400 216800 69800 217200
rect 70200 216800 70600 217200
rect 71000 216800 71400 217200
rect 71800 216800 72200 217200
rect 72600 216800 73000 217200
rect 73400 217000 292200 217200
rect 73400 216800 285400 217000
rect -800 216600 285400 216800
rect 285800 216600 286200 217000
rect 286600 216600 287000 217000
rect 287400 216600 287800 217000
rect 288200 216600 288600 217000
rect 289000 216600 289400 217000
rect 289800 216600 292200 217000
rect -800 216400 292200 216600
rect -800 216000 60000 216400
rect 60400 216000 60800 216400
rect 61200 216000 61600 216400
rect 62000 216000 62400 216400
rect 62800 216000 63200 216400
rect 63600 216000 64000 216400
rect 64400 216000 69000 216400
rect 69400 216000 69800 216400
rect 70200 216000 70600 216400
rect 71000 216000 71400 216400
rect 71800 216000 72200 216400
rect 72600 216000 73000 216400
rect 73400 216200 292200 216400
rect 73400 216000 285400 216200
rect -800 215800 285400 216000
rect 285800 215800 286200 216200
rect 286600 215800 287000 216200
rect 287400 215800 287800 216200
rect 288200 215800 288600 216200
rect 289000 215800 289400 216200
rect 289800 215800 292200 216200
rect -800 215600 292200 215800
rect -800 215200 60000 215600
rect 60400 215200 60800 215600
rect 61200 215200 61600 215600
rect 62000 215200 62400 215600
rect 62800 215200 63200 215600
rect 63600 215200 64000 215600
rect 64400 215200 69000 215600
rect 69400 215200 69800 215600
rect 70200 215200 70600 215600
rect 71000 215200 71400 215600
rect 71800 215200 72200 215600
rect 72600 215200 73000 215600
rect 73400 215400 292200 215600
rect 73400 215200 285400 215400
rect -800 215000 285400 215200
rect 285800 215000 286200 215400
rect 286600 215000 287000 215400
rect 287400 215000 287800 215400
rect 288200 215000 288600 215400
rect 289000 215000 289400 215400
rect 289800 215000 292200 215400
rect -800 214888 292200 215000
rect 0 214800 292200 214888
rect 0 214400 60000 214800
rect 60400 214400 60800 214800
rect 61200 214400 61600 214800
rect 62000 214400 62400 214800
rect 62800 214400 63200 214800
rect 63600 214400 64000 214800
rect 64400 214400 69000 214800
rect 69400 214400 69800 214800
rect 70200 214400 70600 214800
rect 71000 214400 71400 214800
rect 71800 214400 72200 214800
rect 72600 214400 73000 214800
rect 73400 214600 292200 214800
rect 73400 214400 285200 214600
rect 0 214200 285200 214400
rect 285600 214200 286000 214600
rect 286400 214200 286800 214600
rect 287200 214200 287600 214600
rect 288000 214200 288400 214600
rect 288800 214200 289200 214600
rect 289600 214200 292200 214600
rect 0 213800 292200 214200
rect 0 213400 285200 213800
rect 285600 213400 286000 213800
rect 286400 213400 286800 213800
rect 287200 213400 287600 213800
rect 288000 213400 288400 213800
rect 288800 213400 289200 213800
rect 289600 213400 292200 213800
rect 0 213000 292200 213400
rect 0 212600 285200 213000
rect 285600 212600 286000 213000
rect 286400 212600 286800 213000
rect 287200 212600 287600 213000
rect 288000 212600 288400 213000
rect 288800 212600 289200 213000
rect 289600 212600 292200 213000
rect 0 212200 292200 212600
rect 0 211800 285200 212200
rect 285600 211800 286000 212200
rect 286400 211800 286800 212200
rect 287200 211800 287600 212200
rect 288000 211800 288400 212200
rect 288800 211800 289200 212200
rect 289600 211800 292200 212200
rect 0 211400 292200 211800
rect 0 211000 285200 211400
rect 285600 211000 286000 211400
rect 286400 211000 286800 211400
rect 287200 211000 287600 211400
rect 288000 211000 288400 211400
rect 288800 211000 289200 211400
rect 289600 211000 292200 211400
rect 0 210600 292200 211000
rect 0 210200 285200 210600
rect 285600 210200 286000 210600
rect 286400 210200 286800 210600
rect 287200 210200 287600 210600
rect 288000 210200 288400 210600
rect 288800 210200 289200 210600
rect 289600 210200 292200 210600
rect 0 210000 69000 210200
rect 0 209688 60000 210000
rect -800 209600 60000 209688
rect 60400 209600 60800 210000
rect 61200 209600 61600 210000
rect 62000 209600 62400 210000
rect 62800 209600 63200 210000
rect 63600 209600 64000 210000
rect 64400 209800 69000 210000
rect 69400 209800 69800 210200
rect 70200 209800 70600 210200
rect 71000 209800 71400 210200
rect 71800 209800 72200 210200
rect 72600 209800 73000 210200
rect 73400 209800 292200 210200
rect 64400 209600 285200 209800
rect -800 209400 285200 209600
rect 285600 209400 286000 209800
rect 286400 209400 286800 209800
rect 287200 209400 287600 209800
rect 288000 209400 288400 209800
rect 288800 209400 289200 209800
rect 289600 209400 292200 209800
rect -800 209200 69000 209400
rect -800 208800 60000 209200
rect 60400 208800 60800 209200
rect 61200 208800 61600 209200
rect 62000 208800 62400 209200
rect 62800 208800 63200 209200
rect 63600 208800 64000 209200
rect 64400 209000 69000 209200
rect 69400 209000 69800 209400
rect 70200 209000 70600 209400
rect 71000 209000 71400 209400
rect 71800 209000 72200 209400
rect 72600 209000 73000 209400
rect 73400 209000 292200 209400
rect 64400 208800 285200 209000
rect -800 208600 285200 208800
rect 285600 208600 286000 209000
rect 286400 208600 286800 209000
rect 287200 208600 287600 209000
rect 288000 208600 288400 209000
rect 288800 208600 289200 209000
rect 289600 208600 292200 209000
rect -800 208400 69000 208600
rect -800 208000 60000 208400
rect 60400 208000 60800 208400
rect 61200 208000 61600 208400
rect 62000 208000 62400 208400
rect 62800 208000 63200 208400
rect 63600 208000 64000 208400
rect 64400 208200 69000 208400
rect 69400 208200 69800 208600
rect 70200 208200 70600 208600
rect 71000 208200 71400 208600
rect 71800 208200 72200 208600
rect 72600 208200 73000 208600
rect 73400 208200 292200 208600
rect 64400 208000 285200 208200
rect -800 207800 285200 208000
rect 285600 207800 286000 208200
rect 286400 207800 286800 208200
rect 287200 207800 287600 208200
rect 288000 207800 288400 208200
rect 288800 207800 289200 208200
rect 289600 207800 292200 208200
rect -800 207600 69000 207800
rect -800 207200 60000 207600
rect 60400 207200 60800 207600
rect 61200 207200 61600 207600
rect 62000 207200 62400 207600
rect 62800 207200 63200 207600
rect 63600 207200 64000 207600
rect 64400 207400 69000 207600
rect 69400 207400 69800 207800
rect 70200 207400 70600 207800
rect 71000 207400 71400 207800
rect 71800 207400 72200 207800
rect 72600 207400 73000 207800
rect 73400 207400 292200 207800
rect 64400 207200 285200 207400
rect -800 207000 285200 207200
rect 285600 207000 286000 207400
rect 286400 207000 286800 207400
rect 287200 207000 287600 207400
rect 288000 207000 288400 207400
rect 288800 207000 289200 207400
rect 289600 207000 292200 207400
rect -800 206800 69000 207000
rect -800 206400 60000 206800
rect 60400 206400 60800 206800
rect 61200 206400 61600 206800
rect 62000 206400 62400 206800
rect 62800 206400 63200 206800
rect 63600 206400 64000 206800
rect 64400 206600 69000 206800
rect 69400 206600 69800 207000
rect 70200 206600 70600 207000
rect 71000 206600 71400 207000
rect 71800 206600 72200 207000
rect 72600 206600 73000 207000
rect 73400 206600 292200 207000
rect 64400 206400 285200 206600
rect -800 206200 285200 206400
rect 285600 206200 286000 206600
rect 286400 206200 286800 206600
rect 287200 206200 287600 206600
rect 288000 206200 288400 206600
rect 288800 206200 289200 206600
rect 289600 206200 292200 206600
rect -800 206000 69000 206200
rect -800 205600 60000 206000
rect 60400 205600 60800 206000
rect 61200 205600 61600 206000
rect 62000 205600 62400 206000
rect 62800 205600 63200 206000
rect 63600 205600 64000 206000
rect 64400 205800 69000 206000
rect 69400 205800 69800 206200
rect 70200 205800 70600 206200
rect 71000 205800 71400 206200
rect 71800 205800 72200 206200
rect 72600 205800 73000 206200
rect 73400 205800 292200 206200
rect 64400 205600 285200 205800
rect -800 205400 285200 205600
rect 285600 205400 286000 205800
rect 286400 205400 286800 205800
rect 287200 205400 287600 205800
rect 288000 205400 288400 205800
rect 288800 205400 289200 205800
rect 289600 205400 292200 205800
rect -800 204888 292200 205400
rect 0 204800 292200 204888
rect 0 177688 11600 177900
rect -800 172888 11600 177688
rect 0 167688 11600 172888
rect -800 162888 11600 167688
rect 0 162800 11600 162888
rect 13600 177600 306000 177900
rect 13600 177200 86000 177600
rect 86400 177200 86800 177600
rect 87200 177200 87600 177600
rect 88000 177200 88400 177600
rect 88800 177200 89200 177600
rect 89600 177200 90000 177600
rect 90400 177200 299400 177600
rect 299800 177200 300200 177600
rect 300600 177200 301000 177600
rect 301400 177200 301800 177600
rect 302200 177200 302600 177600
rect 303000 177200 303400 177600
rect 303800 177200 306000 177600
rect 13600 176800 306000 177200
rect 13600 176400 86000 176800
rect 86400 176400 86800 176800
rect 87200 176400 87600 176800
rect 88000 176400 88400 176800
rect 88800 176400 89200 176800
rect 89600 176400 90000 176800
rect 90400 176400 299400 176800
rect 299800 176400 300200 176800
rect 300600 176400 301000 176800
rect 301400 176400 301800 176800
rect 302200 176400 302600 176800
rect 303000 176400 303400 176800
rect 303800 176400 306000 176800
rect 13600 176000 306000 176400
rect 13600 175600 86000 176000
rect 86400 175600 86800 176000
rect 87200 175600 87600 176000
rect 88000 175600 88400 176000
rect 88800 175600 89200 176000
rect 89600 175600 90000 176000
rect 90400 175600 299400 176000
rect 299800 175600 300200 176000
rect 300600 175600 301000 176000
rect 301400 175600 301800 176000
rect 302200 175600 302600 176000
rect 303000 175600 303400 176000
rect 303800 175600 306000 176000
rect 13600 175200 306000 175600
rect 13600 174800 86000 175200
rect 86400 174800 86800 175200
rect 87200 174800 87600 175200
rect 88000 174800 88400 175200
rect 88800 174800 89200 175200
rect 89600 174800 90000 175200
rect 90400 174800 299400 175200
rect 299800 174800 300200 175200
rect 300600 174800 301000 175200
rect 301400 174800 301800 175200
rect 302200 174800 302600 175200
rect 303000 174800 303400 175200
rect 303800 174800 306000 175200
rect 13600 174400 306000 174800
rect 13600 174000 86000 174400
rect 86400 174000 86800 174400
rect 87200 174000 87600 174400
rect 88000 174000 88400 174400
rect 88800 174000 89200 174400
rect 89600 174000 90000 174400
rect 90400 174000 299400 174400
rect 299800 174000 300200 174400
rect 300600 174000 301000 174400
rect 301400 174000 301800 174400
rect 302200 174000 302600 174400
rect 303000 174000 303400 174400
rect 303800 174000 306000 174400
rect 13600 173600 306000 174000
rect 13600 173200 86000 173600
rect 86400 173200 86800 173600
rect 87200 173200 87600 173600
rect 88000 173200 88400 173600
rect 88800 173200 89200 173600
rect 89600 173200 90000 173600
rect 90400 173200 299400 173600
rect 299800 173200 300200 173600
rect 300600 173200 301000 173600
rect 301400 173200 301800 173600
rect 302200 173200 302600 173600
rect 303000 173200 303400 173600
rect 303800 173200 306000 173600
rect 13600 172800 306000 173200
rect 13600 172400 86000 172800
rect 86400 172400 86800 172800
rect 87200 172400 87600 172800
rect 88000 172400 88400 172800
rect 88800 172400 89200 172800
rect 89600 172400 90000 172800
rect 90400 172400 299400 172800
rect 299800 172400 300200 172800
rect 300600 172400 301000 172800
rect 301400 172400 301800 172800
rect 302200 172400 302600 172800
rect 303000 172400 303400 172800
rect 303800 172400 306000 172800
rect 13600 172000 306000 172400
rect 13600 171600 86000 172000
rect 86400 171600 86800 172000
rect 87200 171600 87600 172000
rect 88000 171600 88400 172000
rect 88800 171600 89200 172000
rect 89600 171600 90000 172000
rect 90400 171600 299400 172000
rect 299800 171600 300200 172000
rect 300600 171600 301000 172000
rect 301400 171600 301800 172000
rect 302200 171600 302600 172000
rect 303000 171600 303400 172000
rect 303800 171600 306000 172000
rect 13600 171200 306000 171600
rect 13600 170800 86000 171200
rect 86400 170800 86800 171200
rect 87200 170800 87600 171200
rect 88000 170800 88400 171200
rect 88800 170800 89200 171200
rect 89600 170800 90000 171200
rect 90400 170800 299400 171200
rect 299800 170800 300200 171200
rect 300600 170800 301000 171200
rect 301400 170800 301800 171200
rect 302200 170800 302600 171200
rect 303000 170800 303400 171200
rect 303800 170800 306000 171200
rect 13600 170400 306000 170800
rect 13600 170000 86000 170400
rect 86400 170000 86800 170400
rect 87200 170000 87600 170400
rect 88000 170000 88400 170400
rect 88800 170000 89200 170400
rect 89600 170000 90000 170400
rect 90400 170000 299400 170400
rect 299800 170000 300200 170400
rect 300600 170000 301000 170400
rect 301400 170000 301800 170400
rect 302200 170000 302600 170400
rect 303000 170000 303400 170400
rect 303800 170000 306000 170400
rect 13600 169600 306000 170000
rect 13600 169200 86000 169600
rect 86400 169200 86800 169600
rect 87200 169200 87600 169600
rect 88000 169200 88400 169600
rect 88800 169200 89200 169600
rect 89600 169200 90000 169600
rect 90400 169200 299400 169600
rect 299800 169200 300200 169600
rect 300600 169200 301000 169600
rect 301400 169200 301800 169600
rect 302200 169200 302600 169600
rect 303000 169200 303400 169600
rect 303800 169200 306000 169600
rect 13600 168800 306000 169200
rect 13600 168400 86000 168800
rect 86400 168400 86800 168800
rect 87200 168400 87600 168800
rect 88000 168400 88400 168800
rect 88800 168400 89200 168800
rect 89600 168400 90000 168800
rect 90400 168400 299400 168800
rect 299800 168400 300200 168800
rect 300600 168400 301000 168800
rect 301400 168400 301800 168800
rect 302200 168400 302600 168800
rect 303000 168400 303400 168800
rect 303800 168400 306000 168800
rect 13600 168000 306000 168400
rect 13600 167600 86000 168000
rect 86400 167600 86800 168000
rect 87200 167600 87600 168000
rect 88000 167600 88400 168000
rect 88800 167600 89200 168000
rect 89600 167600 90000 168000
rect 90400 167600 299400 168000
rect 299800 167600 300200 168000
rect 300600 167600 301000 168000
rect 301400 167600 301800 168000
rect 302200 167600 302600 168000
rect 303000 167600 303400 168000
rect 303800 167600 306000 168000
rect 13600 167200 306000 167600
rect 13600 166800 86000 167200
rect 86400 166800 86800 167200
rect 87200 166800 87600 167200
rect 88000 166800 88400 167200
rect 88800 166800 89200 167200
rect 89600 166800 90000 167200
rect 90400 166800 299400 167200
rect 299800 166800 300200 167200
rect 300600 166800 301000 167200
rect 301400 166800 301800 167200
rect 302200 166800 302600 167200
rect 303000 166800 303400 167200
rect 303800 166800 306000 167200
rect 13600 166400 306000 166800
rect 13600 166000 86000 166400
rect 86400 166000 86800 166400
rect 87200 166000 87600 166400
rect 88000 166000 88400 166400
rect 88800 166000 89200 166400
rect 89600 166000 90000 166400
rect 90400 166000 299400 166400
rect 299800 166000 300200 166400
rect 300600 166000 301000 166400
rect 301400 166000 301800 166400
rect 302200 166000 302600 166400
rect 303000 166000 303400 166400
rect 303800 166000 306000 166400
rect 13600 165600 306000 166000
rect 13600 165200 86000 165600
rect 86400 165200 86800 165600
rect 87200 165200 87600 165600
rect 88000 165200 88400 165600
rect 88800 165200 89200 165600
rect 89600 165200 90000 165600
rect 90400 165200 299400 165600
rect 299800 165200 300200 165600
rect 300600 165200 301000 165600
rect 301400 165200 301800 165600
rect 302200 165200 302600 165600
rect 303000 165200 303400 165600
rect 303800 165200 306000 165600
rect 13600 164800 306000 165200
rect 13600 164400 86000 164800
rect 86400 164400 86800 164800
rect 87200 164400 87600 164800
rect 88000 164400 88400 164800
rect 88800 164400 89200 164800
rect 89600 164400 90000 164800
rect 90400 164400 299400 164800
rect 299800 164400 300200 164800
rect 300600 164400 301000 164800
rect 301400 164400 301800 164800
rect 302200 164400 302600 164800
rect 303000 164400 303400 164800
rect 303800 164400 306000 164800
rect 13600 164000 306000 164400
rect 13600 163600 86000 164000
rect 86400 163600 86800 164000
rect 87200 163600 87600 164000
rect 88000 163600 88400 164000
rect 88800 163600 89200 164000
rect 89600 163600 90000 164000
rect 90400 163600 299400 164000
rect 299800 163600 300200 164000
rect 300600 163600 301000 164000
rect 301400 163600 301800 164000
rect 302200 163600 302600 164000
rect 303000 163600 303400 164000
rect 303800 163600 306000 164000
rect 13600 162800 306000 163600
rect 311800 129600 317000 342100
rect 0 124888 317000 129600
rect -800 124776 317000 124888
rect 0 124400 317000 124776
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 318000 86300 323200 345500
rect 0 81666 323200 86300
rect -800 81554 323200 81666
rect 0 80900 323200 81554
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 324200 42900 329400 347200
rect 330400 284500 335600 348900
rect 336600 291100 341800 350600
rect 342800 297500 348000 352400
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 564800 313764 584000 314200
rect 564800 313652 584800 313764
rect 564800 311800 584000 313652
rect 564800 308000 567200 311800
rect 556300 306120 561120 306400
rect 556300 306020 559840 306120
rect 559940 306020 559980 306120
rect 560080 306020 560120 306120
rect 560220 306020 560260 306120
rect 560360 306020 560400 306120
rect 560500 306020 560540 306120
rect 560640 306020 560680 306120
rect 560780 306020 560820 306120
rect 560920 306020 560960 306120
rect 561060 306020 561120 306120
rect 556300 305980 561120 306020
rect 556300 305880 559840 305980
rect 559940 305880 559980 305980
rect 560080 305880 560120 305980
rect 560220 305880 560260 305980
rect 560360 305880 560400 305980
rect 560500 305880 560540 305980
rect 560640 305880 560680 305980
rect 560780 305880 560820 305980
rect 560920 305880 560960 305980
rect 561060 305880 561120 305980
rect 556300 305800 561120 305880
rect 562200 306280 568000 308000
rect 562200 306240 570140 306280
rect 562200 306140 569280 306240
rect 569380 306140 569420 306240
rect 569520 306140 569560 306240
rect 569660 306140 569700 306240
rect 569800 306140 569840 306240
rect 569940 306140 569980 306240
rect 570080 306140 570140 306240
rect 562200 305980 570140 306140
rect 562200 305880 569280 305980
rect 569380 305880 569420 305980
rect 569520 305880 569560 305980
rect 569660 305880 569700 305980
rect 569800 305880 569840 305980
rect 569940 305880 569980 305980
rect 570080 305880 570140 305980
rect 562200 305840 570140 305880
rect 556300 301600 557600 305800
rect 562200 302160 568000 305840
rect 511500 301400 557600 301600
rect 511500 301200 511700 301400
rect 511900 301200 512100 301400
rect 512300 301200 512500 301400
rect 512700 301200 512900 301400
rect 513100 301200 513300 301400
rect 513500 301200 513700 301400
rect 513900 301200 514100 301400
rect 514300 301200 514500 301400
rect 514700 301200 514900 301400
rect 515100 301200 515300 301400
rect 515500 301200 515700 301400
rect 515900 301200 516100 301400
rect 516300 301200 516500 301400
rect 516700 301200 557600 301400
rect 511500 301000 557600 301200
rect 511500 300800 511700 301000
rect 511900 300800 512100 301000
rect 512300 300800 512500 301000
rect 512700 300800 512900 301000
rect 513100 300800 513300 301000
rect 513500 300800 513700 301000
rect 513900 300800 514100 301000
rect 514300 300800 514500 301000
rect 514700 300800 514900 301000
rect 515100 300800 515300 301000
rect 515500 300800 515700 301000
rect 515900 300800 516100 301000
rect 516300 300800 516500 301000
rect 516700 300800 557600 301000
rect 511500 300600 557600 300800
rect 511500 300400 511700 300600
rect 511900 300400 512100 300600
rect 512300 300400 512500 300600
rect 512700 300400 512900 300600
rect 513100 300400 513300 300600
rect 513500 300400 513700 300600
rect 513900 300400 514100 300600
rect 514300 300400 514500 300600
rect 514700 300400 514900 300600
rect 515100 300400 515300 300600
rect 515500 300400 515700 300600
rect 515900 300400 516100 300600
rect 516300 300400 516500 300600
rect 516700 300400 557600 300600
rect 511500 300000 557600 300400
rect 559800 302120 568000 302160
rect 559800 302060 559940 302120
rect 560000 302060 560130 302120
rect 560190 302060 560330 302120
rect 560390 302060 560520 302120
rect 560580 302060 560720 302120
rect 560780 302060 560920 302120
rect 560980 302060 568000 302120
rect 559800 301955 568000 302060
rect 559800 301895 559930 301955
rect 559990 301895 560130 301955
rect 560190 301895 560330 301955
rect 560390 301895 560520 301955
rect 560580 301895 560720 301955
rect 560780 301895 560920 301955
rect 560980 301895 568000 301955
rect 559800 301755 568000 301895
rect 559800 301695 559930 301755
rect 559990 301695 560130 301755
rect 560190 301695 560330 301755
rect 560390 301695 560520 301755
rect 560580 301695 560720 301755
rect 560780 301695 560920 301755
rect 560980 301695 568000 301755
rect 559800 301565 568000 301695
rect 559800 301505 559930 301565
rect 559990 301505 560130 301565
rect 560190 301505 560330 301565
rect 560390 301505 560520 301565
rect 560580 301505 560720 301565
rect 560780 301505 560920 301565
rect 560980 301505 568000 301565
rect 559800 301385 568000 301505
rect 559800 301325 559930 301385
rect 559990 301325 560130 301385
rect 560190 301325 560330 301385
rect 560390 301325 560520 301385
rect 560580 301325 560720 301385
rect 560780 301325 560920 301385
rect 560980 301325 568000 301385
rect 559800 301185 568000 301325
rect 559800 301125 559930 301185
rect 559990 301125 560130 301185
rect 560190 301125 560330 301185
rect 560390 301125 560520 301185
rect 560580 301125 560720 301185
rect 560780 301125 560920 301185
rect 560980 301125 568000 301185
rect 559800 300995 568000 301125
rect 559800 300935 559930 300995
rect 559990 300935 560130 300995
rect 560190 300935 560330 300995
rect 560390 300935 560520 300995
rect 560580 300935 560720 300995
rect 560780 300935 560920 300995
rect 560980 300935 568000 300995
rect 559800 300835 568000 300935
rect 559800 300775 559930 300835
rect 559990 300775 560130 300835
rect 560190 300775 560330 300835
rect 560390 300775 560520 300835
rect 560580 300775 560720 300835
rect 560780 300775 560920 300835
rect 560980 300775 568000 300835
rect 559800 300645 568000 300775
rect 559800 300585 559930 300645
rect 559990 300585 560130 300645
rect 560190 300585 560330 300645
rect 560390 300585 560520 300645
rect 560580 300585 560720 300645
rect 560780 300585 560920 300645
rect 560980 300585 568000 300645
rect 559800 300470 568000 300585
rect 559800 300410 559930 300470
rect 559990 300410 560130 300470
rect 560190 300410 560330 300470
rect 560390 300410 560520 300470
rect 560580 300410 560720 300470
rect 560780 300410 560920 300470
rect 560980 300410 568000 300470
rect 559800 300330 568000 300410
rect 559800 300270 559930 300330
rect 559990 300270 560130 300330
rect 560190 300270 560330 300330
rect 560390 300270 560520 300330
rect 560580 300270 560720 300330
rect 560780 300270 560920 300330
rect 560980 300270 568000 300330
rect 559800 300220 568000 300270
rect 530609 298992 531049 299042
rect 530609 298862 530639 298992
rect 530739 298862 530899 298992
rect 530999 298862 531049 298992
rect 550109 298992 550539 299052
rect 342800 294400 530300 297500
rect 342800 294200 528300 294400
rect 528500 294200 528700 294400
rect 528900 294200 529100 294400
rect 529300 294200 529500 294400
rect 529700 294200 529900 294400
rect 530100 294200 530300 294400
rect 342800 294100 530300 294200
rect 342800 293900 528300 294100
rect 528500 293900 528700 294100
rect 528900 293900 529100 294100
rect 529300 293900 529500 294100
rect 529700 293900 529900 294100
rect 530100 293900 530300 294100
rect 342800 293700 530300 293900
rect 342800 293500 528300 293700
rect 528500 293500 528700 293700
rect 528900 293500 529100 293700
rect 529300 293500 529500 293700
rect 529700 293500 529900 293700
rect 530100 293500 530300 293700
rect 342800 293300 530300 293500
rect 342800 293100 528300 293300
rect 528500 293100 528700 293300
rect 528900 293100 529100 293300
rect 529300 293100 529500 293300
rect 529700 293100 529900 293300
rect 530100 293100 530300 293300
rect 342800 292900 530300 293100
rect 342800 292700 528300 292900
rect 528500 292700 528700 292900
rect 528900 292700 529100 292900
rect 529300 292700 529500 292900
rect 529700 292700 529900 292900
rect 530100 292700 530300 292900
rect 342800 292300 530300 292700
rect 530609 292132 531049 298862
rect 533169 298921 536569 298941
rect 533169 298857 533197 298921
rect 536541 298857 536569 298921
rect 533169 295442 536569 298857
rect 536969 298921 540369 298941
rect 536969 298857 536997 298921
rect 540341 298857 540369 298921
rect 536969 295442 540369 298857
rect 540769 298921 544169 298941
rect 540769 298857 540797 298921
rect 544141 298857 544169 298921
rect 540769 295442 544169 298857
rect 544569 298921 547969 298941
rect 544569 298857 544597 298921
rect 547941 298857 547969 298921
rect 544569 295442 547969 298857
rect 550109 298862 550129 298992
rect 550239 298862 550389 298992
rect 550499 298862 550539 298992
rect 535919 294972 547499 295212
rect 535919 294962 542919 294972
rect 535919 294892 537969 294962
rect 538059 294892 538139 294962
rect 538229 294892 540459 294962
rect 540549 294892 540629 294962
rect 540719 294892 542919 294962
rect 542999 294892 543089 294972
rect 543169 294892 547499 294972
rect 535919 294852 547499 294892
rect 537069 294682 537339 294702
rect 537069 294602 537089 294682
rect 537169 294602 537239 294682
rect 537319 294602 537339 294682
rect 537069 294582 537339 294602
rect 539559 294682 539829 294692
rect 539559 294602 539579 294682
rect 539659 294602 539729 294682
rect 539809 294602 539829 294682
rect 539559 294582 539829 294602
rect 542039 294682 542309 294702
rect 542039 294602 542059 294682
rect 542139 294602 542209 294682
rect 542289 294602 542309 294682
rect 542039 294582 542309 294602
rect 537069 294142 537339 294162
rect 537069 294062 537089 294142
rect 537169 294062 537239 294142
rect 537319 294062 537339 294142
rect 537069 294042 537339 294062
rect 539559 294142 539829 294152
rect 539559 294062 539579 294142
rect 539659 294062 539729 294142
rect 539809 294062 539829 294142
rect 539559 294042 539829 294062
rect 542039 294142 542309 294162
rect 542039 294062 542059 294142
rect 542139 294062 542209 294142
rect 542289 294062 542309 294142
rect 542039 294042 542309 294062
rect 547089 293982 547499 294852
rect 535679 293922 547499 293982
rect 535679 293912 540619 293922
rect 535679 293842 537979 293912
rect 538069 293842 538119 293912
rect 538209 293842 540459 293912
rect 540549 293852 540619 293912
rect 540709 293852 542919 293922
rect 542999 293852 543089 293922
rect 543169 293852 547499 293922
rect 540549 293842 547499 293852
rect 535679 293752 547499 293842
rect 537069 293602 537339 293632
rect 537069 293522 537089 293602
rect 537169 293522 537239 293602
rect 537319 293522 537339 293602
rect 537069 293502 537339 293522
rect 539559 293602 539829 293612
rect 539559 293522 539579 293602
rect 539659 293522 539729 293602
rect 539809 293522 539829 293602
rect 539559 293502 539829 293522
rect 542039 293602 542309 293632
rect 542039 293522 542069 293602
rect 542149 293522 542209 293602
rect 542289 293522 542309 293602
rect 542039 293502 542309 293522
rect 547089 293392 547499 293752
rect 536069 293382 547499 293392
rect 536069 293302 537979 293382
rect 538059 293302 538149 293382
rect 538229 293302 540459 293382
rect 540539 293302 540629 293382
rect 540709 293302 542919 293382
rect 542999 293302 543089 293382
rect 543169 293302 547499 293382
rect 536069 293172 547499 293302
rect 538359 293002 538589 293022
rect 538359 292922 538379 293002
rect 538459 292922 538489 293002
rect 538569 292922 538589 293002
rect 538359 292892 538589 292922
rect 540769 293002 540999 293022
rect 540769 292922 540789 293002
rect 540869 292922 540899 293002
rect 540979 292922 540999 293002
rect 540769 292912 540999 292922
rect 543229 292992 543459 293002
rect 543229 292912 543249 292992
rect 543329 292912 543359 292992
rect 543439 292912 543459 292992
rect 543229 292892 543459 292912
rect 540769 292412 540999 292422
rect 538359 292392 538589 292402
rect 538359 292312 538379 292392
rect 538459 292312 538489 292392
rect 538569 292312 538589 292392
rect 540769 292332 540789 292412
rect 540869 292332 540899 292412
rect 540979 292332 540999 292412
rect 540769 292312 540999 292332
rect 543229 292412 543459 292422
rect 543229 292332 543249 292412
rect 543329 292332 543359 292412
rect 543439 292332 543459 292412
rect 543229 292312 543459 292332
rect 538359 292302 538589 292312
rect 547089 292232 547499 293172
rect 530609 291992 530629 292132
rect 530759 291992 530879 292132
rect 531009 291992 531049 292132
rect 535989 292222 547499 292232
rect 535989 292142 537979 292222
rect 538069 292142 538139 292222
rect 538229 292212 547499 292222
rect 538229 292142 540459 292212
rect 540539 292142 540629 292212
rect 540709 292142 542919 292212
rect 542999 292142 543089 292212
rect 543169 292142 547499 292212
rect 550109 292302 550539 298862
rect 562200 295100 568000 300220
rect 569100 302120 570220 302180
rect 569100 302060 569140 302120
rect 569200 302060 569330 302120
rect 569390 302060 569530 302120
rect 569590 302060 569720 302120
rect 569780 302060 569920 302120
rect 569980 302060 570120 302120
rect 570180 302060 570220 302120
rect 569100 302000 570220 302060
rect 569100 301955 569300 302000
rect 569500 301955 569800 302000
rect 570000 301955 570220 302000
rect 569100 301895 569130 301955
rect 569190 301895 569300 301955
rect 569500 301895 569530 301955
rect 569590 301895 569720 301955
rect 569780 301895 569800 301955
rect 570000 301895 570120 301955
rect 570180 301895 570220 301955
rect 569100 301800 569300 301895
rect 569500 301800 569800 301895
rect 570000 301800 570220 301895
rect 569100 301755 570220 301800
rect 569100 301695 569130 301755
rect 569190 301695 569330 301755
rect 569390 301695 569530 301755
rect 569590 301695 569720 301755
rect 569780 301695 569920 301755
rect 569980 301695 570120 301755
rect 570180 301695 570220 301755
rect 569100 301600 570220 301695
rect 569100 301565 569300 301600
rect 569500 301565 569800 301600
rect 570000 301565 570220 301600
rect 569100 301505 569130 301565
rect 569190 301505 569300 301565
rect 569500 301505 569530 301565
rect 569590 301505 569720 301565
rect 569780 301505 569800 301565
rect 570000 301505 570120 301565
rect 570180 301505 570220 301565
rect 569100 301400 569300 301505
rect 569500 301400 569800 301505
rect 570000 301400 570220 301505
rect 569100 301385 570220 301400
rect 569100 301325 569130 301385
rect 569190 301325 569330 301385
rect 569390 301325 569530 301385
rect 569590 301325 569720 301385
rect 569780 301325 569920 301385
rect 569980 301325 570120 301385
rect 570180 301325 570220 301385
rect 569100 301200 570220 301325
rect 569100 301185 569300 301200
rect 569500 301185 569800 301200
rect 570000 301185 570220 301200
rect 569100 301125 569130 301185
rect 569190 301125 569300 301185
rect 569500 301125 569530 301185
rect 569590 301125 569720 301185
rect 569780 301125 569800 301185
rect 570000 301125 570120 301185
rect 570180 301125 570220 301185
rect 569100 301000 569300 301125
rect 569500 301000 569800 301125
rect 570000 301000 570220 301125
rect 569100 300995 570220 301000
rect 569100 300935 569130 300995
rect 569190 300935 569330 300995
rect 569390 300935 569530 300995
rect 569590 300935 569720 300995
rect 569780 300935 569920 300995
rect 569980 300935 570120 300995
rect 570180 300935 570220 300995
rect 569100 300835 570220 300935
rect 569100 300775 569130 300835
rect 569190 300800 569330 300835
rect 569390 300800 569530 300835
rect 569190 300775 569300 300800
rect 569500 300775 569530 300800
rect 569590 300775 569720 300835
rect 569780 300800 569920 300835
rect 569980 300800 570120 300835
rect 569780 300775 569800 300800
rect 570000 300775 570120 300800
rect 570180 300775 570220 300835
rect 569100 300645 569300 300775
rect 569500 300645 569800 300775
rect 570000 300645 570220 300775
rect 569100 300585 569130 300645
rect 569190 300600 569300 300645
rect 569500 300600 569530 300645
rect 569190 300585 569330 300600
rect 569390 300585 569530 300600
rect 569590 300585 569720 300645
rect 569780 300600 569800 300645
rect 570000 300600 570120 300645
rect 569780 300585 569920 300600
rect 569980 300585 570120 300600
rect 570180 300585 570220 300645
rect 569100 300470 570220 300585
rect 569100 300410 569130 300470
rect 569190 300410 569330 300470
rect 569390 300410 569530 300470
rect 569590 300410 569720 300470
rect 569780 300410 569920 300470
rect 569980 300410 570120 300470
rect 570180 300410 570220 300470
rect 569100 300400 570220 300410
rect 569100 300330 569300 300400
rect 569500 300330 569800 300400
rect 570000 300330 570220 300400
rect 569100 300270 569130 300330
rect 569190 300270 569300 300330
rect 569500 300270 569530 300330
rect 569590 300270 569720 300330
rect 569780 300270 569800 300330
rect 570000 300270 570120 300330
rect 570180 300270 570220 300330
rect 569100 300200 569300 300270
rect 569500 300200 569800 300270
rect 570000 300200 570220 300270
rect 569100 300100 570220 300200
rect 562200 294900 562300 295100
rect 562500 294900 562700 295100
rect 562900 294900 563100 295100
rect 563300 294900 563500 295100
rect 563700 294900 563900 295100
rect 564100 294900 564300 295100
rect 564500 294900 564700 295100
rect 564900 294900 565100 295100
rect 565300 294900 565500 295100
rect 565700 294900 565900 295100
rect 566100 294900 566300 295100
rect 566500 294900 566700 295100
rect 566900 294900 567100 295100
rect 567300 294900 567500 295100
rect 567700 294900 568000 295100
rect 562200 294700 568000 294900
rect 562200 294500 562300 294700
rect 562500 294500 562700 294700
rect 562900 294500 563100 294700
rect 563300 294500 563500 294700
rect 563700 294500 563900 294700
rect 564100 294500 564300 294700
rect 564500 294500 564700 294700
rect 564900 294500 565100 294700
rect 565300 294500 565500 294700
rect 565700 294500 565900 294700
rect 566100 294500 566300 294700
rect 566500 294500 566700 294700
rect 566900 294500 567100 294700
rect 567300 294500 567500 294700
rect 567700 294500 568000 294700
rect 562200 294300 568000 294500
rect 562200 294100 562300 294300
rect 562500 294100 562700 294300
rect 562900 294100 563100 294300
rect 563300 294100 563500 294300
rect 563700 294100 563900 294300
rect 564100 294100 564300 294300
rect 564500 294100 564700 294300
rect 564900 294100 565100 294300
rect 565300 294100 565500 294300
rect 565700 294100 565900 294300
rect 566100 294100 566300 294300
rect 566500 294100 566700 294300
rect 566900 294100 567100 294300
rect 567300 294100 567500 294300
rect 567700 294100 568000 294300
rect 562200 293900 568000 294100
rect 562200 293700 562300 293900
rect 562500 293700 562700 293900
rect 562900 293700 563100 293900
rect 563300 293700 563500 293900
rect 563700 293700 563900 293900
rect 564100 293700 564300 293900
rect 564500 293700 564700 293900
rect 564900 293700 565100 293900
rect 565300 293700 565500 293900
rect 565700 293700 565900 293900
rect 566100 293700 566300 293900
rect 566500 293700 566700 293900
rect 566900 293700 567100 293900
rect 567300 293700 567500 293900
rect 567700 293700 568000 293900
rect 562200 293500 568000 293700
rect 562200 293300 562300 293500
rect 562500 293300 562700 293500
rect 562900 293300 563100 293500
rect 563300 293300 563500 293500
rect 563700 293300 563900 293500
rect 564100 293300 564300 293500
rect 564500 293300 564700 293500
rect 564900 293300 565100 293500
rect 565300 293300 565500 293500
rect 565700 293300 565900 293500
rect 566100 293300 566300 293500
rect 566500 293300 566700 293500
rect 566900 293300 567100 293500
rect 567300 293300 567500 293500
rect 567700 293300 568000 293500
rect 562200 293200 568000 293300
rect 550109 292162 550129 292302
rect 550259 292162 550389 292302
rect 550519 292162 550539 292302
rect 550109 292152 550539 292162
rect 535989 292052 547499 292142
rect 530609 291972 531049 291992
rect 538359 291832 538589 291852
rect 538359 291752 538379 291832
rect 538459 291752 538489 291832
rect 538569 291752 538589 291832
rect 538359 291732 538589 291752
rect 540769 291832 540999 291842
rect 540769 291752 540789 291832
rect 540869 291752 540899 291832
rect 540979 291752 540999 291832
rect 540769 291732 540999 291752
rect 543229 291832 543459 291842
rect 543229 291752 543249 291832
rect 543329 291752 543359 291832
rect 543439 291752 543459 291832
rect 543229 291732 543459 291752
rect 534849 291652 535139 291672
rect 534849 291542 534869 291652
rect 534959 291542 535029 291652
rect 535119 291542 535139 291652
rect 534849 291532 535139 291542
rect 544779 291602 545071 291612
rect 544779 291522 544799 291602
rect 544879 291522 544969 291602
rect 545049 291522 545071 291602
rect 544779 291514 545071 291522
rect 547089 291322 547499 292052
rect 533839 291300 547499 291322
rect 533839 291200 547200 291300
rect 533839 291142 545900 291200
rect 546100 291142 546200 291200
rect 336600 290940 533500 291100
rect 533839 291062 536119 291142
rect 536209 291062 536299 291142
rect 536389 291062 538649 291142
rect 538739 291062 538809 291142
rect 538899 291062 541119 291142
rect 541209 291062 541279 291142
rect 541369 291062 543569 291142
rect 543659 291062 543729 291142
rect 543819 291062 545900 291142
rect 546159 291062 546200 291142
rect 533839 291000 545900 291062
rect 546100 291000 546200 291062
rect 546400 291000 546500 291200
rect 546700 291000 546800 291200
rect 547000 291100 547200 291200
rect 547400 291100 547499 291300
rect 547000 291000 547499 291100
rect 533839 290962 547200 291000
rect 336600 290880 533080 290940
rect 533140 290880 533180 290940
rect 533240 290880 533280 290940
rect 533340 290880 533500 290940
rect 336600 290820 533500 290880
rect 336600 290760 533080 290820
rect 533140 290760 533180 290820
rect 533240 290760 533280 290820
rect 533340 290760 533500 290820
rect 336600 290720 533500 290760
rect 336600 290660 533080 290720
rect 533140 290660 533180 290720
rect 533240 290660 533280 290720
rect 533340 290660 533500 290720
rect 336600 290580 533500 290660
rect 336600 290520 533080 290580
rect 533140 290520 533180 290580
rect 533240 290520 533280 290580
rect 533340 290520 533500 290580
rect 336600 290480 533500 290520
rect 336600 290420 533080 290480
rect 533140 290420 533180 290480
rect 533240 290420 533280 290480
rect 533340 290420 533500 290480
rect 336600 290380 533500 290420
rect 336600 290320 533080 290380
rect 533140 290320 533180 290380
rect 533240 290320 533280 290380
rect 533340 290320 533500 290380
rect 336600 290280 533500 290320
rect 336600 290220 533080 290280
rect 533140 290220 533180 290280
rect 533240 290220 533280 290280
rect 533340 290220 533500 290280
rect 336600 289800 533500 290220
rect 547089 290800 547200 290962
rect 547400 290800 547499 291000
rect 547089 290700 547499 290800
rect 547089 290500 547200 290700
rect 547400 290500 547499 290700
rect 547089 290400 547499 290500
rect 547089 290200 547200 290400
rect 547400 290200 547499 290400
rect 547089 290192 547499 290200
rect 534209 290100 547499 290192
rect 534209 290072 545800 290100
rect 534209 290062 536299 290072
rect 534209 289982 536119 290062
rect 536209 289992 536299 290062
rect 536389 290062 545800 290072
rect 536389 289992 538649 290062
rect 536209 289982 538649 289992
rect 538739 289982 538809 290062
rect 538899 289982 541119 290062
rect 541209 289982 541279 290062
rect 541369 289982 543569 290062
rect 543659 289982 543729 290062
rect 543819 289982 545800 290062
rect 534209 289900 545800 289982
rect 546000 290062 546100 290100
rect 546300 290062 546400 290100
rect 546000 289982 546069 290062
rect 546319 289982 546400 290062
rect 546000 289900 546100 289982
rect 546300 289900 546400 289982
rect 546600 289900 546800 290100
rect 547000 289900 547499 290100
rect 534209 289852 547499 289900
rect 336600 285700 511200 289800
rect 531739 289252 532089 289262
rect 531739 289122 531759 289252
rect 531849 289122 531969 289252
rect 532059 289122 532089 289252
rect 549059 289242 549319 289252
rect 549059 289152 549069 289242
rect 549139 289152 549229 289242
rect 549299 289152 549319 289242
rect 531739 288940 532089 289122
rect 538359 289132 538589 289142
rect 538359 289052 538379 289132
rect 538459 289052 538489 289132
rect 538569 289052 538589 289132
rect 538359 289042 538589 289052
rect 540769 289132 540999 289152
rect 540769 289052 540789 289132
rect 540869 289052 540899 289132
rect 540979 289052 540999 289132
rect 543229 289142 543459 289152
rect 543229 289062 543249 289142
rect 543329 289062 543359 289142
rect 543439 289062 543459 289142
rect 543229 289052 543459 289062
rect 540769 289042 540999 289052
rect 511500 288912 536560 288940
rect 549059 288912 549319 289152
rect 511500 288800 550449 288912
rect 511500 288600 511700 288800
rect 511900 288600 512100 288800
rect 512300 288600 512500 288800
rect 512700 288600 512900 288800
rect 513100 288600 513300 288800
rect 513500 288600 513700 288800
rect 513900 288600 514100 288800
rect 514300 288600 514500 288800
rect 514700 288600 514900 288800
rect 515100 288600 515300 288800
rect 515500 288600 515700 288800
rect 515900 288600 516100 288800
rect 516300 288600 516500 288800
rect 516700 288772 550449 288800
rect 516700 288662 538279 288772
rect 538389 288662 539139 288772
rect 539249 288662 540349 288772
rect 540459 288662 541199 288772
rect 541309 288662 542769 288772
rect 542879 288662 543649 288772
rect 543759 288662 550449 288772
rect 516700 288600 550449 288662
rect 511500 288552 550449 288600
rect 511500 288400 536560 288552
rect 545399 288542 550449 288552
rect 572600 288764 574700 288900
rect 572600 288704 572750 288764
rect 572810 288704 572890 288764
rect 572950 288704 573065 288764
rect 573125 288704 573255 288764
rect 573315 288704 573415 288764
rect 573475 288704 573605 288764
rect 573665 288704 573805 288764
rect 573865 288704 573985 288764
rect 574045 288704 574175 288764
rect 574235 288704 574375 288764
rect 574435 288754 574700 288764
rect 574435 288704 574540 288754
rect 572600 288700 574540 288704
rect 572600 288564 572800 288700
rect 573100 288564 573300 288700
rect 573600 288564 573800 288700
rect 574100 288564 574300 288700
rect 511500 288200 511700 288400
rect 511900 288200 512100 288400
rect 512300 288200 512500 288400
rect 512700 288200 512900 288400
rect 513100 288200 513300 288400
rect 513500 288200 513700 288400
rect 513900 288200 514100 288400
rect 514300 288200 514500 288400
rect 514700 288200 514900 288400
rect 515100 288200 515300 288400
rect 515500 288200 515700 288400
rect 515900 288200 516100 288400
rect 516300 288200 516500 288400
rect 516700 288200 536560 288400
rect 539559 288392 539829 288402
rect 537069 288372 537339 288392
rect 537069 288292 537089 288372
rect 537169 288292 537239 288372
rect 537319 288292 537339 288372
rect 539559 288312 539579 288392
rect 539659 288312 539729 288392
rect 539809 288312 539829 288392
rect 539559 288292 539829 288312
rect 542039 288392 542309 288402
rect 542039 288312 542059 288392
rect 542139 288312 542199 288392
rect 542279 288312 542309 288392
rect 542039 288292 542309 288312
rect 537069 288262 537339 288292
rect 511500 288000 536560 288200
rect 511500 287800 511700 288000
rect 511900 287800 512100 288000
rect 512300 287800 512500 288000
rect 512700 287800 512900 288000
rect 513100 287800 513300 288000
rect 513500 287800 513700 288000
rect 513900 287800 514100 288000
rect 514300 287800 514500 288000
rect 514700 287800 514900 288000
rect 515100 287800 515300 288000
rect 515500 287800 515700 288000
rect 515900 287800 516100 288000
rect 516300 287800 516500 288000
rect 516700 287852 536560 288000
rect 545469 287852 545689 288542
rect 516700 287800 545689 287852
rect 511500 287652 545689 287800
rect 511500 287600 537569 287652
rect 511500 287400 511700 287600
rect 511900 287400 512100 287600
rect 512300 287400 512500 287600
rect 512700 287400 512900 287600
rect 513100 287400 513300 287600
rect 513500 287400 513700 287600
rect 513900 287400 514100 287600
rect 514300 287400 514500 287600
rect 514700 287400 514900 287600
rect 515100 287400 515300 287600
rect 515500 287400 515700 287600
rect 515900 287400 516100 287600
rect 516300 287400 516500 287600
rect 516700 287562 537569 287600
rect 537679 287562 542479 287652
rect 542589 287562 545689 287652
rect 572600 288504 572750 288564
rect 573125 288504 573255 288564
rect 573600 288504 573605 288564
rect 573665 288504 573800 288564
rect 574100 288504 574175 288564
rect 574235 288504 574300 288564
rect 572600 288400 572800 288504
rect 573100 288400 573300 288504
rect 573600 288400 573800 288504
rect 574100 288400 574300 288504
rect 574600 288400 574700 288754
rect 572600 288364 574700 288400
rect 572600 288304 572750 288364
rect 572810 288304 572890 288364
rect 572950 288304 573065 288364
rect 573125 288304 573255 288364
rect 573315 288304 573415 288364
rect 573475 288304 573605 288364
rect 573665 288304 573805 288364
rect 573865 288304 573985 288364
rect 574045 288304 574175 288364
rect 574235 288304 574375 288364
rect 574435 288304 574540 288364
rect 574600 288304 574700 288364
rect 572600 288200 574700 288304
rect 572600 288174 572800 288200
rect 573100 288174 573300 288200
rect 573600 288174 573800 288200
rect 574100 288174 574300 288200
rect 572600 288114 572750 288174
rect 573125 288114 573255 288174
rect 573600 288114 573605 288174
rect 573665 288114 573800 288174
rect 574100 288114 574175 288174
rect 574235 288114 574300 288174
rect 572600 287974 572800 288114
rect 573100 287974 573300 288114
rect 573600 287974 573800 288114
rect 574100 287974 574300 288114
rect 572600 287914 572750 287974
rect 573125 287914 573255 287974
rect 573600 287914 573605 287974
rect 573665 287914 573800 287974
rect 574100 287914 574175 287974
rect 574235 287914 574300 287974
rect 572600 287900 572800 287914
rect 573100 287900 573300 287914
rect 573600 287900 573800 287914
rect 574100 287900 574300 287914
rect 574600 287900 574700 288200
rect 572600 287774 574700 287900
rect 572600 287714 572750 287774
rect 572810 287714 572890 287774
rect 572950 287714 573065 287774
rect 573125 287714 573255 287774
rect 573315 287714 573415 287774
rect 573475 287714 573605 287774
rect 573665 287714 573805 287774
rect 573865 287714 573985 287774
rect 574045 287714 574175 287774
rect 574235 287714 574375 287774
rect 574435 287714 574540 287774
rect 574600 287714 574700 287774
rect 572600 287600 574700 287714
rect 578320 288600 578660 288660
rect 578320 288520 578360 288600
rect 578440 288520 578540 288600
rect 578620 288520 578660 288600
rect 578320 288440 578660 288520
rect 578320 288360 578360 288440
rect 578440 288360 578540 288440
rect 578620 288360 578660 288440
rect 578320 288280 578660 288360
rect 578320 288200 578360 288280
rect 578440 288200 578540 288280
rect 578620 288200 578660 288280
rect 578320 288100 578660 288200
rect 578320 288020 578360 288100
rect 578440 288020 578540 288100
rect 578620 288020 578660 288100
rect 578320 287940 578660 288020
rect 578320 287860 578360 287940
rect 578440 287860 578540 287940
rect 578620 287860 578660 287940
rect 516700 287400 545689 287562
rect 511500 287392 545689 287400
rect 511500 287200 536560 287392
rect 511500 287000 511700 287200
rect 511900 287000 512100 287200
rect 512300 287000 512500 287200
rect 512700 287000 512900 287200
rect 513100 287000 513300 287200
rect 513500 287000 513700 287200
rect 513900 287000 514100 287200
rect 514300 287000 514500 287200
rect 514700 287000 514900 287200
rect 515100 287000 515300 287200
rect 515500 287000 515700 287200
rect 515900 287000 516100 287200
rect 516300 287000 516500 287200
rect 516700 287000 536560 287200
rect 511500 286800 536560 287000
rect 511500 286600 511700 286800
rect 511900 286600 512100 286800
rect 512300 286600 512500 286800
rect 512700 286600 512900 286800
rect 513100 286600 513300 286800
rect 513500 286600 513700 286800
rect 513900 286600 514100 286800
rect 514300 286600 514500 286800
rect 514700 286600 514900 286800
rect 515100 286600 515300 286800
rect 515500 286600 515700 286800
rect 515900 286600 516100 286800
rect 516300 286600 516500 286800
rect 516700 286672 536560 286800
rect 545469 286672 545689 287392
rect 578320 287200 578660 287860
rect 516700 286600 545689 286672
rect 511500 286460 545689 286600
rect 511500 286400 511600 286460
rect 535629 286452 545689 286460
rect 535629 286352 537509 286452
rect 537629 286352 538729 286452
rect 538849 286352 539939 286452
rect 540059 286352 541159 286452
rect 541279 286442 543599 286452
rect 541279 286352 542389 286442
rect 535629 286342 542389 286352
rect 542509 286352 543599 286442
rect 543719 286352 545689 286452
rect 542509 286342 545689 286352
rect 535629 286212 545689 286342
rect 557600 286200 582600 287200
rect 557600 286000 557700 286200
rect 557900 286000 558100 286200
rect 558300 286000 558500 286200
rect 558700 286000 558900 286200
rect 559100 286000 559300 286200
rect 559500 286000 582600 286200
rect 537344 285500 543804 285938
rect 557600 285800 582600 286000
rect 557600 285600 557700 285800
rect 557900 285600 558100 285800
rect 558300 285600 558500 285800
rect 558700 285600 558900 285800
rect 559100 285600 559300 285800
rect 559500 285600 582600 285800
rect 537344 285478 549100 285500
rect 537344 285318 537384 285478
rect 537544 285318 538444 285478
rect 538604 285318 539904 285478
rect 540064 285318 541124 285478
rect 541284 285318 542604 285478
rect 542764 285318 543604 285478
rect 543764 285400 549100 285478
rect 543764 285318 545800 285400
rect 537344 285200 545800 285318
rect 546000 285200 546200 285400
rect 546400 285200 546600 285400
rect 546800 285200 547000 285400
rect 547200 285200 547400 285400
rect 547600 285200 547800 285400
rect 548000 285200 548200 285400
rect 548400 285200 548600 285400
rect 548800 285200 549100 285400
rect 537344 285000 549100 285200
rect 537344 284898 545800 285000
rect 537344 284738 537384 284898
rect 537544 284738 538444 284898
rect 538604 284738 539904 284898
rect 540064 284738 541124 284898
rect 541284 284738 542604 284898
rect 542764 284738 543604 284898
rect 543764 284800 545800 284898
rect 546000 284800 546200 285000
rect 546400 284800 546600 285000
rect 546800 284800 547000 285000
rect 547200 284800 547400 285000
rect 547600 284800 547800 285000
rect 548000 284800 548200 285000
rect 548400 284800 548600 285000
rect 548800 284800 549100 285000
rect 543764 284738 549100 284800
rect 537344 284718 549100 284738
rect 543600 284700 549100 284718
rect 557600 285400 582600 285600
rect 557600 285200 557700 285400
rect 557900 285200 558100 285400
rect 558300 285200 558500 285400
rect 558700 285200 558900 285400
rect 559100 285200 559300 285400
rect 559500 285200 582600 285400
rect 557600 285000 582600 285200
rect 557600 284800 557700 285000
rect 557900 284800 558100 285000
rect 558300 284800 558500 285000
rect 558700 284800 558900 285000
rect 559100 284800 559300 285000
rect 559500 284800 582600 285000
rect 557600 284600 582600 284800
rect 330400 284420 540780 284500
rect 330400 284360 540440 284420
rect 540500 284360 540540 284420
rect 540600 284360 540640 284420
rect 540700 284360 540780 284420
rect 330400 284320 540780 284360
rect 330400 284260 540440 284320
rect 540500 284260 540540 284320
rect 540600 284260 540640 284320
rect 540700 284260 540780 284320
rect 330400 284220 540780 284260
rect 330400 284160 540440 284220
rect 540500 284160 540540 284220
rect 540600 284160 540640 284220
rect 540700 284160 540780 284220
rect 330400 284120 540780 284160
rect 330400 284060 540440 284120
rect 540500 284060 540540 284120
rect 540600 284060 540640 284120
rect 540700 284060 540780 284120
rect 330400 284020 540780 284060
rect 557600 284400 557700 284600
rect 557900 284400 558100 284600
rect 558300 284400 558500 284600
rect 558700 284400 558900 284600
rect 559100 284400 559300 284600
rect 559500 284400 582600 284600
rect 557600 284200 582600 284400
rect 330400 279300 511000 284020
rect 557600 284000 557700 284200
rect 557900 284000 558100 284200
rect 558300 284000 558500 284200
rect 558700 284000 558900 284200
rect 559100 284000 559300 284200
rect 559500 284000 582600 284200
rect 557600 283800 582600 284000
rect 557600 283600 557700 283800
rect 557900 283600 558100 283800
rect 558300 283600 558500 283800
rect 558700 283600 558900 283800
rect 559100 283600 559300 283800
rect 559500 283600 582600 283800
rect 511500 283558 537760 283560
rect 511500 283518 543914 283558
rect 511500 283368 539764 283518
rect 539984 283368 540284 283518
rect 540504 283368 540704 283518
rect 540924 283368 541254 283518
rect 541474 283368 543914 283518
rect 511500 283200 543914 283368
rect 511500 283000 511900 283200
rect 512100 283000 512300 283200
rect 512500 283000 512700 283200
rect 512900 283000 513100 283200
rect 513300 283000 513500 283200
rect 513700 283000 513900 283200
rect 514100 283000 514300 283200
rect 514500 283000 514700 283200
rect 514900 283000 515100 283200
rect 515300 283000 515500 283200
rect 515700 283000 515900 283200
rect 516100 283000 516300 283200
rect 516500 283000 516700 283200
rect 516900 283000 543914 283200
rect 511500 282968 543914 283000
rect 511500 282958 539524 282968
rect 511500 282828 537404 282958
rect 537584 282828 538544 282958
rect 538724 282838 539524 282958
rect 539704 282838 540294 282968
rect 540474 282838 540734 282968
rect 540914 282958 542524 282968
rect 540914 282838 541454 282958
rect 538724 282828 541454 282838
rect 541634 282838 542524 282958
rect 542704 282838 543524 282968
rect 543704 282838 543914 282968
rect 541634 282828 543914 282838
rect 511500 282800 543914 282828
rect 511500 282600 511900 282800
rect 512100 282600 512300 282800
rect 512500 282600 512700 282800
rect 512900 282600 513100 282800
rect 513300 282600 513500 282800
rect 513700 282600 513900 282800
rect 514100 282600 514300 282800
rect 514500 282600 514700 282800
rect 514900 282600 515100 282800
rect 515300 282600 515500 282800
rect 515700 282600 515900 282800
rect 516100 282600 516300 282800
rect 516500 282600 516700 282800
rect 516900 282798 543914 282800
rect 516900 282600 537760 282798
rect 511500 282400 537760 282600
rect 511500 282200 511900 282400
rect 512100 282200 512300 282400
rect 512500 282200 512700 282400
rect 512900 282200 513100 282400
rect 513300 282200 513500 282400
rect 513700 282200 513900 282400
rect 514100 282200 514300 282400
rect 514500 282200 514700 282400
rect 514900 282200 515100 282400
rect 515300 282200 515500 282400
rect 515700 282200 515900 282400
rect 516100 282200 516300 282400
rect 516500 282200 516700 282400
rect 516900 282200 537760 282400
rect 511500 282000 537760 282200
rect 511500 281800 511900 282000
rect 512100 281800 512300 282000
rect 512500 281800 512700 282000
rect 512900 281800 513100 282000
rect 513300 281800 513500 282000
rect 513700 281800 513900 282000
rect 514100 281800 514300 282000
rect 514500 281800 514700 282000
rect 514900 281800 515100 282000
rect 515300 281800 515500 282000
rect 515700 281800 515900 282000
rect 516100 281800 516300 282000
rect 516500 281800 516700 282000
rect 516900 281800 537760 282000
rect 511500 281600 537760 281800
rect 511500 281400 511900 281600
rect 512100 281400 512300 281600
rect 512500 281400 512700 281600
rect 512900 281400 513100 281600
rect 513300 281400 513500 281600
rect 513700 281400 513900 281600
rect 514100 281400 514300 281600
rect 514500 281400 514700 281600
rect 514900 281400 515100 281600
rect 515300 281400 515500 281600
rect 515700 281400 515900 281600
rect 516100 281400 516300 281600
rect 516500 281400 516700 281600
rect 516900 281400 537760 281600
rect 511500 281200 537760 281400
rect 511500 281000 511900 281200
rect 512100 281000 512300 281200
rect 512500 281000 512700 281200
rect 512900 281000 513100 281200
rect 513300 281000 513500 281200
rect 513700 281000 513900 281200
rect 514100 281000 514300 281200
rect 514500 281000 514700 281200
rect 514900 281000 515100 281200
rect 515300 281000 515500 281200
rect 515700 281000 515900 281200
rect 516100 281000 516300 281200
rect 516500 281000 516700 281200
rect 516900 281058 537760 281200
rect 516900 281000 537364 281058
rect 511500 280938 537364 281000
rect 537484 280938 537760 281058
rect 511500 280800 537760 280938
rect 511500 280600 511900 280800
rect 512100 280600 512300 280800
rect 512500 280600 512700 280800
rect 512900 280600 513100 280800
rect 513300 280600 513500 280800
rect 513700 280600 513900 280800
rect 514100 280600 514300 280800
rect 514500 280600 514700 280800
rect 514900 280600 515100 280800
rect 515300 280600 515500 280800
rect 515700 280600 515900 280800
rect 516100 280600 516300 280800
rect 516500 280600 516700 280800
rect 516900 280600 537760 280800
rect 511500 280460 537760 280600
rect 543594 281400 543914 282798
rect 557600 283400 582600 283600
rect 557600 283200 557700 283400
rect 557900 283200 558100 283400
rect 558300 283200 558500 283400
rect 558700 283200 558900 283400
rect 559100 283200 559300 283400
rect 559500 283200 582600 283400
rect 557600 283000 582600 283200
rect 557600 282800 557700 283000
rect 557900 282800 558100 283000
rect 558300 282800 558500 283000
rect 558700 282800 558900 283000
rect 559100 282800 559300 283000
rect 559500 282800 582600 283000
rect 557600 282600 582600 282800
rect 557600 282400 557700 282600
rect 557900 282400 558100 282600
rect 558300 282400 558500 282600
rect 558700 282400 558900 282600
rect 559100 282400 559300 282600
rect 559500 282400 582600 282600
rect 557600 281800 582600 282400
rect 543594 281300 568280 281400
rect 543594 281100 567900 281300
rect 568100 281100 568280 281300
rect 543594 281058 568280 281100
rect 543594 280938 543734 281058
rect 543854 281000 568280 281058
rect 543854 280938 567900 281000
rect 543594 280800 567900 280938
rect 568100 280800 568280 281000
rect 543594 280700 568280 280800
rect 543594 280500 567900 280700
rect 568100 280500 568280 280700
rect 537294 278058 537614 280460
rect 537294 277938 537364 278058
rect 537484 277938 537614 278058
rect 537294 275058 537614 277938
rect 537294 274938 537364 275058
rect 537484 274938 537614 275058
rect 537294 272058 537614 274938
rect 537294 271938 537364 272058
rect 537484 271938 537614 272058
rect 537294 269058 537614 271938
rect 537294 268938 537364 269058
rect 537484 268938 537614 269058
rect 537294 267758 537614 268938
rect 543594 280400 568280 280500
rect 543594 280200 567900 280400
rect 568100 280200 568280 280400
rect 543594 280100 568280 280200
rect 572700 281284 574700 281800
rect 572700 281224 572770 281284
rect 572830 281224 572910 281284
rect 572970 281224 573085 281284
rect 573145 281224 573275 281284
rect 573335 281224 573435 281284
rect 573495 281224 573625 281284
rect 573685 281224 573825 281284
rect 573885 281224 574005 281284
rect 574065 281224 574195 281284
rect 574255 281224 574395 281284
rect 574455 281274 574700 281284
rect 574455 281224 574560 281274
rect 572700 281214 574560 281224
rect 574620 281214 574700 281274
rect 572700 281084 574700 281214
rect 572700 281024 572770 281084
rect 572830 281024 572910 281084
rect 572970 281024 573085 281084
rect 573145 281024 573275 281084
rect 573335 281024 573435 281084
rect 573495 281024 573625 281084
rect 573685 281024 573825 281084
rect 573885 281024 574005 281084
rect 574065 281024 574195 281084
rect 574255 281024 574395 281084
rect 574455 281024 574560 281084
rect 574620 281024 574700 281084
rect 572700 280884 574700 281024
rect 572700 280824 572770 280884
rect 572830 280824 572910 280884
rect 572970 280824 573085 280884
rect 573145 280824 573275 280884
rect 573335 280824 573435 280884
rect 573495 280824 573625 280884
rect 573685 280824 573825 280884
rect 573885 280824 574005 280884
rect 574065 280824 574195 280884
rect 574255 280824 574395 280884
rect 574455 280824 574560 280884
rect 574620 280824 574700 280884
rect 572700 280694 574700 280824
rect 572700 280634 572770 280694
rect 572830 280634 572910 280694
rect 572970 280634 573085 280694
rect 573145 280634 573275 280694
rect 573335 280634 573435 280694
rect 573495 280634 573625 280694
rect 573685 280634 573825 280694
rect 573885 280634 574005 280694
rect 574065 280634 574195 280694
rect 574255 280634 574395 280694
rect 574455 280634 574560 280694
rect 574620 280634 574700 280694
rect 572700 280494 574700 280634
rect 572700 280434 572770 280494
rect 572830 280434 572910 280494
rect 572970 280434 573085 280494
rect 573145 280434 573275 280494
rect 573335 280434 573435 280494
rect 573495 280434 573625 280494
rect 573685 280434 573825 280494
rect 573885 280434 574005 280494
rect 574065 280434 574195 280494
rect 574255 280434 574395 280494
rect 574455 280434 574560 280494
rect 574620 280434 574700 280494
rect 572700 280294 574700 280434
rect 572700 280234 572770 280294
rect 572830 280234 572910 280294
rect 572970 280234 573085 280294
rect 573145 280234 573275 280294
rect 573335 280234 573435 280294
rect 573495 280234 573625 280294
rect 573685 280234 573825 280294
rect 573885 280234 574005 280294
rect 574065 280234 574195 280294
rect 574255 280234 574395 280294
rect 574455 280234 574560 280294
rect 574620 280234 574700 280294
rect 572700 280100 574700 280234
rect 543594 278058 543914 280100
rect 543594 277938 543734 278058
rect 543854 277938 543914 278058
rect 543594 275058 543914 277938
rect 543594 274938 543734 275058
rect 543854 274938 543914 275058
rect 543594 272058 543914 274938
rect 543594 271938 543734 272058
rect 543854 271938 543914 272058
rect 543594 269058 543914 271938
rect 543594 268938 543734 269058
rect 543854 268938 543914 269058
rect 543594 267758 543914 268938
rect 537294 267738 543914 267758
rect 537294 267728 542294 267738
rect 537294 267318 537744 267728
rect 538914 267318 539254 267728
rect 540424 267318 540774 267728
rect 541944 267328 542294 267728
rect 543464 267328 543914 267738
rect 541944 267318 543914 267328
rect 537294 267278 543914 267318
rect 580200 269600 582600 281800
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 580200 269342 584000 269600
rect 580200 269230 584800 269342
rect 580200 267200 584000 269230
rect 545600 248600 584000 248800
rect 545600 248400 546000 248600
rect 546200 248400 546400 248600
rect 546600 248400 546800 248600
rect 547000 248400 547200 248600
rect 547400 248400 547600 248600
rect 547800 248400 548000 248600
rect 548200 248400 548400 248600
rect 548600 248400 548800 248600
rect 549000 248400 584000 248600
rect 545600 248200 584000 248400
rect 545600 248000 546000 248200
rect 546200 248000 546400 248200
rect 546600 248000 546800 248200
rect 547000 248000 547200 248200
rect 547400 248000 547600 248200
rect 547800 248000 548000 248200
rect 548200 248000 548400 248200
rect 548600 248000 548800 248200
rect 549000 248000 584000 248200
rect 545600 247800 584000 248000
rect 545600 247600 546000 247800
rect 546200 247600 546400 247800
rect 546600 247600 546800 247800
rect 547000 247600 547200 247800
rect 547400 247600 547600 247800
rect 547800 247600 548000 247800
rect 548200 247600 548400 247800
rect 548600 247600 548800 247800
rect 549000 247600 584000 247800
rect 545600 247400 584000 247600
rect 545600 247200 546000 247400
rect 546200 247200 546400 247400
rect 546600 247200 546800 247400
rect 547000 247200 547200 247400
rect 547400 247200 547600 247400
rect 547800 247200 548000 247400
rect 548200 247200 548400 247400
rect 548600 247200 548800 247400
rect 549000 247200 584000 247400
rect 545600 247000 584000 247200
rect 545600 246800 546000 247000
rect 546200 246800 546400 247000
rect 546600 246800 546800 247000
rect 547000 246800 547200 247000
rect 547400 246800 547600 247000
rect 547800 246800 548000 247000
rect 548200 246800 548400 247000
rect 548600 246800 548800 247000
rect 549000 246800 584000 247000
rect 545600 246600 584000 246800
rect 545600 246400 546000 246600
rect 546200 246400 546400 246600
rect 546600 246400 546800 246600
rect 547000 246400 547200 246600
rect 547400 246400 547600 246600
rect 547800 246400 548000 246600
rect 548200 246400 548400 246600
rect 548600 246400 548800 246600
rect 549000 246400 584000 246600
rect 545600 246200 584000 246400
rect 545600 246000 546000 246200
rect 546200 246000 546400 246200
rect 546600 246000 546800 246200
rect 547000 246000 547200 246200
rect 547400 246000 547600 246200
rect 547800 246000 548000 246200
rect 548200 246000 548400 246200
rect 548600 246000 548800 246200
rect 549000 246000 584000 246200
rect 545600 245800 584000 246000
rect 545600 245600 546000 245800
rect 546200 245600 546400 245800
rect 546600 245600 546800 245800
rect 547000 245600 547200 245800
rect 547400 245600 547600 245800
rect 547800 245600 548000 245800
rect 548200 245600 548400 245800
rect 548600 245600 548800 245800
rect 549000 245600 584000 245800
rect 545600 245400 584000 245600
rect 545600 245200 546000 245400
rect 546200 245200 546400 245400
rect 546600 245200 546800 245400
rect 547000 245200 547200 245400
rect 547400 245200 547600 245400
rect 547800 245200 548000 245400
rect 548200 245200 548400 245400
rect 548600 245200 548800 245400
rect 549000 245200 584000 245400
rect 545600 245000 584000 245200
rect 545600 244800 546000 245000
rect 546200 244800 546400 245000
rect 546600 244800 546800 245000
rect 547000 244800 547200 245000
rect 547400 244800 547600 245000
rect 547800 244800 548000 245000
rect 548200 244800 548400 245000
rect 548600 244800 548800 245000
rect 549000 244800 584000 245000
rect 545600 244600 584000 244800
rect 545600 244400 546000 244600
rect 546200 244400 546400 244600
rect 546600 244400 546800 244600
rect 547000 244400 547200 244600
rect 547400 244400 547600 244600
rect 547800 244400 548000 244600
rect 548200 244400 548400 244600
rect 548600 244400 548800 244600
rect 549000 244400 584000 244600
rect 545600 244200 584000 244400
rect 545600 244000 546000 244200
rect 546200 244000 546400 244200
rect 546600 244000 546800 244200
rect 547000 244000 547200 244200
rect 547400 244000 547600 244200
rect 547800 244000 548000 244200
rect 548200 244000 548400 244200
rect 548600 244000 548800 244200
rect 549000 244000 584000 244200
rect 545600 243800 584000 244000
rect 545600 243600 546000 243800
rect 546200 243600 546400 243800
rect 546600 243600 546800 243800
rect 547000 243600 547200 243800
rect 547400 243600 547600 243800
rect 547800 243600 548000 243800
rect 548200 243600 548400 243800
rect 548600 243600 548800 243800
rect 549000 243600 584000 243800
rect 545600 243400 584000 243600
rect 545600 243200 546000 243400
rect 546200 243200 546400 243400
rect 546600 243200 546800 243400
rect 547000 243200 547200 243400
rect 547400 243200 547600 243400
rect 547800 243200 548000 243400
rect 548200 243200 548400 243400
rect 548600 243200 548800 243400
rect 549000 243200 584000 243400
rect 545600 243000 584000 243200
rect 545600 242800 546000 243000
rect 546200 242800 546400 243000
rect 546600 242800 546800 243000
rect 547000 242800 547200 243000
rect 547400 242800 547600 243000
rect 547800 242800 548000 243000
rect 548200 242800 548400 243000
rect 548600 242800 548800 243000
rect 549000 242800 584000 243000
rect 545600 242600 584000 242800
rect 545600 242400 546000 242600
rect 546200 242400 546400 242600
rect 546600 242400 546800 242600
rect 547000 242400 547200 242600
rect 547400 242400 547600 242600
rect 547800 242400 548000 242600
rect 548200 242400 548400 242600
rect 548600 242400 548800 242600
rect 549000 242400 584000 242600
rect 545600 242200 584000 242400
rect 545600 242000 546000 242200
rect 546200 242000 546400 242200
rect 546600 242000 546800 242200
rect 547000 242000 547200 242200
rect 547400 242000 547600 242200
rect 547800 242000 548000 242200
rect 548200 242000 548400 242200
rect 548600 242000 548800 242200
rect 549000 242000 584000 242200
rect 545600 241800 584000 242000
rect 545600 241600 546000 241800
rect 546200 241600 546400 241800
rect 546600 241600 546800 241800
rect 547000 241600 547200 241800
rect 547400 241600 547600 241800
rect 547800 241600 548000 241800
rect 548200 241600 548400 241800
rect 548600 241600 548800 241800
rect 549000 241600 584000 241800
rect 545600 241400 584000 241600
rect 545600 241200 546000 241400
rect 546200 241200 546400 241400
rect 546600 241200 546800 241400
rect 547000 241200 547200 241400
rect 547400 241200 547600 241400
rect 547800 241200 548000 241400
rect 548200 241200 548400 241400
rect 548600 241200 548800 241400
rect 549000 241200 584000 241400
rect 545600 241000 584000 241200
rect 545600 240800 546000 241000
rect 546200 240800 546400 241000
rect 546600 240800 546800 241000
rect 547000 240800 547200 241000
rect 547400 240800 547600 241000
rect 547800 240800 548000 241000
rect 548200 240800 548400 241000
rect 548600 240800 548800 241000
rect 549000 240800 584000 241000
rect 545600 240600 584000 240800
rect 545600 240400 546000 240600
rect 546200 240400 546400 240600
rect 546600 240400 546800 240600
rect 547000 240400 547200 240600
rect 547400 240400 547600 240600
rect 547800 240400 548000 240600
rect 548200 240400 548400 240600
rect 548600 240400 548800 240600
rect 549000 240400 584000 240600
rect 545600 240200 584000 240400
rect 545600 240000 546000 240200
rect 546200 240000 546400 240200
rect 546600 240000 546800 240200
rect 547000 240000 547200 240200
rect 547400 240000 547600 240200
rect 547800 240000 548000 240200
rect 548200 240000 548400 240200
rect 548600 240000 548800 240200
rect 549000 240030 584000 240200
rect 549000 240000 584800 240030
rect 545600 239800 584800 240000
rect 545600 239600 546000 239800
rect 546200 239600 546400 239800
rect 546600 239600 546800 239800
rect 547000 239600 547200 239800
rect 547400 239600 547600 239800
rect 547800 239600 548000 239800
rect 548200 239600 548400 239800
rect 548600 239600 548800 239800
rect 549000 239600 584800 239800
rect 545600 239400 584800 239600
rect 545600 239200 546000 239400
rect 546200 239200 546400 239400
rect 546600 239200 546800 239400
rect 547000 239200 547200 239400
rect 547400 239200 547600 239400
rect 547800 239200 548000 239400
rect 548200 239200 548400 239400
rect 548600 239200 548800 239400
rect 549000 239200 584800 239400
rect 545600 239000 584800 239200
rect 545600 238800 546000 239000
rect 546200 238800 546400 239000
rect 546600 238800 546800 239000
rect 547000 238800 547200 239000
rect 547400 238800 547600 239000
rect 547800 238800 548000 239000
rect 548200 238800 548400 239000
rect 548600 238800 548800 239000
rect 549000 238800 584800 239000
rect 545600 238600 584800 238800
rect 545600 238400 546000 238600
rect 546200 238400 546400 238600
rect 546600 238400 546800 238600
rect 547000 238400 547200 238600
rect 547400 238400 547600 238600
rect 547800 238400 548000 238600
rect 548200 238400 548400 238600
rect 548600 238400 548800 238600
rect 549000 238400 584800 238600
rect 545600 238200 584800 238400
rect 545600 238000 546000 238200
rect 546200 238000 546400 238200
rect 546600 238000 546800 238200
rect 547000 238000 547200 238200
rect 547400 238000 547600 238200
rect 547800 238000 548000 238200
rect 548200 238000 548400 238200
rect 548600 238000 548800 238200
rect 549000 238000 584800 238200
rect 545600 237800 584800 238000
rect 545600 237600 546000 237800
rect 546200 237600 546400 237800
rect 546600 237600 546800 237800
rect 547000 237600 547200 237800
rect 547400 237600 547600 237800
rect 547800 237600 548000 237800
rect 548200 237600 548400 237800
rect 548600 237600 548800 237800
rect 549000 237600 584800 237800
rect 545600 237400 584800 237600
rect 545600 237200 546000 237400
rect 546200 237200 546400 237400
rect 546600 237200 546800 237400
rect 547000 237200 547200 237400
rect 547400 237200 547600 237400
rect 547800 237200 548000 237400
rect 548200 237200 548400 237400
rect 548600 237200 548800 237400
rect 549000 237200 584800 237400
rect 545600 237000 584800 237200
rect 545600 236800 546000 237000
rect 546200 236800 546400 237000
rect 546600 236800 546800 237000
rect 547000 236800 547200 237000
rect 547400 236800 547600 237000
rect 547800 236800 548000 237000
rect 548200 236800 548400 237000
rect 548600 236800 548800 237000
rect 549000 236800 584800 237000
rect 545600 236600 584800 236800
rect 545600 236400 546000 236600
rect 546200 236400 546400 236600
rect 546600 236400 546800 236600
rect 547000 236400 547200 236600
rect 547400 236400 547600 236600
rect 547800 236400 548000 236600
rect 548200 236400 548400 236600
rect 548600 236400 548800 236600
rect 549000 236400 584800 236600
rect 545600 236200 584800 236400
rect 545600 236000 546000 236200
rect 546200 236000 546400 236200
rect 546600 236000 546800 236200
rect 547000 236000 547200 236200
rect 547400 236000 547600 236200
rect 547800 236000 548000 236200
rect 548200 236000 548400 236200
rect 548600 236000 548800 236200
rect 549000 236000 584800 236200
rect 545600 235800 584800 236000
rect 545600 235600 546000 235800
rect 546200 235600 546400 235800
rect 546600 235600 546800 235800
rect 547000 235600 547200 235800
rect 547400 235600 547600 235800
rect 547800 235600 548000 235800
rect 548200 235600 548400 235800
rect 548600 235600 548800 235800
rect 549000 235600 584800 235800
rect 545600 235400 584800 235600
rect 545600 235200 546000 235400
rect 546200 235200 546400 235400
rect 546600 235200 546800 235400
rect 547000 235200 547200 235400
rect 547400 235200 547600 235400
rect 547800 235200 548000 235400
rect 548200 235200 548400 235400
rect 548600 235200 548800 235400
rect 549000 235230 584800 235400
rect 549000 235200 584000 235230
rect 545600 235000 584000 235200
rect 545600 234800 546000 235000
rect 546200 234800 546400 235000
rect 546600 234800 546800 235000
rect 547000 234800 547200 235000
rect 547400 234800 547600 235000
rect 547800 234800 548000 235000
rect 548200 234800 548400 235000
rect 548600 234800 548800 235000
rect 549000 234800 584000 235000
rect 545600 234700 584000 234800
rect 545600 234500 546000 234700
rect 546200 234500 546400 234700
rect 546600 234500 546800 234700
rect 547000 234500 547200 234700
rect 547400 234500 547600 234700
rect 547800 234500 548000 234700
rect 548200 234500 548400 234700
rect 548600 234500 548800 234700
rect 549000 234500 584000 234700
rect 545600 234400 584000 234500
rect 545600 234200 546000 234400
rect 546200 234200 546400 234400
rect 546600 234200 546800 234400
rect 547000 234200 547200 234400
rect 547400 234200 547600 234400
rect 547800 234200 548000 234400
rect 548200 234200 548400 234400
rect 548600 234200 548800 234400
rect 549000 234200 584000 234400
rect 545600 234000 584000 234200
rect 545600 233800 546000 234000
rect 546200 233800 546400 234000
rect 546600 233800 546800 234000
rect 547000 233800 547200 234000
rect 547400 233800 547600 234000
rect 547800 233800 548000 234000
rect 548200 233800 548400 234000
rect 548600 233800 548800 234000
rect 549000 233800 584000 234000
rect 545600 233400 584000 233800
rect 574600 230030 584000 233400
rect 574600 225230 584800 230030
rect 574600 225100 584000 225230
rect 511500 195600 572000 196500
rect 511500 195200 512000 195600
rect 512400 195200 512800 195600
rect 513200 195200 513600 195600
rect 514000 195200 514400 195600
rect 514800 195200 515200 195600
rect 515600 195200 516000 195600
rect 516400 195200 572000 195600
rect 511500 194800 572000 195200
rect 511500 194400 512000 194800
rect 512400 194400 512800 194800
rect 513200 194400 513600 194800
rect 514000 194400 514400 194800
rect 514800 194400 515200 194800
rect 515600 194400 516000 194800
rect 516400 194400 572000 194800
rect 511500 194000 572000 194400
rect 511500 193600 512000 194000
rect 512400 193600 512800 194000
rect 513200 193600 513600 194000
rect 514000 193600 514400 194000
rect 514800 193600 515200 194000
rect 515600 193600 516000 194000
rect 516400 193600 572000 194000
rect 511500 193200 572000 193600
rect 511500 192800 512000 193200
rect 512400 192800 512800 193200
rect 513200 192800 513600 193200
rect 514000 192800 514400 193200
rect 514800 192800 515200 193200
rect 515600 192800 516000 193200
rect 516400 192800 572000 193200
rect 511500 192400 572000 192800
rect 511500 192000 512000 192400
rect 512400 192000 512800 192400
rect 513200 192000 513600 192400
rect 514000 192000 514400 192400
rect 514800 192000 515200 192400
rect 515600 192000 516000 192400
rect 516400 192000 572000 192400
rect 511500 191600 572000 192000
rect 511500 191200 512000 191600
rect 512400 191200 512800 191600
rect 513200 191200 513600 191600
rect 514000 191200 514400 191600
rect 514800 191200 515200 191600
rect 515600 191200 516000 191600
rect 516400 191200 572000 191600
rect 511500 190800 572000 191200
rect 511500 190400 512000 190800
rect 512400 190400 512800 190800
rect 513200 190400 513600 190800
rect 514000 190400 514400 190800
rect 514800 190400 515200 190800
rect 515600 190400 516000 190800
rect 516400 190400 572000 190800
rect 511500 190000 572000 190400
rect 511500 189600 512000 190000
rect 512400 189600 512800 190000
rect 513200 189600 513600 190000
rect 514000 189600 514400 190000
rect 514800 189600 515200 190000
rect 515600 189600 516000 190000
rect 516400 189600 572000 190000
rect 511500 189200 572000 189600
rect 511500 188800 512000 189200
rect 512400 188800 512800 189200
rect 513200 188800 513600 189200
rect 514000 188800 514400 189200
rect 514800 188800 515200 189200
rect 515600 188800 516000 189200
rect 516400 188800 572000 189200
rect 511500 188400 572000 188800
rect 511500 188000 512000 188400
rect 512400 188000 512800 188400
rect 513200 188000 513600 188400
rect 514000 188000 514400 188400
rect 514800 188000 515200 188400
rect 515600 188000 516000 188400
rect 516400 188000 572000 188400
rect 511500 187600 572000 188000
rect 511500 187200 512000 187600
rect 512400 187200 512800 187600
rect 513200 187200 513600 187600
rect 514000 187200 514400 187600
rect 514800 187200 515200 187600
rect 515600 187200 516000 187600
rect 516400 187200 572000 187600
rect 511500 186800 572000 187200
rect 511500 186400 512000 186800
rect 512400 186400 512800 186800
rect 513200 186400 513600 186800
rect 514000 186400 514400 186800
rect 514800 186400 515200 186800
rect 515600 186400 516000 186800
rect 516400 186400 572000 186800
rect 511500 186000 572000 186400
rect 511500 185600 512000 186000
rect 512400 185600 512800 186000
rect 513200 185600 513600 186000
rect 514000 185600 514400 186000
rect 514800 185600 515200 186000
rect 515600 185600 516000 186000
rect 516400 185600 572000 186000
rect 511500 185200 572000 185600
rect 511500 184800 512000 185200
rect 512400 184800 512800 185200
rect 513200 184800 513600 185200
rect 514000 184800 514400 185200
rect 514800 184800 515200 185200
rect 515600 184800 516000 185200
rect 516400 184800 572000 185200
rect 511500 184400 572000 184800
rect 511500 184000 512000 184400
rect 512400 184000 512800 184400
rect 513200 184000 513600 184400
rect 514000 184000 514400 184400
rect 514800 184000 515200 184400
rect 515600 184000 516000 184400
rect 516400 184000 572000 184400
rect 511500 183600 572000 184000
rect 511500 183200 512000 183600
rect 512400 183200 512800 183600
rect 513200 183200 513600 183600
rect 514000 183200 514400 183600
rect 514800 183200 515200 183600
rect 515600 183200 516000 183600
rect 516400 183200 572000 183600
rect 511500 182800 572000 183200
rect 511500 182400 512000 182800
rect 512400 182400 512800 182800
rect 513200 182400 513600 182800
rect 514000 182400 514400 182800
rect 514800 182400 515200 182800
rect 515600 182400 516000 182800
rect 516400 182400 572000 182800
rect 511500 182000 572000 182400
rect 511500 181600 512000 182000
rect 512400 181600 512800 182000
rect 513200 181600 513600 182000
rect 514000 181600 514400 182000
rect 514800 181600 515200 182000
rect 515600 181600 516000 182000
rect 516400 181600 572000 182000
rect 511500 181100 572000 181600
rect 573000 196230 584000 196500
rect 573000 191430 584800 196230
rect 573000 186230 584000 191430
rect 573000 181430 584800 186230
rect 573000 181100 584000 181430
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 0 38444 329400 42900
rect -800 38332 329400 38444
rect 0 37700 329400 38332
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 12020 549400 12540 564300
rect 11600 162800 13600 177900
rect 572000 181100 573000 196500
<< via3 >>
rect 16400 702000 16600 702200
rect 16800 702000 17000 702200
rect 17200 702000 17400 702200
rect 17600 702000 17800 702200
rect 18000 702000 18200 702200
rect 18400 702000 18600 702200
rect 18800 702000 19000 702200
rect 19200 702000 19400 702200
rect 19600 702000 19800 702200
rect 20000 702000 20200 702200
rect 20400 702000 20600 702200
rect 20800 702000 21000 702200
rect 23400 702060 23520 702180
rect 23600 702060 23720 702180
rect 23800 702060 23920 702180
rect 24000 702060 24120 702180
rect 24200 702060 24320 702180
rect 65060 702080 65240 702260
rect 65400 702080 65580 702260
rect 65740 702080 65920 702260
rect 16400 701600 16600 701800
rect 16800 701600 17000 701800
rect 17200 701600 17400 701800
rect 17600 701600 17800 701800
rect 18000 701600 18200 701800
rect 18400 701600 18600 701800
rect 18800 701600 19000 701800
rect 19200 701600 19400 701800
rect 19600 701600 19800 701800
rect 20000 701600 20200 701800
rect 20400 701600 20600 701800
rect 20800 701600 21000 701800
rect 16400 701200 16600 701400
rect 16800 701200 17000 701400
rect 17200 701200 17400 701400
rect 17600 701200 17800 701400
rect 18000 701200 18200 701400
rect 18400 701200 18600 701400
rect 18800 701200 19000 701400
rect 19200 701200 19400 701400
rect 19600 701200 19800 701400
rect 20000 701200 20200 701400
rect 20400 701200 20600 701400
rect 20800 701200 21000 701400
rect 16400 700800 16600 701000
rect 16800 700800 17000 701000
rect 17200 700800 17400 701000
rect 17600 700800 17800 701000
rect 18000 700800 18200 701000
rect 18400 700800 18600 701000
rect 18800 700800 19000 701000
rect 19200 700800 19400 701000
rect 19600 700800 19800 701000
rect 20000 700800 20200 701000
rect 20400 700800 20600 701000
rect 20800 700800 21000 701000
rect 16400 700400 16600 700600
rect 16800 700400 17000 700600
rect 17200 700400 17400 700600
rect 17600 700400 17800 700600
rect 18000 700400 18200 700600
rect 18400 700400 18600 700600
rect 18800 700400 19000 700600
rect 19200 700400 19400 700600
rect 19600 700400 19800 700600
rect 20000 700400 20200 700600
rect 20400 700400 20600 700600
rect 20800 700400 21000 700600
rect 16400 700000 16600 700200
rect 16800 700000 17000 700200
rect 17200 700000 17400 700200
rect 17600 700000 17800 700200
rect 18000 700000 18200 700200
rect 18400 700000 18600 700200
rect 18800 700000 19000 700200
rect 19200 700000 19400 700200
rect 19600 700000 19800 700200
rect 20000 700000 20200 700200
rect 20400 700000 20600 700200
rect 20800 700000 21000 700200
rect 68400 702000 68600 702200
rect 68800 702000 69000 702200
rect 69200 702000 69400 702200
rect 69600 702000 69800 702200
rect 70000 702000 70200 702200
rect 70400 702000 70600 702200
rect 70800 702000 71000 702200
rect 71200 702000 71400 702200
rect 71600 702000 71800 702200
rect 72000 702000 72200 702200
rect 72400 702000 72600 702200
rect 72800 702000 73000 702200
rect 68400 701600 68600 701800
rect 68800 701600 69000 701800
rect 69200 701600 69400 701800
rect 69600 701600 69800 701800
rect 70000 701600 70200 701800
rect 70400 701600 70600 701800
rect 70800 701600 71000 701800
rect 71200 701600 71400 701800
rect 71600 701600 71800 701800
rect 72000 701600 72200 701800
rect 72400 701600 72600 701800
rect 72800 701600 73000 701800
rect 68400 701200 68600 701400
rect 68800 701200 69000 701400
rect 69200 701200 69400 701400
rect 69600 701200 69800 701400
rect 70000 701200 70200 701400
rect 70400 701200 70600 701400
rect 70800 701200 71000 701400
rect 71200 701200 71400 701400
rect 71600 701200 71800 701400
rect 72000 701200 72200 701400
rect 72400 701200 72600 701400
rect 72800 701200 73000 701400
rect 68400 700800 68600 701000
rect 68800 700800 69000 701000
rect 69200 700800 69400 701000
rect 69600 700800 69800 701000
rect 70000 700800 70200 701000
rect 70400 700800 70600 701000
rect 70800 700800 71000 701000
rect 71200 700800 71400 701000
rect 71600 700800 71800 701000
rect 72000 700800 72200 701000
rect 72400 700800 72600 701000
rect 72800 700800 73000 701000
rect 68400 700400 68600 700600
rect 68800 700400 69000 700600
rect 69200 700400 69400 700600
rect 69600 700400 69800 700600
rect 70000 700400 70200 700600
rect 70400 700400 70600 700600
rect 70800 700400 71000 700600
rect 71200 700400 71400 700600
rect 71600 700400 71800 700600
rect 72000 700400 72200 700600
rect 72400 700400 72600 700600
rect 72800 700400 73000 700600
rect 68400 700000 68600 700200
rect 68800 700000 69000 700200
rect 69200 700000 69400 700200
rect 69600 700000 69800 700200
rect 70000 700000 70200 700200
rect 70400 700000 70600 700200
rect 70800 700000 71000 700200
rect 71200 700000 71400 700200
rect 71600 700000 71800 700200
rect 72000 700000 72200 700200
rect 72400 700000 72600 700200
rect 72800 700000 73000 700200
rect 13000 698000 13200 698200
rect 13600 698000 13800 698200
rect 23400 698000 23600 698200
rect 23800 698000 24000 698200
rect 24200 698000 24400 698200
rect 65000 698000 65200 698200
rect 65600 698000 65800 698200
rect 75400 698000 75600 698200
rect 76000 698000 76200 698200
rect 13000 697600 13200 697800
rect 13600 697600 13800 697800
rect 23400 697600 23600 697800
rect 23800 697600 24000 697800
rect 24200 697600 24400 697800
rect 65000 697600 65200 697800
rect 65600 697600 65800 697800
rect 75400 697600 75600 697800
rect 76000 697600 76200 697800
rect 23400 697200 23600 697400
rect 23800 697200 24000 697400
rect 24200 697200 24400 697400
rect 65000 697200 65200 697400
rect 65600 697200 65800 697400
rect 75400 697200 75600 697400
rect 76000 697200 76200 697400
rect 13000 697000 13200 697200
rect 13600 697000 13800 697200
rect 23400 696800 23600 697000
rect 23800 696800 24000 697000
rect 24200 696800 24400 697000
rect 65000 696800 65200 697000
rect 65600 696800 65800 697000
rect 75400 696800 75600 697000
rect 76000 696800 76200 697000
rect 13000 696600 13200 696800
rect 13600 696600 13800 696800
rect 23400 696400 23600 696600
rect 23800 696400 24000 696600
rect 24200 696400 24400 696600
rect 65000 696400 65200 696600
rect 65600 696400 65800 696600
rect 75400 696400 75600 696600
rect 76000 696400 76200 696600
rect 38700 692840 38860 693000
rect 39120 692840 39280 693000
rect 38700 692620 38860 692780
rect 39120 692620 39280 692780
rect 49960 692860 50100 693000
rect 50180 692860 50320 693000
rect 50400 692860 50540 693000
rect 49960 692660 50100 692800
rect 50180 692660 50320 692800
rect 50400 692660 50540 692800
rect 38700 692400 38860 692560
rect 39120 692400 39280 692560
rect 38700 692180 38860 692340
rect 39120 692180 39280 692340
rect 12900 691700 13100 691900
rect 13200 691700 13400 691900
rect 13500 691700 13700 691900
rect 13800 691700 14000 691900
rect 58000 691700 58200 691900
rect 58400 691700 58600 691900
rect 58800 691700 59000 691900
rect 59200 691700 59400 691900
rect 59600 691700 59800 691900
rect 60000 691700 60200 691900
rect 60400 691700 60600 691900
rect 60800 691700 61000 691900
rect 61200 691700 61400 691900
rect 61600 691700 61800 691900
rect 515700 701400 515900 701600
rect 516100 701400 516300 701600
rect 516500 701400 516700 701600
rect 516900 701400 517100 701600
rect 517300 701400 517500 701600
rect 517700 701400 517900 701600
rect 518100 701400 518300 701600
rect 518500 701400 518700 701600
rect 518900 701400 519100 701600
rect 519300 701400 519500 701600
rect 519700 701400 519900 701600
rect 520100 701400 520300 701600
rect 520500 701400 520700 701600
rect 515700 701000 515900 701200
rect 516100 701000 516300 701200
rect 516500 701000 516700 701200
rect 516900 701000 517100 701200
rect 517300 701000 517500 701200
rect 517700 701000 517900 701200
rect 518100 701000 518300 701200
rect 518500 701000 518700 701200
rect 518900 701000 519100 701200
rect 519300 701000 519500 701200
rect 519700 701000 519900 701200
rect 520100 701000 520300 701200
rect 520500 701000 520700 701200
rect 515700 700600 515900 700800
rect 516100 700600 516300 700800
rect 516500 700600 516700 700800
rect 516900 700600 517100 700800
rect 517300 700600 517500 700800
rect 517700 700600 517900 700800
rect 518100 700600 518300 700800
rect 518500 700600 518700 700800
rect 518900 700600 519100 700800
rect 519300 700600 519500 700800
rect 519700 700600 519900 700800
rect 520100 700600 520300 700800
rect 520500 700600 520700 700800
rect 515700 700200 515900 700400
rect 516100 700200 516300 700400
rect 516500 700200 516700 700400
rect 516900 700200 517100 700400
rect 517300 700200 517500 700400
rect 517700 700200 517900 700400
rect 518100 700200 518300 700400
rect 518500 700200 518700 700400
rect 518900 700200 519100 700400
rect 519300 700200 519500 700400
rect 519700 700200 519900 700400
rect 520100 700200 520300 700400
rect 520500 700200 520700 700400
rect 515700 699800 515900 700000
rect 516100 699800 516300 700000
rect 516500 699800 516700 700000
rect 516900 699800 517100 700000
rect 517300 699800 517500 700000
rect 517700 699800 517900 700000
rect 518100 699800 518300 700000
rect 518500 699800 518700 700000
rect 518900 699800 519100 700000
rect 519300 699800 519500 700000
rect 519700 699800 519900 700000
rect 520100 699800 520300 700000
rect 520500 699800 520700 700000
rect 515700 699400 515900 699600
rect 516100 699400 516300 699600
rect 516500 699400 516700 699600
rect 516900 699400 517100 699600
rect 517300 699400 517500 699600
rect 517700 699400 517900 699600
rect 518100 699400 518300 699600
rect 518500 699400 518700 699600
rect 518900 699400 519100 699600
rect 519300 699400 519500 699600
rect 519700 699400 519900 699600
rect 520100 699400 520300 699600
rect 520500 699400 520700 699600
rect 515700 699000 515900 699200
rect 516100 699000 516300 699200
rect 516500 699000 516700 699200
rect 516900 699000 517100 699200
rect 517300 699000 517500 699200
rect 517700 699000 517900 699200
rect 518100 699000 518300 699200
rect 518500 699000 518700 699200
rect 518900 699000 519100 699200
rect 519300 699000 519500 699200
rect 519700 699000 519900 699200
rect 520100 699000 520300 699200
rect 520500 699000 520700 699200
rect 515700 697200 515900 697400
rect 516100 697200 516300 697400
rect 516500 697200 516700 697400
rect 516900 697200 517100 697400
rect 517300 697200 517500 697400
rect 517700 697200 517900 697400
rect 518100 697200 518300 697400
rect 518500 697200 518700 697400
rect 518900 697200 519100 697400
rect 519300 697200 519500 697400
rect 519700 697200 519900 697400
rect 520100 697200 520300 697400
rect 520500 697200 520700 697400
rect 515700 696800 515900 697000
rect 516100 696800 516300 697000
rect 516500 696800 516700 697000
rect 516900 696800 517100 697000
rect 517300 696800 517500 697000
rect 517700 696800 517900 697000
rect 518100 696800 518300 697000
rect 518500 696800 518700 697000
rect 518900 696800 519100 697000
rect 519300 696800 519500 697000
rect 519700 696800 519900 697000
rect 520100 696800 520300 697000
rect 520500 696800 520700 697000
rect 515700 696400 515900 696600
rect 516100 696400 516300 696600
rect 516500 696400 516700 696600
rect 516900 696400 517100 696600
rect 517300 696400 517500 696600
rect 517700 696400 517900 696600
rect 518100 696400 518300 696600
rect 518500 696400 518700 696600
rect 518900 696400 519100 696600
rect 519300 696400 519500 696600
rect 519700 696400 519900 696600
rect 520100 696400 520300 696600
rect 520500 696400 520700 696600
rect 573300 697800 573500 698000
rect 573800 697800 574000 698000
rect 573300 697400 573500 697600
rect 573800 697400 574000 697600
rect 573300 697000 573500 697200
rect 573800 697000 574000 697200
rect 573300 696600 573500 696800
rect 573800 696600 574000 696800
rect 573300 696200 573500 696400
rect 573800 696200 574000 696400
rect 68400 690000 68600 690200
rect 68800 690000 69000 690200
rect 69200 690000 69400 690200
rect 69600 690000 69800 690200
rect 70000 690000 70200 690200
rect 70400 690000 70600 690200
rect 70800 690000 71000 690200
rect 71200 690000 71400 690200
rect 71600 690000 71800 690200
rect 72000 690000 72200 690200
rect 72400 690000 72600 690200
rect 72800 690000 73000 690200
rect 68400 689600 68600 689800
rect 68800 689600 69000 689800
rect 69200 689600 69400 689800
rect 69600 689600 69800 689800
rect 70000 689600 70200 689800
rect 70400 689600 70600 689800
rect 70800 689600 71000 689800
rect 71200 689600 71400 689800
rect 71600 689600 71800 689800
rect 72000 689600 72200 689800
rect 72400 689600 72600 689800
rect 72800 689600 73000 689800
rect 532300 690200 532500 690400
rect 532700 690200 532900 690400
rect 533100 690200 533300 690400
rect 533500 690200 533700 690400
rect 533900 690200 534100 690400
rect 532300 689900 532500 690100
rect 532700 689900 532900 690100
rect 533100 689900 533300 690100
rect 533500 689900 533700 690100
rect 533900 689900 534100 690100
rect 532300 689500 532500 689700
rect 532700 689500 532900 689700
rect 533100 689500 533300 689700
rect 533500 689500 533700 689700
rect 533900 689500 534100 689700
rect 532300 689100 532500 689300
rect 532700 689100 532900 689300
rect 533100 689100 533300 689300
rect 533500 689100 533700 689300
rect 533900 689100 534100 689300
rect 16400 688500 16600 688700
rect 16800 688500 17000 688700
rect 17200 688500 17400 688700
rect 17600 688500 17800 688700
rect 18000 688500 18200 688700
rect 18400 688500 18600 688700
rect 18800 688500 19000 688700
rect 19200 688500 19400 688700
rect 19600 688500 19800 688700
rect 20000 688500 20200 688700
rect 20400 688500 20600 688700
rect 20800 688500 21000 688700
rect 532300 688700 532500 688900
rect 532700 688700 532900 688900
rect 533100 688700 533300 688900
rect 533500 688700 533700 688900
rect 533900 688700 534100 688900
rect 16400 688100 16600 688300
rect 16800 688100 17000 688300
rect 17200 688100 17400 688300
rect 17600 688100 17800 688300
rect 18000 688100 18200 688300
rect 18400 688100 18600 688300
rect 18800 688100 19000 688300
rect 19200 688100 19400 688300
rect 19600 688100 19800 688300
rect 20000 688100 20200 688300
rect 20400 688100 20600 688300
rect 20800 688100 21000 688300
rect 36800 687100 37000 687300
rect 37200 687100 37400 687300
rect 37600 687100 37800 687300
rect 38000 687100 38200 687300
rect 549900 687000 550100 687200
rect 550200 687000 550400 687200
rect 550500 687000 550700 687200
rect 550800 687000 551000 687200
rect 551200 687100 551400 687300
rect 551200 686800 551400 687000
rect 551200 686500 551400 686700
rect 551200 686200 551400 686400
rect 549800 685900 550000 686100
rect 550100 685900 550300 686100
rect 550400 685900 550600 686100
rect 550800 685900 551000 686100
rect 36800 685100 37000 685300
rect 37200 685100 37400 685300
rect 37600 685100 37800 685300
rect 38000 685100 38200 685300
rect 36800 684700 37000 684900
rect 37200 684700 37400 684900
rect 37600 684700 37800 684900
rect 38000 684700 38200 684900
rect 36800 684300 37000 684500
rect 37200 684300 37400 684500
rect 37600 684300 37800 684500
rect 38000 684300 38200 684500
rect 36800 683900 37000 684100
rect 37200 683900 37400 684100
rect 37600 683900 37800 684100
rect 38000 683900 38200 684100
rect 36800 683500 37000 683700
rect 37200 683500 37400 683700
rect 37600 683500 37800 683700
rect 38000 683500 38200 683700
rect 36800 683100 37000 683300
rect 37200 683100 37400 683300
rect 37600 683100 37800 683300
rect 38000 683100 38200 683300
rect 515700 684600 515900 684800
rect 516100 684600 516300 684800
rect 516500 684600 516700 684800
rect 516900 684600 517100 684800
rect 517300 684600 517500 684800
rect 517700 684600 517900 684800
rect 518100 684600 518300 684800
rect 518500 684600 518700 684800
rect 518900 684600 519100 684800
rect 519300 684600 519500 684800
rect 519700 684600 519900 684800
rect 520100 684600 520300 684800
rect 520500 684600 520700 684800
rect 515700 684200 515900 684400
rect 516100 684200 516300 684400
rect 516500 684200 516700 684400
rect 516900 684200 517100 684400
rect 517300 684200 517500 684400
rect 517700 684200 517900 684400
rect 518100 684200 518300 684400
rect 518500 684200 518700 684400
rect 518900 684200 519100 684400
rect 519300 684200 519500 684400
rect 519700 684200 519900 684400
rect 520100 684200 520300 684400
rect 520500 684200 520700 684400
rect 515700 683800 515900 684000
rect 516100 683800 516300 684000
rect 516500 683800 516700 684000
rect 516900 683800 517100 684000
rect 517300 683800 517500 684000
rect 517700 683800 517900 684000
rect 518100 683800 518300 684000
rect 518500 683800 518700 684000
rect 518900 683800 519100 684000
rect 519300 683800 519500 684000
rect 519700 683800 519900 684000
rect 520100 683800 520300 684000
rect 520500 683800 520700 684000
rect 576800 684400 577100 684700
rect 577300 684400 577600 684700
rect 577800 684400 578100 684700
rect 578300 684400 578600 684700
rect 576800 683900 577100 684200
rect 577300 683900 577600 684200
rect 577800 683900 578100 684200
rect 578300 683900 578600 684200
rect 515700 683400 515900 683600
rect 516100 683400 516300 683600
rect 516500 683400 516700 683600
rect 516900 683400 517100 683600
rect 517300 683400 517500 683600
rect 517700 683400 517900 683600
rect 518100 683400 518300 683600
rect 518500 683400 518700 683600
rect 518900 683400 519100 683600
rect 519300 683400 519500 683600
rect 519700 683400 519900 683600
rect 520100 683400 520300 683600
rect 520500 683400 520700 683600
rect 36800 682700 37000 682900
rect 37200 682700 37400 682900
rect 37600 682700 37800 682900
rect 38000 682700 38200 682900
rect 36800 682300 37000 682500
rect 37200 682300 37400 682500
rect 37600 682300 37800 682500
rect 38000 682300 38200 682500
rect 515700 683000 515900 683200
rect 516100 683000 516300 683200
rect 516500 683000 516700 683200
rect 516900 683000 517100 683200
rect 517300 683000 517500 683200
rect 517700 683000 517900 683200
rect 518100 683000 518300 683200
rect 518500 683000 518700 683200
rect 518900 683000 519100 683200
rect 519300 683000 519500 683200
rect 519700 683000 519900 683200
rect 520100 683000 520300 683200
rect 520500 683000 520700 683200
rect 515700 682600 515900 682800
rect 516100 682600 516300 682800
rect 516500 682600 516700 682800
rect 516900 682600 517100 682800
rect 517300 682600 517500 682800
rect 517700 682600 517900 682800
rect 518100 682600 518300 682800
rect 518500 682600 518700 682800
rect 518900 682600 519100 682800
rect 519300 682600 519500 682800
rect 519700 682600 519900 682800
rect 520100 682600 520300 682800
rect 520500 682600 520700 682800
rect 36800 681900 37000 682100
rect 37200 681900 37400 682100
rect 37600 681900 37800 682100
rect 38000 681900 38200 682100
rect 58000 682000 58200 682200
rect 58400 682000 58600 682200
rect 58800 682000 59000 682200
rect 59200 682000 59400 682200
rect 59600 682000 59800 682200
rect 60000 682000 60200 682200
rect 60400 682000 60600 682200
rect 60800 682000 61000 682200
rect 61200 682000 61400 682200
rect 61600 682000 61800 682200
rect 36800 681500 37000 681700
rect 37200 681500 37400 681700
rect 37600 681500 37800 681700
rect 38000 681500 38200 681700
rect 36800 681100 37000 681300
rect 37200 681100 37400 681300
rect 37600 681100 37800 681300
rect 38000 681100 38200 681300
rect 36800 680700 37000 680900
rect 37200 680700 37400 680900
rect 37600 680700 37800 680900
rect 38000 680700 38200 680900
rect 549800 681200 550000 681400
rect 550200 681200 550400 681400
rect 550600 681200 550800 681400
rect 551000 681200 551200 681400
rect 551400 681200 551600 681400
rect 551800 681200 552000 681400
rect 552200 681200 552400 681400
rect 552600 681200 552800 681400
rect 549800 680800 550000 681000
rect 550200 680800 550400 681000
rect 550600 680800 550800 681000
rect 551000 680800 551200 681000
rect 551400 680800 551600 681000
rect 551800 680800 552000 681000
rect 552200 680800 552400 681000
rect 552600 680800 552800 681000
rect 36800 680300 37000 680500
rect 37200 680300 37400 680500
rect 37600 680300 37800 680500
rect 38000 680300 38200 680500
rect 515900 679000 516100 679200
rect 516300 679000 516500 679200
rect 516700 679000 516900 679200
rect 517100 679000 517300 679200
rect 517500 679000 517700 679200
rect 517900 679000 518100 679200
rect 518300 679000 518500 679200
rect 518700 679000 518900 679200
rect 519100 679000 519300 679200
rect 519500 679000 519700 679200
rect 519900 679000 520100 679200
rect 520300 679000 520500 679200
rect 520700 679000 520900 679200
rect 515900 678600 516100 678800
rect 516300 678600 516500 678800
rect 516700 678600 516900 678800
rect 517100 678600 517300 678800
rect 517500 678600 517700 678800
rect 517900 678600 518100 678800
rect 518300 678600 518500 678800
rect 518700 678600 518900 678800
rect 519100 678600 519300 678800
rect 519500 678600 519700 678800
rect 519900 678600 520100 678800
rect 520300 678600 520500 678800
rect 520700 678600 520900 678800
rect 515900 678200 516100 678400
rect 516300 678200 516500 678400
rect 516700 678200 516900 678400
rect 517100 678200 517300 678400
rect 517500 678200 517700 678400
rect 517900 678200 518100 678400
rect 518300 678200 518500 678400
rect 518700 678200 518900 678400
rect 519100 678200 519300 678400
rect 519500 678200 519700 678400
rect 519900 678200 520100 678400
rect 520300 678200 520500 678400
rect 520700 678200 520900 678400
rect 515900 677800 516100 678000
rect 516300 677800 516500 678000
rect 516700 677800 516900 678000
rect 517100 677800 517300 678000
rect 517500 677800 517700 678000
rect 517900 677800 518100 678000
rect 518300 677800 518500 678000
rect 518700 677800 518900 678000
rect 519100 677800 519300 678000
rect 519500 677800 519700 678000
rect 519900 677800 520100 678000
rect 520300 677800 520500 678000
rect 520700 677800 520900 678000
rect 515900 677400 516100 677600
rect 516300 677400 516500 677600
rect 516700 677400 516900 677600
rect 517100 677400 517300 677600
rect 517500 677400 517700 677600
rect 517900 677400 518100 677600
rect 518300 677400 518500 677600
rect 518700 677400 518900 677600
rect 519100 677400 519300 677600
rect 519500 677400 519700 677600
rect 519900 677400 520100 677600
rect 520300 677400 520500 677600
rect 520700 677400 520900 677600
rect 515900 677000 516100 677200
rect 516300 677000 516500 677200
rect 516700 677000 516900 677200
rect 517100 677000 517300 677200
rect 517500 677000 517700 677200
rect 517900 677000 518100 677200
rect 518300 677000 518500 677200
rect 518700 677000 518900 677200
rect 519100 677000 519300 677200
rect 519500 677000 519700 677200
rect 519900 677000 520100 677200
rect 520300 677000 520500 677200
rect 520700 677000 520900 677200
rect 515900 676600 516100 676800
rect 516300 676600 516500 676800
rect 516700 676600 516900 676800
rect 517100 676600 517300 676800
rect 517500 676600 517700 676800
rect 517900 676600 518100 676800
rect 518300 676600 518500 676800
rect 518700 676600 518900 676800
rect 519100 676600 519300 676800
rect 519500 676600 519700 676800
rect 519900 676600 520100 676800
rect 520300 676600 520500 676800
rect 520700 676600 520900 676800
rect 32800 663000 33100 663300
rect 33300 663000 33600 663300
rect 33800 663000 34100 663300
rect 34300 663000 34600 663300
rect 34800 663000 35100 663300
rect 35300 663000 35600 663300
rect 35800 663000 36100 663300
rect 36300 663000 36600 663300
rect 36800 663000 37100 663300
rect 37300 663000 37600 663300
rect 37800 663000 38100 663300
rect 38300 663000 38600 663300
rect 38800 663000 39100 663300
rect 39300 663000 39600 663300
rect 39800 663000 40100 663300
rect 40300 663000 40600 663300
rect 2500 648300 2800 648600
rect 3000 648300 3300 648600
rect 3500 648300 3800 648600
rect 2500 647800 2800 648100
rect 3000 647800 3300 648100
rect 3500 647800 3800 648100
rect 2500 647300 2800 647600
rect 3000 647300 3300 647600
rect 3500 647300 3800 647600
rect 2500 646800 2800 647100
rect 3000 646800 3300 647100
rect 3500 646800 3800 647100
rect 2500 646300 2800 646600
rect 3000 646300 3300 646600
rect 3500 646300 3800 646600
rect 2500 645800 2800 646100
rect 3000 645800 3300 646100
rect 3500 645800 3800 646100
rect 2500 645300 2800 645600
rect 3000 645300 3300 645600
rect 3500 645300 3800 645600
rect 2500 644800 2800 645100
rect 3000 644800 3300 645100
rect 3500 644800 3800 645100
rect 2500 644300 2800 644600
rect 3000 644300 3300 644600
rect 3500 644300 3800 644600
rect 2500 643800 2800 644100
rect 3000 643800 3300 644100
rect 3500 643800 3800 644100
rect 2500 643300 2800 643600
rect 3000 643300 3300 643600
rect 3500 643300 3800 643600
rect 2500 642800 2800 643100
rect 3000 642800 3300 643100
rect 3500 642800 3800 643100
rect 2500 642300 2800 642600
rect 3000 642300 3300 642600
rect 3500 642300 3800 642600
rect 2500 641800 2800 642100
rect 3000 641800 3300 642100
rect 3500 641800 3800 642100
rect 2500 641300 2800 641600
rect 3000 641300 3300 641600
rect 3500 641300 3800 641600
rect 2500 640800 2800 641100
rect 3000 640800 3300 641100
rect 3500 640800 3800 641100
rect 2500 640300 2800 640600
rect 3000 640300 3300 640600
rect 3500 640300 3800 640600
rect 2500 639800 2800 640100
rect 3000 639800 3300 640100
rect 3500 639800 3800 640100
rect 2500 639300 2800 639600
rect 3000 639300 3300 639600
rect 3500 639300 3800 639600
rect 2500 638800 2800 639100
rect 3000 638800 3300 639100
rect 3500 638800 3800 639100
rect 2500 638300 2800 638600
rect 3000 638300 3300 638600
rect 3500 638300 3800 638600
rect 2500 637800 2800 638100
rect 3000 637800 3300 638100
rect 3500 637800 3800 638100
rect 2500 637300 2800 637600
rect 3000 637300 3300 637600
rect 3500 637300 3800 637600
rect 2500 636800 2800 637100
rect 3000 636800 3300 637100
rect 3500 636800 3800 637100
rect 2500 636300 2800 636600
rect 3000 636300 3300 636600
rect 3500 636300 3800 636600
rect 2500 635800 2800 636100
rect 3000 635800 3300 636100
rect 3500 635800 3800 636100
rect 2500 635300 2800 635600
rect 3000 635300 3300 635600
rect 3500 635300 3800 635600
rect 2500 634800 2800 635100
rect 3000 634800 3300 635100
rect 3500 634800 3800 635100
rect 2500 634300 2800 634600
rect 3000 634300 3300 634600
rect 3500 634300 3800 634600
rect 550000 644400 550200 644600
rect 550400 644400 550600 644600
rect 550800 644400 551000 644600
rect 551200 644400 551400 644600
rect 551600 644400 551800 644600
rect 552000 644400 552200 644600
rect 552400 644400 552600 644600
rect 552800 644400 553000 644600
rect 550000 644000 550200 644200
rect 550400 644000 550600 644200
rect 550800 644000 551000 644200
rect 551200 644000 551400 644200
rect 551600 644000 551800 644200
rect 552000 644000 552200 644200
rect 552400 644000 552600 644200
rect 552800 644000 553000 644200
rect 550000 643600 550200 643800
rect 550400 643600 550600 643800
rect 550800 643600 551000 643800
rect 551200 643600 551400 643800
rect 551600 643600 551800 643800
rect 552000 643600 552200 643800
rect 552400 643600 552600 643800
rect 552800 643600 553000 643800
rect 550000 643200 550200 643400
rect 550400 643200 550600 643400
rect 550800 643200 551000 643400
rect 551200 643200 551400 643400
rect 551600 643200 551800 643400
rect 552000 643200 552200 643400
rect 552400 643200 552600 643400
rect 552800 643200 553000 643400
rect 550000 642800 550200 643000
rect 550400 642800 550600 643000
rect 550800 642800 551000 643000
rect 551200 642800 551400 643000
rect 551600 642800 551800 643000
rect 552000 642800 552200 643000
rect 552400 642800 552600 643000
rect 552800 642800 553000 643000
rect 550000 642400 550200 642600
rect 550400 642400 550600 642600
rect 550800 642400 551000 642600
rect 551200 642400 551400 642600
rect 551600 642400 551800 642600
rect 552000 642400 552200 642600
rect 552400 642400 552600 642600
rect 552800 642400 553000 642600
rect 550000 642000 550200 642200
rect 550400 642000 550600 642200
rect 550800 642000 551000 642200
rect 551200 642000 551400 642200
rect 551600 642000 551800 642200
rect 552000 642000 552200 642200
rect 552400 642000 552600 642200
rect 552800 642000 553000 642200
rect 550000 641600 550200 641800
rect 550400 641600 550600 641800
rect 550800 641600 551000 641800
rect 551200 641600 551400 641800
rect 551600 641600 551800 641800
rect 552000 641600 552200 641800
rect 552400 641600 552600 641800
rect 552800 641600 553000 641800
rect 550000 641200 550200 641400
rect 550400 641200 550600 641400
rect 550800 641200 551000 641400
rect 551200 641200 551400 641400
rect 551600 641200 551800 641400
rect 552000 641200 552200 641400
rect 552400 641200 552600 641400
rect 552800 641200 553000 641400
rect 550000 640800 550200 641000
rect 550400 640800 550600 641000
rect 550800 640800 551000 641000
rect 551200 640800 551400 641000
rect 551600 640800 551800 641000
rect 552000 640800 552200 641000
rect 552400 640800 552600 641000
rect 552800 640800 553000 641000
rect 550000 640400 550200 640600
rect 550400 640400 550600 640600
rect 550800 640400 551000 640600
rect 551200 640400 551400 640600
rect 551600 640400 551800 640600
rect 552000 640400 552200 640600
rect 552400 640400 552600 640600
rect 552800 640400 553000 640600
rect 550000 640000 550200 640200
rect 550400 640000 550600 640200
rect 550800 640000 551000 640200
rect 551200 640000 551400 640200
rect 551600 640000 551800 640200
rect 552000 640000 552200 640200
rect 552400 640000 552600 640200
rect 552800 640000 553000 640200
rect 550000 639600 550200 639800
rect 550400 639600 550600 639800
rect 550800 639600 551000 639800
rect 551200 639600 551400 639800
rect 551600 639600 551800 639800
rect 552000 639600 552200 639800
rect 552400 639600 552600 639800
rect 552800 639600 553000 639800
rect 550000 639200 550200 639400
rect 550400 639200 550600 639400
rect 550800 639200 551000 639400
rect 551200 639200 551400 639400
rect 551600 639200 551800 639400
rect 552000 639200 552200 639400
rect 552400 639200 552600 639400
rect 552800 639200 553000 639400
rect 550000 638800 550200 639000
rect 550400 638800 550600 639000
rect 550800 638800 551000 639000
rect 551200 638800 551400 639000
rect 551600 638800 551800 639000
rect 552000 638800 552200 639000
rect 552400 638800 552600 639000
rect 552800 638800 553000 639000
rect 550000 638400 550200 638600
rect 550400 638400 550600 638600
rect 550800 638400 551000 638600
rect 551200 638400 551400 638600
rect 551600 638400 551800 638600
rect 552000 638400 552200 638600
rect 552400 638400 552600 638600
rect 552800 638400 553000 638600
rect 550000 638000 550200 638200
rect 550400 638000 550600 638200
rect 550800 638000 551000 638200
rect 551200 638000 551400 638200
rect 551600 638000 551800 638200
rect 552000 638000 552200 638200
rect 552400 638000 552600 638200
rect 552800 638000 553000 638200
rect 550000 637600 550200 637800
rect 550400 637600 550600 637800
rect 550800 637600 551000 637800
rect 551200 637600 551400 637800
rect 551600 637600 551800 637800
rect 552000 637600 552200 637800
rect 552400 637600 552600 637800
rect 552800 637600 553000 637800
rect 550000 637200 550200 637400
rect 550400 637200 550600 637400
rect 550800 637200 551000 637400
rect 551200 637200 551400 637400
rect 551600 637200 551800 637400
rect 552000 637200 552200 637400
rect 552400 637200 552600 637400
rect 552800 637200 553000 637400
rect 550000 636800 550200 637000
rect 550400 636800 550600 637000
rect 550800 636800 551000 637000
rect 551200 636800 551400 637000
rect 551600 636800 551800 637000
rect 552000 636800 552200 637000
rect 552400 636800 552600 637000
rect 552800 636800 553000 637000
rect 550000 636400 550200 636600
rect 550400 636400 550600 636600
rect 550800 636400 551000 636600
rect 551200 636400 551400 636600
rect 551600 636400 551800 636600
rect 552000 636400 552200 636600
rect 552400 636400 552600 636600
rect 552800 636400 553000 636600
rect 550000 636000 550200 636200
rect 550400 636000 550600 636200
rect 550800 636000 551000 636200
rect 551200 636000 551400 636200
rect 551600 636000 551800 636200
rect 552000 636000 552200 636200
rect 552400 636000 552600 636200
rect 552800 636000 553000 636200
rect 550000 635600 550200 635800
rect 550400 635600 550600 635800
rect 550800 635600 551000 635800
rect 551200 635600 551400 635800
rect 551600 635600 551800 635800
rect 552000 635600 552200 635800
rect 552400 635600 552600 635800
rect 552800 635600 553000 635800
rect 550000 635200 550200 635400
rect 550400 635200 550600 635400
rect 550800 635200 551000 635400
rect 551200 635200 551400 635400
rect 551600 635200 551800 635400
rect 552000 635200 552200 635400
rect 552400 635200 552600 635400
rect 552800 635200 553000 635400
rect 550000 634800 550200 635000
rect 550400 634800 550600 635000
rect 550800 634800 551000 635000
rect 551200 634800 551400 635000
rect 551600 634800 551800 635000
rect 552000 634800 552200 635000
rect 552400 634800 552600 635000
rect 552800 634800 553000 635000
rect 550000 634400 550200 634600
rect 550400 634400 550600 634600
rect 550800 634400 551000 634600
rect 551200 634400 551400 634600
rect 551600 634400 551800 634600
rect 552000 634400 552200 634600
rect 552400 634400 552600 634600
rect 552800 634400 553000 634600
rect 550000 634000 550200 634200
rect 550400 634000 550600 634200
rect 550800 634000 551000 634200
rect 551200 634000 551400 634200
rect 551600 634000 551800 634200
rect 552000 634000 552200 634200
rect 552400 634000 552600 634200
rect 552800 634000 553000 634200
rect 550000 633600 550200 633800
rect 550400 633600 550600 633800
rect 550800 633600 551000 633800
rect 551200 633600 551400 633800
rect 551600 633600 551800 633800
rect 552000 633600 552200 633800
rect 552400 633600 552600 633800
rect 552800 633600 553000 633800
rect 550000 633200 550200 633400
rect 550400 633200 550600 633400
rect 550800 633200 551000 633400
rect 551200 633200 551400 633400
rect 551600 633200 551800 633400
rect 552000 633200 552200 633400
rect 552400 633200 552600 633400
rect 552800 633200 553000 633400
rect 550000 632800 550200 633000
rect 550400 632800 550600 633000
rect 550800 632800 551000 633000
rect 551200 632800 551400 633000
rect 551600 632800 551800 633000
rect 552000 632800 552200 633000
rect 552400 632800 552600 633000
rect 552800 632800 553000 633000
rect 550000 632400 550200 632600
rect 550400 632400 550600 632600
rect 550800 632400 551000 632600
rect 551200 632400 551400 632600
rect 551600 632400 551800 632600
rect 552000 632400 552200 632600
rect 552400 632400 552600 632600
rect 552800 632400 553000 632600
rect 550000 632000 550200 632200
rect 550400 632000 550600 632200
rect 550800 632000 551000 632200
rect 551200 632000 551400 632200
rect 551600 632000 551800 632200
rect 552000 632000 552200 632200
rect 552400 632000 552600 632200
rect 552800 632000 553000 632200
rect 550000 631600 550200 631800
rect 550400 631600 550600 631800
rect 550800 631600 551000 631800
rect 551200 631600 551400 631800
rect 551600 631600 551800 631800
rect 552000 631600 552200 631800
rect 552400 631600 552600 631800
rect 552800 631600 553000 631800
rect 550000 631200 550200 631400
rect 550400 631200 550600 631400
rect 550800 631200 551000 631400
rect 551200 631200 551400 631400
rect 551600 631200 551800 631400
rect 552000 631200 552200 631400
rect 552400 631200 552600 631400
rect 552800 631200 553000 631400
rect 550000 630800 550200 631000
rect 550400 630800 550600 631000
rect 550800 630800 551000 631000
rect 551200 630800 551400 631000
rect 551600 630800 551800 631000
rect 552000 630800 552200 631000
rect 552400 630800 552600 631000
rect 552800 630800 553000 631000
rect 550000 630500 550200 630700
rect 550400 630500 550600 630700
rect 550800 630500 551000 630700
rect 551200 630500 551400 630700
rect 551600 630500 551800 630700
rect 552000 630500 552200 630700
rect 552400 630500 552600 630700
rect 552800 630500 553000 630700
rect 550000 630200 550200 630400
rect 550400 630200 550600 630400
rect 550800 630200 551000 630400
rect 551200 630200 551400 630400
rect 551600 630200 551800 630400
rect 552000 630200 552200 630400
rect 552400 630200 552600 630400
rect 552800 630200 553000 630400
rect 550000 629800 550200 630000
rect 550400 629800 550600 630000
rect 550800 629800 551000 630000
rect 551200 629800 551400 630000
rect 551600 629800 551800 630000
rect 552000 629800 552200 630000
rect 552400 629800 552600 630000
rect 552800 629800 553000 630000
rect 282400 583400 282800 583800
rect 283200 583400 283600 583800
rect 282400 582600 282800 583000
rect 283200 582600 283600 583000
rect 282400 581800 282800 582200
rect 283200 581800 283600 582200
rect 282400 581000 282800 581400
rect 283200 581000 283600 581400
rect 282400 580200 282800 580600
rect 283200 580200 283600 580600
rect 282400 579400 282800 579800
rect 283200 579400 283600 579800
rect 32800 563900 33000 564100
rect 33200 563900 33400 564100
rect 33600 563900 33800 564100
rect 34000 563900 34200 564100
rect 34400 563900 34600 564100
rect 34800 563900 35000 564100
rect 35200 563900 35400 564100
rect 35600 563900 35800 564100
rect 36000 563900 36200 564100
rect 36400 563900 36600 564100
rect 36800 563900 37000 564100
rect 37200 563900 37400 564100
rect 37600 563900 37800 564100
rect 38000 563900 38200 564100
rect 38400 563900 38600 564100
rect 38800 563900 39000 564100
rect 39200 563900 39400 564100
rect 39600 563900 39800 564100
rect 40000 563900 40200 564100
rect 40400 563900 40600 564100
rect 32800 563500 33000 563700
rect 33200 563500 33400 563700
rect 33600 563500 33800 563700
rect 34000 563500 34200 563700
rect 34400 563500 34600 563700
rect 34800 563500 35000 563700
rect 35200 563500 35400 563700
rect 35600 563500 35800 563700
rect 36000 563500 36200 563700
rect 36400 563500 36600 563700
rect 36800 563500 37000 563700
rect 37200 563500 37400 563700
rect 37600 563500 37800 563700
rect 38000 563500 38200 563700
rect 38400 563500 38600 563700
rect 38800 563500 39000 563700
rect 39200 563500 39400 563700
rect 39600 563500 39800 563700
rect 40000 563500 40200 563700
rect 40400 563500 40600 563700
rect 32800 563100 33000 563300
rect 33200 563100 33400 563300
rect 33600 563100 33800 563300
rect 34000 563100 34200 563300
rect 34400 563100 34600 563300
rect 34800 563100 35000 563300
rect 35200 563100 35400 563300
rect 35600 563100 35800 563300
rect 36000 563100 36200 563300
rect 36400 563100 36600 563300
rect 36800 563100 37000 563300
rect 37200 563100 37400 563300
rect 37600 563100 37800 563300
rect 38000 563100 38200 563300
rect 38400 563100 38600 563300
rect 38800 563100 39000 563300
rect 39200 563100 39400 563300
rect 39600 563100 39800 563300
rect 40000 563100 40200 563300
rect 40400 563100 40600 563300
rect 32800 562700 33000 562900
rect 33200 562700 33400 562900
rect 33600 562700 33800 562900
rect 34000 562700 34200 562900
rect 34400 562700 34600 562900
rect 34800 562700 35000 562900
rect 35200 562700 35400 562900
rect 35600 562700 35800 562900
rect 36000 562700 36200 562900
rect 36400 562700 36600 562900
rect 36800 562700 37000 562900
rect 37200 562700 37400 562900
rect 37600 562700 37800 562900
rect 38000 562700 38200 562900
rect 38400 562700 38600 562900
rect 38800 562700 39000 562900
rect 39200 562700 39400 562900
rect 39600 562700 39800 562900
rect 40000 562700 40200 562900
rect 40400 562700 40600 562900
rect 32800 562300 33000 562500
rect 33200 562300 33400 562500
rect 33600 562300 33800 562500
rect 34000 562300 34200 562500
rect 34400 562300 34600 562500
rect 34800 562300 35000 562500
rect 35200 562300 35400 562500
rect 35600 562300 35800 562500
rect 36000 562300 36200 562500
rect 36400 562300 36600 562500
rect 36800 562300 37000 562500
rect 37200 562300 37400 562500
rect 37600 562300 37800 562500
rect 38000 562300 38200 562500
rect 38400 562300 38600 562500
rect 38800 562300 39000 562500
rect 39200 562300 39400 562500
rect 39600 562300 39800 562500
rect 40000 562300 40200 562500
rect 40400 562300 40600 562500
rect 32800 561900 33000 562100
rect 33200 561900 33400 562100
rect 33600 561900 33800 562100
rect 34000 561900 34200 562100
rect 34400 561900 34600 562100
rect 34800 561900 35000 562100
rect 35200 561900 35400 562100
rect 35600 561900 35800 562100
rect 36000 561900 36200 562100
rect 36400 561900 36600 562100
rect 36800 561900 37000 562100
rect 37200 561900 37400 562100
rect 37600 561900 37800 562100
rect 38000 561900 38200 562100
rect 38400 561900 38600 562100
rect 38800 561900 39000 562100
rect 39200 561900 39400 562100
rect 39600 561900 39800 562100
rect 40000 561900 40200 562100
rect 40400 561900 40600 562100
rect 32800 561500 33000 561700
rect 33200 561500 33400 561700
rect 33600 561500 33800 561700
rect 34000 561500 34200 561700
rect 34400 561500 34600 561700
rect 34800 561500 35000 561700
rect 35200 561500 35400 561700
rect 35600 561500 35800 561700
rect 36000 561500 36200 561700
rect 36400 561500 36600 561700
rect 36800 561500 37000 561700
rect 37200 561500 37400 561700
rect 37600 561500 37800 561700
rect 38000 561500 38200 561700
rect 38400 561500 38600 561700
rect 38800 561500 39000 561700
rect 39200 561500 39400 561700
rect 39600 561500 39800 561700
rect 40000 561500 40200 561700
rect 40400 561500 40600 561700
rect 32800 561100 33000 561300
rect 33200 561100 33400 561300
rect 33600 561100 33800 561300
rect 34000 561100 34200 561300
rect 34400 561100 34600 561300
rect 34800 561100 35000 561300
rect 35200 561100 35400 561300
rect 35600 561100 35800 561300
rect 36000 561100 36200 561300
rect 36400 561100 36600 561300
rect 36800 561100 37000 561300
rect 37200 561100 37400 561300
rect 37600 561100 37800 561300
rect 38000 561100 38200 561300
rect 38400 561100 38600 561300
rect 38800 561100 39000 561300
rect 39200 561100 39400 561300
rect 39600 561100 39800 561300
rect 40000 561100 40200 561300
rect 40400 561100 40600 561300
rect 32800 560700 33000 560900
rect 33200 560700 33400 560900
rect 33600 560700 33800 560900
rect 34000 560700 34200 560900
rect 34400 560700 34600 560900
rect 34800 560700 35000 560900
rect 35200 560700 35400 560900
rect 35600 560700 35800 560900
rect 36000 560700 36200 560900
rect 36400 560700 36600 560900
rect 36800 560700 37000 560900
rect 37200 560700 37400 560900
rect 37600 560700 37800 560900
rect 38000 560700 38200 560900
rect 38400 560700 38600 560900
rect 38800 560700 39000 560900
rect 39200 560700 39400 560900
rect 39600 560700 39800 560900
rect 40000 560700 40200 560900
rect 40400 560700 40600 560900
rect 32800 560300 33000 560500
rect 33200 560300 33400 560500
rect 33600 560300 33800 560500
rect 34000 560300 34200 560500
rect 34400 560300 34600 560500
rect 34800 560300 35000 560500
rect 35200 560300 35400 560500
rect 35600 560300 35800 560500
rect 36000 560300 36200 560500
rect 36400 560300 36600 560500
rect 36800 560300 37000 560500
rect 37200 560300 37400 560500
rect 37600 560300 37800 560500
rect 38000 560300 38200 560500
rect 38400 560300 38600 560500
rect 38800 560300 39000 560500
rect 39200 560300 39400 560500
rect 39600 560300 39800 560500
rect 40000 560300 40200 560500
rect 40400 560300 40600 560500
rect 32800 559900 33000 560100
rect 33200 559900 33400 560100
rect 33600 559900 33800 560100
rect 34000 559900 34200 560100
rect 34400 559900 34600 560100
rect 34800 559900 35000 560100
rect 35200 559900 35400 560100
rect 35600 559900 35800 560100
rect 36000 559900 36200 560100
rect 36400 559900 36600 560100
rect 36800 559900 37000 560100
rect 37200 559900 37400 560100
rect 37600 559900 37800 560100
rect 38000 559900 38200 560100
rect 38400 559900 38600 560100
rect 38800 559900 39000 560100
rect 39200 559900 39400 560100
rect 39600 559900 39800 560100
rect 40000 559900 40200 560100
rect 40400 559900 40600 560100
rect 32800 559500 33000 559700
rect 33200 559500 33400 559700
rect 33600 559500 33800 559700
rect 34000 559500 34200 559700
rect 34400 559500 34600 559700
rect 34800 559500 35000 559700
rect 35200 559500 35400 559700
rect 35600 559500 35800 559700
rect 36000 559500 36200 559700
rect 36400 559500 36600 559700
rect 36800 559500 37000 559700
rect 37200 559500 37400 559700
rect 37600 559500 37800 559700
rect 38000 559500 38200 559700
rect 38400 559500 38600 559700
rect 38800 559500 39000 559700
rect 39200 559500 39400 559700
rect 39600 559500 39800 559700
rect 40000 559500 40200 559700
rect 40400 559500 40600 559700
rect 32800 559100 33000 559300
rect 33200 559100 33400 559300
rect 33600 559100 33800 559300
rect 34000 559100 34200 559300
rect 34400 559100 34600 559300
rect 34800 559100 35000 559300
rect 35200 559100 35400 559300
rect 35600 559100 35800 559300
rect 36000 559100 36200 559300
rect 36400 559100 36600 559300
rect 36800 559100 37000 559300
rect 37200 559100 37400 559300
rect 37600 559100 37800 559300
rect 38000 559100 38200 559300
rect 38400 559100 38600 559300
rect 38800 559100 39000 559300
rect 39200 559100 39400 559300
rect 39600 559100 39800 559300
rect 40000 559100 40200 559300
rect 40400 559100 40600 559300
rect 32800 558700 33000 558900
rect 33200 558700 33400 558900
rect 33600 558700 33800 558900
rect 34000 558700 34200 558900
rect 34400 558700 34600 558900
rect 34800 558700 35000 558900
rect 35200 558700 35400 558900
rect 35600 558700 35800 558900
rect 36000 558700 36200 558900
rect 36400 558700 36600 558900
rect 36800 558700 37000 558900
rect 37200 558700 37400 558900
rect 37600 558700 37800 558900
rect 38000 558700 38200 558900
rect 38400 558700 38600 558900
rect 38800 558700 39000 558900
rect 39200 558700 39400 558900
rect 39600 558700 39800 558900
rect 40000 558700 40200 558900
rect 40400 558700 40600 558900
rect 32800 558300 33000 558500
rect 33200 558300 33400 558500
rect 33600 558300 33800 558500
rect 34000 558300 34200 558500
rect 34400 558300 34600 558500
rect 34800 558300 35000 558500
rect 35200 558300 35400 558500
rect 35600 558300 35800 558500
rect 36000 558300 36200 558500
rect 36400 558300 36600 558500
rect 36800 558300 37000 558500
rect 37200 558300 37400 558500
rect 37600 558300 37800 558500
rect 38000 558300 38200 558500
rect 38400 558300 38600 558500
rect 38800 558300 39000 558500
rect 39200 558300 39400 558500
rect 39600 558300 39800 558500
rect 40000 558300 40200 558500
rect 40400 558300 40600 558500
rect 32800 557900 33000 558100
rect 33200 557900 33400 558100
rect 33600 557900 33800 558100
rect 34000 557900 34200 558100
rect 34400 557900 34600 558100
rect 34800 557900 35000 558100
rect 35200 557900 35400 558100
rect 35600 557900 35800 558100
rect 36000 557900 36200 558100
rect 36400 557900 36600 558100
rect 36800 557900 37000 558100
rect 37200 557900 37400 558100
rect 37600 557900 37800 558100
rect 38000 557900 38200 558100
rect 38400 557900 38600 558100
rect 38800 557900 39000 558100
rect 39200 557900 39400 558100
rect 39600 557900 39800 558100
rect 40000 557900 40200 558100
rect 40400 557900 40600 558100
rect 32800 557500 33000 557700
rect 33200 557500 33400 557700
rect 33600 557500 33800 557700
rect 34000 557500 34200 557700
rect 34400 557500 34600 557700
rect 34800 557500 35000 557700
rect 35200 557500 35400 557700
rect 35600 557500 35800 557700
rect 36000 557500 36200 557700
rect 36400 557500 36600 557700
rect 36800 557500 37000 557700
rect 37200 557500 37400 557700
rect 37600 557500 37800 557700
rect 38000 557500 38200 557700
rect 38400 557500 38600 557700
rect 38800 557500 39000 557700
rect 39200 557500 39400 557700
rect 39600 557500 39800 557700
rect 40000 557500 40200 557700
rect 40400 557500 40600 557700
rect 32800 557100 33000 557300
rect 33200 557100 33400 557300
rect 33600 557100 33800 557300
rect 34000 557100 34200 557300
rect 34400 557100 34600 557300
rect 34800 557100 35000 557300
rect 35200 557100 35400 557300
rect 35600 557100 35800 557300
rect 36000 557100 36200 557300
rect 36400 557100 36600 557300
rect 36800 557100 37000 557300
rect 37200 557100 37400 557300
rect 37600 557100 37800 557300
rect 38000 557100 38200 557300
rect 38400 557100 38600 557300
rect 38800 557100 39000 557300
rect 39200 557100 39400 557300
rect 39600 557100 39800 557300
rect 40000 557100 40200 557300
rect 40400 557100 40600 557300
rect 32800 556700 33000 556900
rect 33200 556700 33400 556900
rect 33600 556700 33800 556900
rect 34000 556700 34200 556900
rect 34400 556700 34600 556900
rect 34800 556700 35000 556900
rect 35200 556700 35400 556900
rect 35600 556700 35800 556900
rect 36000 556700 36200 556900
rect 36400 556700 36600 556900
rect 36800 556700 37000 556900
rect 37200 556700 37400 556900
rect 37600 556700 37800 556900
rect 38000 556700 38200 556900
rect 38400 556700 38600 556900
rect 38800 556700 39000 556900
rect 39200 556700 39400 556900
rect 39600 556700 39800 556900
rect 40000 556700 40200 556900
rect 40400 556700 40600 556900
rect 32800 556300 33000 556500
rect 33200 556300 33400 556500
rect 33600 556300 33800 556500
rect 34000 556300 34200 556500
rect 34400 556300 34600 556500
rect 34800 556300 35000 556500
rect 35200 556300 35400 556500
rect 35600 556300 35800 556500
rect 36000 556300 36200 556500
rect 36400 556300 36600 556500
rect 36800 556300 37000 556500
rect 37200 556300 37400 556500
rect 37600 556300 37800 556500
rect 38000 556300 38200 556500
rect 38400 556300 38600 556500
rect 38800 556300 39000 556500
rect 39200 556300 39400 556500
rect 39600 556300 39800 556500
rect 40000 556300 40200 556500
rect 40400 556300 40600 556500
rect 32800 555900 33000 556100
rect 33200 555900 33400 556100
rect 33600 555900 33800 556100
rect 34000 555900 34200 556100
rect 34400 555900 34600 556100
rect 34800 555900 35000 556100
rect 35200 555900 35400 556100
rect 35600 555900 35800 556100
rect 36000 555900 36200 556100
rect 36400 555900 36600 556100
rect 36800 555900 37000 556100
rect 37200 555900 37400 556100
rect 37600 555900 37800 556100
rect 38000 555900 38200 556100
rect 38400 555900 38600 556100
rect 38800 555900 39000 556100
rect 39200 555900 39400 556100
rect 39600 555900 39800 556100
rect 40000 555900 40200 556100
rect 40400 555900 40600 556100
rect 32800 555500 33000 555700
rect 33200 555500 33400 555700
rect 33600 555500 33800 555700
rect 34000 555500 34200 555700
rect 34400 555500 34600 555700
rect 34800 555500 35000 555700
rect 35200 555500 35400 555700
rect 35600 555500 35800 555700
rect 36000 555500 36200 555700
rect 36400 555500 36600 555700
rect 36800 555500 37000 555700
rect 37200 555500 37400 555700
rect 37600 555500 37800 555700
rect 38000 555500 38200 555700
rect 38400 555500 38600 555700
rect 38800 555500 39000 555700
rect 39200 555500 39400 555700
rect 39600 555500 39800 555700
rect 40000 555500 40200 555700
rect 40400 555500 40600 555700
rect 32800 555100 33000 555300
rect 33200 555100 33400 555300
rect 33600 555100 33800 555300
rect 34000 555100 34200 555300
rect 34400 555100 34600 555300
rect 34800 555100 35000 555300
rect 35200 555100 35400 555300
rect 35600 555100 35800 555300
rect 36000 555100 36200 555300
rect 36400 555100 36600 555300
rect 36800 555100 37000 555300
rect 37200 555100 37400 555300
rect 37600 555100 37800 555300
rect 38000 555100 38200 555300
rect 38400 555100 38600 555300
rect 38800 555100 39000 555300
rect 39200 555100 39400 555300
rect 39600 555100 39800 555300
rect 40000 555100 40200 555300
rect 40400 555100 40600 555300
rect 32800 554700 33000 554900
rect 33200 554700 33400 554900
rect 33600 554700 33800 554900
rect 34000 554700 34200 554900
rect 34400 554700 34600 554900
rect 34800 554700 35000 554900
rect 35200 554700 35400 554900
rect 35600 554700 35800 554900
rect 36000 554700 36200 554900
rect 36400 554700 36600 554900
rect 36800 554700 37000 554900
rect 37200 554700 37400 554900
rect 37600 554700 37800 554900
rect 38000 554700 38200 554900
rect 38400 554700 38600 554900
rect 38800 554700 39000 554900
rect 39200 554700 39400 554900
rect 39600 554700 39800 554900
rect 40000 554700 40200 554900
rect 40400 554700 40600 554900
rect 32800 554300 33000 554500
rect 33200 554300 33400 554500
rect 33600 554300 33800 554500
rect 34000 554300 34200 554500
rect 34400 554300 34600 554500
rect 34800 554300 35000 554500
rect 35200 554300 35400 554500
rect 35600 554300 35800 554500
rect 36000 554300 36200 554500
rect 36400 554300 36600 554500
rect 36800 554300 37000 554500
rect 37200 554300 37400 554500
rect 37600 554300 37800 554500
rect 38000 554300 38200 554500
rect 38400 554300 38600 554500
rect 38800 554300 39000 554500
rect 39200 554300 39400 554500
rect 39600 554300 39800 554500
rect 40000 554300 40200 554500
rect 40400 554300 40600 554500
rect 32800 553900 33000 554100
rect 33200 553900 33400 554100
rect 33600 553900 33800 554100
rect 34000 553900 34200 554100
rect 34400 553900 34600 554100
rect 34800 553900 35000 554100
rect 35200 553900 35400 554100
rect 35600 553900 35800 554100
rect 36000 553900 36200 554100
rect 36400 553900 36600 554100
rect 36800 553900 37000 554100
rect 37200 553900 37400 554100
rect 37600 553900 37800 554100
rect 38000 553900 38200 554100
rect 38400 553900 38600 554100
rect 38800 553900 39000 554100
rect 39200 553900 39400 554100
rect 39600 553900 39800 554100
rect 40000 553900 40200 554100
rect 40400 553900 40600 554100
rect 32800 553500 33000 553700
rect 33200 553500 33400 553700
rect 33600 553500 33800 553700
rect 34000 553500 34200 553700
rect 34400 553500 34600 553700
rect 34800 553500 35000 553700
rect 35200 553500 35400 553700
rect 35600 553500 35800 553700
rect 36000 553500 36200 553700
rect 36400 553500 36600 553700
rect 36800 553500 37000 553700
rect 37200 553500 37400 553700
rect 37600 553500 37800 553700
rect 38000 553500 38200 553700
rect 38400 553500 38600 553700
rect 38800 553500 39000 553700
rect 39200 553500 39400 553700
rect 39600 553500 39800 553700
rect 40000 553500 40200 553700
rect 40400 553500 40600 553700
rect 32800 553100 33000 553300
rect 33200 553100 33400 553300
rect 33600 553100 33800 553300
rect 34000 553100 34200 553300
rect 34400 553100 34600 553300
rect 34800 553100 35000 553300
rect 35200 553100 35400 553300
rect 35600 553100 35800 553300
rect 36000 553100 36200 553300
rect 36400 553100 36600 553300
rect 36800 553100 37000 553300
rect 37200 553100 37400 553300
rect 37600 553100 37800 553300
rect 38000 553100 38200 553300
rect 38400 553100 38600 553300
rect 38800 553100 39000 553300
rect 39200 553100 39400 553300
rect 39600 553100 39800 553300
rect 40000 553100 40200 553300
rect 40400 553100 40600 553300
rect 32800 552700 33000 552900
rect 33200 552700 33400 552900
rect 33600 552700 33800 552900
rect 34000 552700 34200 552900
rect 34400 552700 34600 552900
rect 34800 552700 35000 552900
rect 35200 552700 35400 552900
rect 35600 552700 35800 552900
rect 36000 552700 36200 552900
rect 36400 552700 36600 552900
rect 36800 552700 37000 552900
rect 37200 552700 37400 552900
rect 37600 552700 37800 552900
rect 38000 552700 38200 552900
rect 38400 552700 38600 552900
rect 38800 552700 39000 552900
rect 39200 552700 39400 552900
rect 39600 552700 39800 552900
rect 40000 552700 40200 552900
rect 40400 552700 40600 552900
rect 32800 552300 33000 552500
rect 33200 552300 33400 552500
rect 33600 552300 33800 552500
rect 34000 552300 34200 552500
rect 34400 552300 34600 552500
rect 34800 552300 35000 552500
rect 35200 552300 35400 552500
rect 35600 552300 35800 552500
rect 36000 552300 36200 552500
rect 36400 552300 36600 552500
rect 36800 552300 37000 552500
rect 37200 552300 37400 552500
rect 37600 552300 37800 552500
rect 38000 552300 38200 552500
rect 38400 552300 38600 552500
rect 38800 552300 39000 552500
rect 39200 552300 39400 552500
rect 39600 552300 39800 552500
rect 40000 552300 40200 552500
rect 40400 552300 40600 552500
rect 32800 551900 33000 552100
rect 33200 551900 33400 552100
rect 33600 551900 33800 552100
rect 34000 551900 34200 552100
rect 34400 551900 34600 552100
rect 34800 551900 35000 552100
rect 35200 551900 35400 552100
rect 35600 551900 35800 552100
rect 36000 551900 36200 552100
rect 36400 551900 36600 552100
rect 36800 551900 37000 552100
rect 37200 551900 37400 552100
rect 37600 551900 37800 552100
rect 38000 551900 38200 552100
rect 38400 551900 38600 552100
rect 38800 551900 39000 552100
rect 39200 551900 39400 552100
rect 39600 551900 39800 552100
rect 40000 551900 40200 552100
rect 40400 551900 40600 552100
rect 32800 551500 33000 551700
rect 33200 551500 33400 551700
rect 33600 551500 33800 551700
rect 34000 551500 34200 551700
rect 34400 551500 34600 551700
rect 34800 551500 35000 551700
rect 35200 551500 35400 551700
rect 35600 551500 35800 551700
rect 36000 551500 36200 551700
rect 36400 551500 36600 551700
rect 36800 551500 37000 551700
rect 37200 551500 37400 551700
rect 37600 551500 37800 551700
rect 38000 551500 38200 551700
rect 38400 551500 38600 551700
rect 38800 551500 39000 551700
rect 39200 551500 39400 551700
rect 39600 551500 39800 551700
rect 40000 551500 40200 551700
rect 40400 551500 40600 551700
rect 32800 551100 33000 551300
rect 33200 551100 33400 551300
rect 33600 551100 33800 551300
rect 34000 551100 34200 551300
rect 34400 551100 34600 551300
rect 34800 551100 35000 551300
rect 35200 551100 35400 551300
rect 35600 551100 35800 551300
rect 36000 551100 36200 551300
rect 36400 551100 36600 551300
rect 36800 551100 37000 551300
rect 37200 551100 37400 551300
rect 37600 551100 37800 551300
rect 38000 551100 38200 551300
rect 38400 551100 38600 551300
rect 38800 551100 39000 551300
rect 39200 551100 39400 551300
rect 39600 551100 39800 551300
rect 40000 551100 40200 551300
rect 40400 551100 40600 551300
rect 32800 550700 33000 550900
rect 33200 550700 33400 550900
rect 33600 550700 33800 550900
rect 34000 550700 34200 550900
rect 34400 550700 34600 550900
rect 34800 550700 35000 550900
rect 35200 550700 35400 550900
rect 35600 550700 35800 550900
rect 36000 550700 36200 550900
rect 36400 550700 36600 550900
rect 36800 550700 37000 550900
rect 37200 550700 37400 550900
rect 37600 550700 37800 550900
rect 38000 550700 38200 550900
rect 38400 550700 38600 550900
rect 38800 550700 39000 550900
rect 39200 550700 39400 550900
rect 39600 550700 39800 550900
rect 40000 550700 40200 550900
rect 40400 550700 40600 550900
rect 32800 550300 33000 550500
rect 33200 550300 33400 550500
rect 33600 550300 33800 550500
rect 34000 550300 34200 550500
rect 34400 550300 34600 550500
rect 34800 550300 35000 550500
rect 35200 550300 35400 550500
rect 35600 550300 35800 550500
rect 36000 550300 36200 550500
rect 36400 550300 36600 550500
rect 36800 550300 37000 550500
rect 37200 550300 37400 550500
rect 37600 550300 37800 550500
rect 38000 550300 38200 550500
rect 38400 550300 38600 550500
rect 38800 550300 39000 550500
rect 39200 550300 39400 550500
rect 39600 550300 39800 550500
rect 40000 550300 40200 550500
rect 40400 550300 40600 550500
rect 32800 549900 33000 550100
rect 33200 549900 33400 550100
rect 33600 549900 33800 550100
rect 34000 549900 34200 550100
rect 34400 549900 34600 550100
rect 34800 549900 35000 550100
rect 35200 549900 35400 550100
rect 35600 549900 35800 550100
rect 36000 549900 36200 550100
rect 36400 549900 36600 550100
rect 36800 549900 37000 550100
rect 37200 549900 37400 550100
rect 37600 549900 37800 550100
rect 38000 549900 38200 550100
rect 38400 549900 38600 550100
rect 38800 549900 39000 550100
rect 39200 549900 39400 550100
rect 39600 549900 39800 550100
rect 40000 549900 40200 550100
rect 40400 549900 40600 550100
rect 32800 549500 33000 549700
rect 33200 549500 33400 549700
rect 33600 549500 33800 549700
rect 34000 549500 34200 549700
rect 34400 549500 34600 549700
rect 34800 549500 35000 549700
rect 35200 549500 35400 549700
rect 35600 549500 35800 549700
rect 36000 549500 36200 549700
rect 36400 549500 36600 549700
rect 36800 549500 37000 549700
rect 37200 549500 37400 549700
rect 37600 549500 37800 549700
rect 38000 549500 38200 549700
rect 38400 549500 38600 549700
rect 38800 549500 39000 549700
rect 39200 549500 39400 549700
rect 39600 549500 39800 549700
rect 40000 549500 40200 549700
rect 40400 549500 40600 549700
rect 285400 493800 285800 494200
rect 286200 493800 286600 494200
rect 285400 493000 285800 493400
rect 286200 493000 286600 493400
rect 285400 492200 285800 492600
rect 286200 492200 286600 492600
rect 285400 491400 285800 491800
rect 286200 491400 286600 491800
rect 285400 490600 285800 491000
rect 286200 490600 286600 491000
rect 285400 489800 285800 490200
rect 286200 489800 286600 490200
rect 288400 449400 288800 449800
rect 289200 449400 289600 449800
rect 288400 448600 288800 449000
rect 289200 448600 289600 449000
rect 288400 447800 288800 448200
rect 289200 447800 289600 448200
rect 288400 447000 288800 447400
rect 289200 447000 289600 447400
rect 288400 446200 288800 446600
rect 289200 446200 289600 446600
rect 288400 445400 288800 445800
rect 289200 445400 289600 445800
rect 291400 405000 291800 405400
rect 292200 405000 292600 405400
rect 291400 404200 291800 404600
rect 292200 404200 292600 404600
rect 291400 403400 291800 403800
rect 292200 403400 292600 403800
rect 291400 402600 291800 403000
rect 292200 402600 292600 403000
rect 291400 401800 291800 402200
rect 292200 401800 292600 402200
rect 291400 401000 291800 401400
rect 292200 401000 292600 401400
rect 294400 358600 294800 359000
rect 295200 358600 295600 359000
rect 294400 357800 294800 358200
rect 295200 357800 295600 358200
rect 294400 357000 294800 357400
rect 295200 357000 295600 357400
rect 294400 356200 294800 356600
rect 295200 356200 295600 356600
rect 294400 355400 294800 355800
rect 295200 355400 295600 355800
rect 294400 354600 294800 355000
rect 295200 354600 295600 355000
rect 9800 304180 10000 304200
rect 10200 304180 10400 304200
rect 10600 304180 10800 304200
rect 11000 304180 11200 304200
rect 11400 304180 11600 304200
rect 9800 304120 9845 304180
rect 9845 304120 9905 304180
rect 9905 304120 10000 304180
rect 10200 304120 10235 304180
rect 10235 304120 10295 304180
rect 10295 304120 10400 304180
rect 10600 304120 10615 304180
rect 10615 304120 10675 304180
rect 10675 304120 10800 304180
rect 11000 304120 11025 304180
rect 11025 304120 11155 304180
rect 11155 304120 11200 304180
rect 11400 304120 11470 304180
rect 11470 304120 11530 304180
rect 11530 304120 11600 304180
rect 9800 304000 10000 304120
rect 10200 304000 10400 304120
rect 10600 304000 10800 304120
rect 11000 304000 11200 304120
rect 11400 304000 11600 304120
rect 9800 303590 10000 303600
rect 10200 303590 10400 303600
rect 10600 303590 10800 303600
rect 11000 303590 11200 303600
rect 11400 303590 11600 303600
rect 9800 303530 9845 303590
rect 9845 303530 9905 303590
rect 9905 303530 10000 303590
rect 10200 303530 10235 303590
rect 10235 303530 10295 303590
rect 10295 303530 10400 303590
rect 10600 303530 10615 303590
rect 10615 303530 10675 303590
rect 10675 303530 10800 303590
rect 11000 303530 11025 303590
rect 11025 303530 11155 303590
rect 11155 303530 11200 303590
rect 11400 303530 11470 303590
rect 11470 303530 11530 303590
rect 11530 303530 11600 303590
rect 9800 303400 10000 303530
rect 10200 303400 10400 303530
rect 10600 303400 10800 303530
rect 11000 303400 11200 303530
rect 11400 303400 11600 303530
rect 5800 300800 6000 301000
rect 6200 300800 6400 301000
rect 6600 300800 6800 301000
rect 7000 300800 7200 301000
rect 7400 300800 7600 301000
rect 7800 300800 8000 301000
rect 5800 300400 6000 300600
rect 6200 300400 6400 300600
rect 6600 300400 6800 300600
rect 7000 300400 7200 300600
rect 7400 300400 7600 300600
rect 7800 300400 8000 300600
rect 5800 300000 6000 300200
rect 6200 300000 6400 300200
rect 6600 300000 6800 300200
rect 7000 300000 7200 300200
rect 7400 300000 7600 300200
rect 7800 300000 8000 300200
rect 5800 299600 6000 299800
rect 6200 299600 6400 299800
rect 6600 299600 6800 299800
rect 7000 299600 7200 299800
rect 7400 299600 7600 299800
rect 7800 299600 8000 299800
rect 5800 299200 6000 299400
rect 6200 299200 6400 299400
rect 6600 299200 6800 299400
rect 7000 299200 7200 299400
rect 7400 299200 7600 299400
rect 7800 299200 8000 299400
rect 5800 298800 6000 299000
rect 6200 298800 6400 299000
rect 6600 298800 6800 299000
rect 7000 298800 7200 299000
rect 7400 298800 7600 299000
rect 7800 298800 8000 299000
rect 5800 298400 6000 298600
rect 6200 298400 6400 298600
rect 6600 298400 6800 298600
rect 7000 298400 7200 298600
rect 7400 298400 7600 298600
rect 7800 298400 8000 298600
rect 5800 298000 6000 298200
rect 6200 298000 6400 298200
rect 6600 298000 6800 298200
rect 7000 298000 7200 298200
rect 7400 298000 7600 298200
rect 7800 298000 8000 298200
rect 5800 297600 6000 297800
rect 6200 297600 6400 297800
rect 6600 297600 6800 297800
rect 7000 297600 7200 297800
rect 7400 297600 7600 297800
rect 7800 297600 8000 297800
rect 5800 297200 6000 297400
rect 6200 297200 6400 297400
rect 6600 297200 6800 297400
rect 7000 297200 7200 297400
rect 7400 297200 7600 297400
rect 7800 297200 8000 297400
rect 5800 296800 6000 297000
rect 6200 296800 6400 297000
rect 6600 296800 6800 297000
rect 7000 296800 7200 297000
rect 7400 296800 7600 297000
rect 7800 296800 8000 297000
rect 5800 296400 6000 296600
rect 6200 296400 6400 296600
rect 6600 296400 6800 296600
rect 7000 296400 7200 296600
rect 7400 296400 7600 296600
rect 7800 296400 8000 296600
rect 17800 300800 18000 301000
rect 18200 300800 18400 301000
rect 17800 300400 18000 300600
rect 18200 300400 18400 300600
rect 17800 300000 18000 300200
rect 18200 300000 18400 300200
rect 17800 299600 18000 299800
rect 18200 299600 18400 299800
rect 17800 299200 18000 299400
rect 18200 299200 18400 299400
rect 294800 343900 295100 344200
rect 17800 298800 18000 299000
rect 18200 298800 18400 299000
rect 17800 298400 18000 298600
rect 18200 298400 18400 298600
rect 17800 298000 18000 298200
rect 18200 298000 18400 298200
rect 17800 297600 18000 297800
rect 18200 297600 18400 297800
rect 17800 297200 18000 297400
rect 18200 297200 18400 297400
rect 17800 296800 18000 297000
rect 18200 296800 18400 297000
rect 17800 296400 18000 296600
rect 18200 296400 18400 296600
rect 5740 293740 5920 293920
rect 9800 293780 10000 293800
rect 10200 293780 10400 293800
rect 10600 293780 10800 293800
rect 11000 293780 11200 293800
rect 11400 293780 11600 293800
rect 9800 293720 9845 293780
rect 9845 293720 9905 293780
rect 9905 293720 10000 293780
rect 10200 293720 10235 293780
rect 10235 293720 10295 293780
rect 10295 293720 10400 293780
rect 10600 293720 10615 293780
rect 10615 293720 10675 293780
rect 10675 293720 10800 293780
rect 11000 293720 11025 293780
rect 11025 293720 11155 293780
rect 11155 293720 11200 293780
rect 11400 293720 11470 293780
rect 11470 293720 11530 293780
rect 11530 293720 11600 293780
rect 9800 293600 10000 293720
rect 10200 293600 10400 293720
rect 10600 293600 10800 293720
rect 11000 293600 11200 293720
rect 11400 293600 11600 293720
rect 5740 293400 5920 293580
rect 5740 293060 5920 293240
rect 9800 293190 10000 293200
rect 10200 293190 10400 293200
rect 10600 293190 10800 293200
rect 11000 293190 11200 293200
rect 11400 293190 11600 293200
rect 9800 293130 9845 293190
rect 9845 293130 9905 293190
rect 9905 293130 10000 293190
rect 10200 293130 10235 293190
rect 10235 293130 10295 293190
rect 10295 293130 10400 293190
rect 10600 293130 10615 293190
rect 10615 293130 10675 293190
rect 10675 293130 10800 293190
rect 11000 293130 11025 293190
rect 11025 293130 11155 293190
rect 11155 293130 11200 293190
rect 11400 293130 11470 293190
rect 11470 293130 11530 293190
rect 11530 293130 11600 293190
rect 9800 293000 10000 293130
rect 10200 293000 10400 293130
rect 10600 293000 10800 293130
rect 11000 293000 11200 293130
rect 11400 293000 11600 293130
rect 13190 280430 13260 280500
rect 13080 280320 13150 280390
rect 6891 276678 6955 280022
rect 14540 278370 14640 278550
rect 15000 278400 15140 278540
rect 15200 278400 15340 278540
rect 15000 278180 15140 278320
rect 15200 278180 15340 278320
rect 14540 277950 14640 278130
rect 15000 277960 15140 278100
rect 15200 277960 15340 278100
rect 16100 289600 16300 289800
rect 16100 289200 16300 289400
rect 16100 288800 16300 289000
rect 16100 288400 16300 288600
rect 16100 288000 16300 288200
rect 16100 287600 16300 287800
rect 16100 287200 16300 287400
rect 16100 286800 16300 287000
rect 16100 286400 16300 286600
rect 16100 286000 16300 286200
rect 14040 276510 14140 276600
rect 14040 276320 14140 276410
rect 6891 272878 6955 276222
rect 12870 275220 13120 275470
rect 12360 273060 12630 273330
rect 12870 273320 13120 273570
rect 6891 269078 6955 272422
rect 12360 272010 12630 272280
rect 12870 271740 13120 271990
rect 12860 269850 13110 270090
rect 12860 269840 12910 269850
rect 12910 269840 13080 269850
rect 13080 269840 13110 269850
rect 14520 274120 14580 274130
rect 14580 274120 14720 274130
rect 14720 274120 14780 274130
rect 14520 273880 14780 274120
rect 14520 273870 14580 273880
rect 14580 273870 14720 273880
rect 14720 273870 14780 273880
rect 14000 273060 14270 273330
rect 14520 272860 14580 272870
rect 14580 272860 14720 272870
rect 14720 272860 14780 272870
rect 14520 272610 14780 272860
rect 14000 272010 14270 272280
rect 14520 271590 14580 271600
rect 14580 271590 14720 271600
rect 14720 271590 14780 271600
rect 14520 271350 14780 271590
rect 14520 271340 14580 271350
rect 14580 271340 14720 271350
rect 14720 271340 14780 271350
rect 25800 289600 26000 289800
rect 25800 289200 26000 289400
rect 25800 288800 26000 289000
rect 25800 288400 26000 288600
rect 25800 288000 26000 288200
rect 25800 287600 26000 287800
rect 25800 287200 26000 287400
rect 25800 286800 26000 287000
rect 25800 286400 26000 286600
rect 25800 286000 26000 286200
rect 16070 274120 16130 274130
rect 16130 274120 16270 274130
rect 16270 274120 16330 274130
rect 16070 273880 16330 274120
rect 16070 273870 16130 273880
rect 16130 273870 16270 273880
rect 16270 273870 16330 273880
rect 15610 273280 15870 273540
rect 16070 272860 16130 272870
rect 16130 272860 16270 272870
rect 16270 272860 16330 272870
rect 16070 272610 16330 272860
rect 15610 271780 15870 272040
rect 16070 271590 16130 271600
rect 16130 271590 16270 271600
rect 16270 271590 16330 271600
rect 16070 271350 16330 271590
rect 16070 271340 16130 271350
rect 16130 271340 16270 271350
rect 16270 271340 16330 271350
rect 18710 272520 18970 272780
rect 20230 272520 20490 272780
rect 21330 273560 21580 273810
rect 21750 272530 22000 272780
rect 21330 271500 21580 271750
rect 14040 268900 14140 268990
rect 14040 268710 14140 268800
rect 6891 265278 6955 268622
rect 14540 267120 14640 267300
rect 15000 267120 15160 267280
rect 15220 267120 15380 267280
rect 15440 267120 15600 267280
rect 15660 267120 15820 267280
rect 14540 266700 14640 266880
rect 15000 266700 15160 266860
rect 15220 266700 15380 266860
rect 15440 266700 15600 266860
rect 15660 266700 15820 266860
rect 13080 264930 13150 265000
rect 13190 264820 13260 264890
rect 9800 252380 10000 252400
rect 10200 252380 10400 252400
rect 10600 252380 10800 252400
rect 11000 252380 11200 252400
rect 11400 252380 11600 252400
rect 5820 252200 5940 252320
rect 9800 252320 9845 252380
rect 9845 252320 9905 252380
rect 9905 252320 10000 252380
rect 10200 252320 10235 252380
rect 10235 252320 10295 252380
rect 10295 252320 10400 252380
rect 10600 252320 10615 252380
rect 10615 252320 10675 252380
rect 10675 252320 10800 252380
rect 11000 252320 11025 252380
rect 11025 252320 11155 252380
rect 11155 252320 11200 252380
rect 11400 252320 11470 252380
rect 11470 252320 11530 252380
rect 11530 252320 11600 252380
rect 9800 252200 10000 252320
rect 10200 252200 10400 252320
rect 10600 252200 10800 252320
rect 11000 252200 11200 252320
rect 11400 252200 11600 252320
rect 5820 252000 5940 252120
rect 9800 251980 10000 252000
rect 10200 251980 10400 252000
rect 10600 251980 10800 252000
rect 11000 251980 11200 252000
rect 11400 251980 11600 252000
rect 5820 251800 5940 251920
rect 9800 251920 9845 251980
rect 9845 251920 9905 251980
rect 9905 251920 10000 251980
rect 10200 251920 10235 251980
rect 10235 251920 10295 251980
rect 10295 251920 10400 251980
rect 10600 251920 10615 251980
rect 10615 251920 10675 251980
rect 10675 251920 10800 251980
rect 11000 251920 11025 251980
rect 11025 251920 11155 251980
rect 11155 251920 11200 251980
rect 11400 251920 11470 251980
rect 11470 251920 11530 251980
rect 11530 251920 11600 251980
rect 9800 251800 10000 251920
rect 10200 251800 10400 251920
rect 10600 251800 10800 251920
rect 11000 251800 11200 251920
rect 11400 251800 11600 251920
rect 5820 251600 5940 251720
rect 9800 251590 10000 251600
rect 10200 251590 10400 251600
rect 10600 251590 10800 251600
rect 11000 251590 11200 251600
rect 11400 251590 11600 251600
rect 9800 251530 9845 251590
rect 9845 251530 9905 251590
rect 9905 251530 10000 251590
rect 10200 251530 10235 251590
rect 10235 251530 10295 251590
rect 10295 251530 10400 251590
rect 10600 251530 10615 251590
rect 10615 251530 10675 251590
rect 10675 251530 10800 251590
rect 11000 251530 11025 251590
rect 11025 251530 11155 251590
rect 11155 251530 11200 251590
rect 11400 251530 11470 251590
rect 11470 251530 11530 251590
rect 11530 251530 11600 251590
rect 5820 251400 5940 251520
rect 9800 251400 10000 251530
rect 10200 251400 10400 251530
rect 10600 251400 10800 251530
rect 11000 251400 11200 251530
rect 11400 251400 11600 251530
rect 5800 248800 6000 249000
rect 6200 248800 6400 249000
rect 6600 248800 6800 249000
rect 7000 248800 7200 249000
rect 7400 248800 7600 249000
rect 7800 248800 8000 249000
rect 5800 248400 6000 248600
rect 6200 248400 6400 248600
rect 6600 248400 6800 248600
rect 7000 248400 7200 248600
rect 7400 248400 7600 248600
rect 7800 248400 8000 248600
rect 5800 248000 6000 248200
rect 6200 248000 6400 248200
rect 6600 248000 6800 248200
rect 7000 248000 7200 248200
rect 7400 248000 7600 248200
rect 7800 248000 8000 248200
rect 5800 247600 6000 247800
rect 6200 247600 6400 247800
rect 6600 247600 6800 247800
rect 7000 247600 7200 247800
rect 7400 247600 7600 247800
rect 7800 247600 8000 247800
rect 5800 247200 6000 247400
rect 6200 247200 6400 247400
rect 6600 247200 6800 247400
rect 7000 247200 7200 247400
rect 7400 247200 7600 247400
rect 7800 247200 8000 247400
rect 5800 246800 6000 247000
rect 6200 246800 6400 247000
rect 6600 246800 6800 247000
rect 7000 246800 7200 247000
rect 7400 246800 7600 247000
rect 7800 246800 8000 247000
rect 5800 246400 6000 246600
rect 6200 246400 6400 246600
rect 6600 246400 6800 246600
rect 7000 246400 7200 246600
rect 7400 246400 7600 246600
rect 7800 246400 8000 246600
rect 5800 246000 6000 246200
rect 6200 246000 6400 246200
rect 6600 246000 6800 246200
rect 7000 246000 7200 246200
rect 7400 246000 7600 246200
rect 7800 246000 8000 246200
rect 5800 245600 6000 245800
rect 6200 245600 6400 245800
rect 6600 245600 6800 245800
rect 7000 245600 7200 245800
rect 7400 245600 7600 245800
rect 7800 245600 8000 245800
rect 5800 245200 6000 245400
rect 6200 245200 6400 245400
rect 6600 245200 6800 245400
rect 7000 245200 7200 245400
rect 7400 245200 7600 245400
rect 7800 245200 8000 245400
rect 5800 244800 6000 245000
rect 6200 244800 6400 245000
rect 6600 244800 6800 245000
rect 7000 244800 7200 245000
rect 7400 244800 7600 245000
rect 7800 244800 8000 245000
rect 5800 244400 6000 244600
rect 6200 244400 6400 244600
rect 6600 244400 6800 244600
rect 7000 244400 7200 244600
rect 7400 244400 7600 244600
rect 7800 244400 8000 244600
rect 22850 273820 23100 274070
rect 24400 273390 24480 273470
rect 24400 272870 24480 272950
rect 23280 272530 23530 272780
rect 24400 272350 24480 272430
rect 24380 271920 24500 271930
rect 24380 271840 24400 271920
rect 24400 271840 24480 271920
rect 24480 271840 24500 271920
rect 24380 271810 24500 271840
rect 34460 275900 34700 276140
rect 37660 275900 37900 276140
rect 40980 275900 41220 276140
rect 25860 273590 25940 273670
rect 26080 273590 26160 273670
rect 26220 273590 26300 273670
rect 22850 271240 23100 271490
rect 27470 272890 27590 273010
rect 28370 272590 28460 272680
rect 27480 272270 27600 272390
rect 28750 272580 28840 272670
rect 30190 272580 30280 272670
rect 288300 340500 288600 340800
rect 25860 271630 25940 271710
rect 26080 271630 26160 271710
rect 26220 271630 26300 271710
rect 34460 269200 34700 269440
rect 37660 269200 37900 269440
rect 40980 269200 41220 269440
rect 44700 268300 45000 268600
rect 44700 267800 45000 268100
rect 44700 267300 45000 267600
rect 44700 266800 45000 267100
rect 20700 266000 20900 266200
rect 20700 265600 20900 265800
rect 20700 265200 20900 265400
rect 20700 264800 20900 265000
rect 44700 266300 45000 266600
rect 22700 266000 22900 266200
rect 23100 266000 23300 266200
rect 23500 266000 23700 266200
rect 23900 266000 24100 266200
rect 24300 266000 24500 266200
rect 24700 266000 24900 266200
rect 25100 266000 25300 266200
rect 25500 266000 25700 266200
rect 25900 266000 26100 266200
rect 26300 266000 26500 266200
rect 26700 266000 26900 266200
rect 27100 266000 27300 266200
rect 27500 266000 27700 266200
rect 22700 265600 22900 265800
rect 23100 265600 23300 265800
rect 23500 265600 23700 265800
rect 23900 265600 24100 265800
rect 24300 265600 24500 265800
rect 24700 265600 24900 265800
rect 25100 265600 25300 265800
rect 25500 265600 25700 265800
rect 25900 265600 26100 265800
rect 26300 265600 26500 265800
rect 26700 265600 26900 265800
rect 27100 265600 27300 265800
rect 27500 265600 27700 265800
rect 44700 265800 45000 266100
rect 22700 265200 22900 265400
rect 23100 265200 23300 265400
rect 23500 265200 23700 265400
rect 23900 265200 24100 265400
rect 24300 265200 24500 265400
rect 24700 265200 24900 265400
rect 25100 265200 25300 265400
rect 25500 265200 25700 265400
rect 25900 265200 26100 265400
rect 26300 265200 26500 265400
rect 26700 265200 26900 265400
rect 27100 265200 27300 265400
rect 27500 265200 27700 265400
rect 44700 265300 45000 265600
rect 22700 264800 22900 265000
rect 23100 264800 23300 265000
rect 23500 264800 23700 265000
rect 23900 264800 24100 265000
rect 24300 264800 24500 265000
rect 24700 264800 24900 265000
rect 25100 264800 25300 265000
rect 25500 264800 25700 265000
rect 25900 264800 26100 265000
rect 26300 264800 26500 265000
rect 26700 264800 26900 265000
rect 27100 264800 27300 265000
rect 27500 264800 27700 265000
rect 19300 248800 19500 249000
rect 19700 248800 19900 249000
rect 19300 248400 19500 248600
rect 19700 248400 19900 248600
rect 19300 248000 19500 248200
rect 19700 248000 19900 248200
rect 19300 247600 19500 247800
rect 19700 247600 19900 247800
rect 19300 247200 19500 247400
rect 19700 247200 19900 247400
rect 19300 246800 19500 247000
rect 19700 246800 19900 247000
rect 19300 246400 19500 246600
rect 19700 246400 19900 246600
rect 19300 246000 19500 246200
rect 19700 246000 19900 246200
rect 19300 245600 19500 245800
rect 19700 245600 19900 245800
rect 19300 245200 19500 245400
rect 19700 245200 19900 245400
rect 19300 244800 19500 245000
rect 19700 244800 19900 245000
rect 19300 244400 19500 244600
rect 19700 244400 19900 244600
rect 44700 264800 45000 265100
rect 44700 264300 45000 264600
rect 44700 263800 45000 264100
rect 44700 263300 45000 263600
rect 44700 262800 45000 263100
rect 44700 262300 45000 262600
rect 44700 261800 45000 262100
rect 44700 261300 45000 261600
rect 44700 260800 45000 261100
rect 9800 241780 10000 241800
rect 10200 241780 10400 241800
rect 10800 241780 11000 241800
rect 11200 241780 11400 241800
rect 16100 241800 16300 242000
rect 9800 241720 9845 241780
rect 9845 241720 9905 241780
rect 9905 241720 10000 241780
rect 10200 241720 10235 241780
rect 10235 241720 10295 241780
rect 10295 241720 10400 241780
rect 10800 241720 10805 241780
rect 10805 241720 10865 241780
rect 10865 241720 10965 241780
rect 10965 241720 11000 241780
rect 11200 241720 11215 241780
rect 11215 241720 11330 241780
rect 11330 241720 11390 241780
rect 11390 241720 11400 241780
rect 9800 241600 10000 241720
rect 10200 241600 10400 241720
rect 10800 241600 11000 241720
rect 11200 241600 11400 241720
rect 16100 241500 16300 241700
rect 9800 241190 10000 241200
rect 10200 241190 10400 241200
rect 10800 241190 11000 241200
rect 11200 241190 11400 241200
rect 16100 241200 16300 241400
rect 9800 241130 9845 241190
rect 9845 241130 9905 241190
rect 9905 241130 10000 241190
rect 10200 241130 10235 241190
rect 10235 241130 10295 241190
rect 10295 241130 10400 241190
rect 10800 241130 10805 241190
rect 10805 241130 10865 241190
rect 10865 241130 10965 241190
rect 10965 241130 11000 241190
rect 11200 241130 11215 241190
rect 11215 241130 11330 241190
rect 11330 241130 11390 241190
rect 11390 241130 11400 241190
rect 9800 241000 10000 241130
rect 10200 241000 10400 241130
rect 10800 241000 11000 241130
rect 11200 241000 11400 241130
rect 16100 240900 16300 241100
rect 285400 219000 285800 219400
rect 286200 219000 286600 219400
rect 287000 219000 287400 219400
rect 287800 219000 288200 219400
rect 288600 219000 289000 219400
rect 289400 219000 289800 219400
rect 60000 218400 60400 218800
rect 60800 218400 61200 218800
rect 61600 218400 62000 218800
rect 62400 218400 62800 218800
rect 63200 218400 63600 218800
rect 64000 218400 64400 218800
rect 69000 218400 69400 218800
rect 69800 218400 70200 218800
rect 70600 218400 71000 218800
rect 71400 218400 71800 218800
rect 72200 218400 72600 218800
rect 73000 218400 73400 218800
rect 285400 218200 285800 218600
rect 286200 218200 286600 218600
rect 287000 218200 287400 218600
rect 287800 218200 288200 218600
rect 288600 218200 289000 218600
rect 289400 218200 289800 218600
rect 60000 217600 60400 218000
rect 60800 217600 61200 218000
rect 61600 217600 62000 218000
rect 62400 217600 62800 218000
rect 63200 217600 63600 218000
rect 64000 217600 64400 218000
rect 69000 217600 69400 218000
rect 69800 217600 70200 218000
rect 70600 217600 71000 218000
rect 71400 217600 71800 218000
rect 72200 217600 72600 218000
rect 73000 217600 73400 218000
rect 285400 217400 285800 217800
rect 286200 217400 286600 217800
rect 287000 217400 287400 217800
rect 287800 217400 288200 217800
rect 288600 217400 289000 217800
rect 289400 217400 289800 217800
rect 60000 216800 60400 217200
rect 60800 216800 61200 217200
rect 61600 216800 62000 217200
rect 62400 216800 62800 217200
rect 63200 216800 63600 217200
rect 64000 216800 64400 217200
rect 69000 216800 69400 217200
rect 69800 216800 70200 217200
rect 70600 216800 71000 217200
rect 71400 216800 71800 217200
rect 72200 216800 72600 217200
rect 73000 216800 73400 217200
rect 285400 216600 285800 217000
rect 286200 216600 286600 217000
rect 287000 216600 287400 217000
rect 287800 216600 288200 217000
rect 288600 216600 289000 217000
rect 289400 216600 289800 217000
rect 60000 216000 60400 216400
rect 60800 216000 61200 216400
rect 61600 216000 62000 216400
rect 62400 216000 62800 216400
rect 63200 216000 63600 216400
rect 64000 216000 64400 216400
rect 69000 216000 69400 216400
rect 69800 216000 70200 216400
rect 70600 216000 71000 216400
rect 71400 216000 71800 216400
rect 72200 216000 72600 216400
rect 73000 216000 73400 216400
rect 285400 215800 285800 216200
rect 286200 215800 286600 216200
rect 287000 215800 287400 216200
rect 287800 215800 288200 216200
rect 288600 215800 289000 216200
rect 289400 215800 289800 216200
rect 60000 215200 60400 215600
rect 60800 215200 61200 215600
rect 61600 215200 62000 215600
rect 62400 215200 62800 215600
rect 63200 215200 63600 215600
rect 64000 215200 64400 215600
rect 69000 215200 69400 215600
rect 69800 215200 70200 215600
rect 70600 215200 71000 215600
rect 71400 215200 71800 215600
rect 72200 215200 72600 215600
rect 73000 215200 73400 215600
rect 285400 215000 285800 215400
rect 286200 215000 286600 215400
rect 287000 215000 287400 215400
rect 287800 215000 288200 215400
rect 288600 215000 289000 215400
rect 289400 215000 289800 215400
rect 60000 214400 60400 214800
rect 60800 214400 61200 214800
rect 61600 214400 62000 214800
rect 62400 214400 62800 214800
rect 63200 214400 63600 214800
rect 64000 214400 64400 214800
rect 69000 214400 69400 214800
rect 69800 214400 70200 214800
rect 70600 214400 71000 214800
rect 71400 214400 71800 214800
rect 72200 214400 72600 214800
rect 73000 214400 73400 214800
rect 285200 214200 285600 214600
rect 286000 214200 286400 214600
rect 286800 214200 287200 214600
rect 287600 214200 288000 214600
rect 288400 214200 288800 214600
rect 289200 214200 289600 214600
rect 285200 213400 285600 213800
rect 286000 213400 286400 213800
rect 286800 213400 287200 213800
rect 287600 213400 288000 213800
rect 288400 213400 288800 213800
rect 289200 213400 289600 213800
rect 285200 212600 285600 213000
rect 286000 212600 286400 213000
rect 286800 212600 287200 213000
rect 287600 212600 288000 213000
rect 288400 212600 288800 213000
rect 289200 212600 289600 213000
rect 285200 211800 285600 212200
rect 286000 211800 286400 212200
rect 286800 211800 287200 212200
rect 287600 211800 288000 212200
rect 288400 211800 288800 212200
rect 289200 211800 289600 212200
rect 285200 211000 285600 211400
rect 286000 211000 286400 211400
rect 286800 211000 287200 211400
rect 287600 211000 288000 211400
rect 288400 211000 288800 211400
rect 289200 211000 289600 211400
rect 285200 210200 285600 210600
rect 286000 210200 286400 210600
rect 286800 210200 287200 210600
rect 287600 210200 288000 210600
rect 288400 210200 288800 210600
rect 289200 210200 289600 210600
rect 60000 209600 60400 210000
rect 60800 209600 61200 210000
rect 61600 209600 62000 210000
rect 62400 209600 62800 210000
rect 63200 209600 63600 210000
rect 64000 209600 64400 210000
rect 69000 209800 69400 210200
rect 69800 209800 70200 210200
rect 70600 209800 71000 210200
rect 71400 209800 71800 210200
rect 72200 209800 72600 210200
rect 73000 209800 73400 210200
rect 285200 209400 285600 209800
rect 286000 209400 286400 209800
rect 286800 209400 287200 209800
rect 287600 209400 288000 209800
rect 288400 209400 288800 209800
rect 289200 209400 289600 209800
rect 60000 208800 60400 209200
rect 60800 208800 61200 209200
rect 61600 208800 62000 209200
rect 62400 208800 62800 209200
rect 63200 208800 63600 209200
rect 64000 208800 64400 209200
rect 69000 209000 69400 209400
rect 69800 209000 70200 209400
rect 70600 209000 71000 209400
rect 71400 209000 71800 209400
rect 72200 209000 72600 209400
rect 73000 209000 73400 209400
rect 285200 208600 285600 209000
rect 286000 208600 286400 209000
rect 286800 208600 287200 209000
rect 287600 208600 288000 209000
rect 288400 208600 288800 209000
rect 289200 208600 289600 209000
rect 60000 208000 60400 208400
rect 60800 208000 61200 208400
rect 61600 208000 62000 208400
rect 62400 208000 62800 208400
rect 63200 208000 63600 208400
rect 64000 208000 64400 208400
rect 69000 208200 69400 208600
rect 69800 208200 70200 208600
rect 70600 208200 71000 208600
rect 71400 208200 71800 208600
rect 72200 208200 72600 208600
rect 73000 208200 73400 208600
rect 285200 207800 285600 208200
rect 286000 207800 286400 208200
rect 286800 207800 287200 208200
rect 287600 207800 288000 208200
rect 288400 207800 288800 208200
rect 289200 207800 289600 208200
rect 60000 207200 60400 207600
rect 60800 207200 61200 207600
rect 61600 207200 62000 207600
rect 62400 207200 62800 207600
rect 63200 207200 63600 207600
rect 64000 207200 64400 207600
rect 69000 207400 69400 207800
rect 69800 207400 70200 207800
rect 70600 207400 71000 207800
rect 71400 207400 71800 207800
rect 72200 207400 72600 207800
rect 73000 207400 73400 207800
rect 285200 207000 285600 207400
rect 286000 207000 286400 207400
rect 286800 207000 287200 207400
rect 287600 207000 288000 207400
rect 288400 207000 288800 207400
rect 289200 207000 289600 207400
rect 60000 206400 60400 206800
rect 60800 206400 61200 206800
rect 61600 206400 62000 206800
rect 62400 206400 62800 206800
rect 63200 206400 63600 206800
rect 64000 206400 64400 206800
rect 69000 206600 69400 207000
rect 69800 206600 70200 207000
rect 70600 206600 71000 207000
rect 71400 206600 71800 207000
rect 72200 206600 72600 207000
rect 73000 206600 73400 207000
rect 285200 206200 285600 206600
rect 286000 206200 286400 206600
rect 286800 206200 287200 206600
rect 287600 206200 288000 206600
rect 288400 206200 288800 206600
rect 289200 206200 289600 206600
rect 60000 205600 60400 206000
rect 60800 205600 61200 206000
rect 61600 205600 62000 206000
rect 62400 205600 62800 206000
rect 63200 205600 63600 206000
rect 64000 205600 64400 206000
rect 69000 205800 69400 206200
rect 69800 205800 70200 206200
rect 70600 205800 71000 206200
rect 71400 205800 71800 206200
rect 72200 205800 72600 206200
rect 73000 205800 73400 206200
rect 285200 205400 285600 205800
rect 286000 205400 286400 205800
rect 286800 205400 287200 205800
rect 287600 205400 288000 205800
rect 288400 205400 288800 205800
rect 289200 205400 289600 205800
rect 86000 177200 86400 177600
rect 86800 177200 87200 177600
rect 87600 177200 88000 177600
rect 88400 177200 88800 177600
rect 89200 177200 89600 177600
rect 90000 177200 90400 177600
rect 299400 177200 299800 177600
rect 300200 177200 300600 177600
rect 301000 177200 301400 177600
rect 301800 177200 302200 177600
rect 302600 177200 303000 177600
rect 303400 177200 303800 177600
rect 86000 176400 86400 176800
rect 86800 176400 87200 176800
rect 87600 176400 88000 176800
rect 88400 176400 88800 176800
rect 89200 176400 89600 176800
rect 90000 176400 90400 176800
rect 299400 176400 299800 176800
rect 300200 176400 300600 176800
rect 301000 176400 301400 176800
rect 301800 176400 302200 176800
rect 302600 176400 303000 176800
rect 303400 176400 303800 176800
rect 86000 175600 86400 176000
rect 86800 175600 87200 176000
rect 87600 175600 88000 176000
rect 88400 175600 88800 176000
rect 89200 175600 89600 176000
rect 90000 175600 90400 176000
rect 299400 175600 299800 176000
rect 300200 175600 300600 176000
rect 301000 175600 301400 176000
rect 301800 175600 302200 176000
rect 302600 175600 303000 176000
rect 303400 175600 303800 176000
rect 86000 174800 86400 175200
rect 86800 174800 87200 175200
rect 87600 174800 88000 175200
rect 88400 174800 88800 175200
rect 89200 174800 89600 175200
rect 90000 174800 90400 175200
rect 299400 174800 299800 175200
rect 300200 174800 300600 175200
rect 301000 174800 301400 175200
rect 301800 174800 302200 175200
rect 302600 174800 303000 175200
rect 303400 174800 303800 175200
rect 86000 174000 86400 174400
rect 86800 174000 87200 174400
rect 87600 174000 88000 174400
rect 88400 174000 88800 174400
rect 89200 174000 89600 174400
rect 90000 174000 90400 174400
rect 299400 174000 299800 174400
rect 300200 174000 300600 174400
rect 301000 174000 301400 174400
rect 301800 174000 302200 174400
rect 302600 174000 303000 174400
rect 303400 174000 303800 174400
rect 86000 173200 86400 173600
rect 86800 173200 87200 173600
rect 87600 173200 88000 173600
rect 88400 173200 88800 173600
rect 89200 173200 89600 173600
rect 90000 173200 90400 173600
rect 299400 173200 299800 173600
rect 300200 173200 300600 173600
rect 301000 173200 301400 173600
rect 301800 173200 302200 173600
rect 302600 173200 303000 173600
rect 303400 173200 303800 173600
rect 86000 172400 86400 172800
rect 86800 172400 87200 172800
rect 87600 172400 88000 172800
rect 88400 172400 88800 172800
rect 89200 172400 89600 172800
rect 90000 172400 90400 172800
rect 299400 172400 299800 172800
rect 300200 172400 300600 172800
rect 301000 172400 301400 172800
rect 301800 172400 302200 172800
rect 302600 172400 303000 172800
rect 303400 172400 303800 172800
rect 86000 171600 86400 172000
rect 86800 171600 87200 172000
rect 87600 171600 88000 172000
rect 88400 171600 88800 172000
rect 89200 171600 89600 172000
rect 90000 171600 90400 172000
rect 299400 171600 299800 172000
rect 300200 171600 300600 172000
rect 301000 171600 301400 172000
rect 301800 171600 302200 172000
rect 302600 171600 303000 172000
rect 303400 171600 303800 172000
rect 86000 170800 86400 171200
rect 86800 170800 87200 171200
rect 87600 170800 88000 171200
rect 88400 170800 88800 171200
rect 89200 170800 89600 171200
rect 90000 170800 90400 171200
rect 299400 170800 299800 171200
rect 300200 170800 300600 171200
rect 301000 170800 301400 171200
rect 301800 170800 302200 171200
rect 302600 170800 303000 171200
rect 303400 170800 303800 171200
rect 86000 170000 86400 170400
rect 86800 170000 87200 170400
rect 87600 170000 88000 170400
rect 88400 170000 88800 170400
rect 89200 170000 89600 170400
rect 90000 170000 90400 170400
rect 299400 170000 299800 170400
rect 300200 170000 300600 170400
rect 301000 170000 301400 170400
rect 301800 170000 302200 170400
rect 302600 170000 303000 170400
rect 303400 170000 303800 170400
rect 86000 169200 86400 169600
rect 86800 169200 87200 169600
rect 87600 169200 88000 169600
rect 88400 169200 88800 169600
rect 89200 169200 89600 169600
rect 90000 169200 90400 169600
rect 299400 169200 299800 169600
rect 300200 169200 300600 169600
rect 301000 169200 301400 169600
rect 301800 169200 302200 169600
rect 302600 169200 303000 169600
rect 303400 169200 303800 169600
rect 86000 168400 86400 168800
rect 86800 168400 87200 168800
rect 87600 168400 88000 168800
rect 88400 168400 88800 168800
rect 89200 168400 89600 168800
rect 90000 168400 90400 168800
rect 299400 168400 299800 168800
rect 300200 168400 300600 168800
rect 301000 168400 301400 168800
rect 301800 168400 302200 168800
rect 302600 168400 303000 168800
rect 303400 168400 303800 168800
rect 86000 167600 86400 168000
rect 86800 167600 87200 168000
rect 87600 167600 88000 168000
rect 88400 167600 88800 168000
rect 89200 167600 89600 168000
rect 90000 167600 90400 168000
rect 299400 167600 299800 168000
rect 300200 167600 300600 168000
rect 301000 167600 301400 168000
rect 301800 167600 302200 168000
rect 302600 167600 303000 168000
rect 303400 167600 303800 168000
rect 86000 166800 86400 167200
rect 86800 166800 87200 167200
rect 87600 166800 88000 167200
rect 88400 166800 88800 167200
rect 89200 166800 89600 167200
rect 90000 166800 90400 167200
rect 299400 166800 299800 167200
rect 300200 166800 300600 167200
rect 301000 166800 301400 167200
rect 301800 166800 302200 167200
rect 302600 166800 303000 167200
rect 303400 166800 303800 167200
rect 86000 166000 86400 166400
rect 86800 166000 87200 166400
rect 87600 166000 88000 166400
rect 88400 166000 88800 166400
rect 89200 166000 89600 166400
rect 90000 166000 90400 166400
rect 299400 166000 299800 166400
rect 300200 166000 300600 166400
rect 301000 166000 301400 166400
rect 301800 166000 302200 166400
rect 302600 166000 303000 166400
rect 303400 166000 303800 166400
rect 86000 165200 86400 165600
rect 86800 165200 87200 165600
rect 87600 165200 88000 165600
rect 88400 165200 88800 165600
rect 89200 165200 89600 165600
rect 90000 165200 90400 165600
rect 299400 165200 299800 165600
rect 300200 165200 300600 165600
rect 301000 165200 301400 165600
rect 301800 165200 302200 165600
rect 302600 165200 303000 165600
rect 303400 165200 303800 165600
rect 86000 164400 86400 164800
rect 86800 164400 87200 164800
rect 87600 164400 88000 164800
rect 88400 164400 88800 164800
rect 89200 164400 89600 164800
rect 90000 164400 90400 164800
rect 299400 164400 299800 164800
rect 300200 164400 300600 164800
rect 301000 164400 301400 164800
rect 301800 164400 302200 164800
rect 302600 164400 303000 164800
rect 303400 164400 303800 164800
rect 86000 163600 86400 164000
rect 86800 163600 87200 164000
rect 87600 163600 88000 164000
rect 88400 163600 88800 164000
rect 89200 163600 89600 164000
rect 90000 163600 90400 164000
rect 299400 163600 299800 164000
rect 300200 163600 300600 164000
rect 301000 163600 301400 164000
rect 301800 163600 302200 164000
rect 302600 163600 303000 164000
rect 303400 163600 303800 164000
rect 511700 301200 511900 301400
rect 512100 301200 512300 301400
rect 512500 301200 512700 301400
rect 512900 301200 513100 301400
rect 513300 301200 513500 301400
rect 513700 301200 513900 301400
rect 514100 301200 514300 301400
rect 514500 301200 514700 301400
rect 514900 301200 515100 301400
rect 515300 301200 515500 301400
rect 515700 301200 515900 301400
rect 516100 301200 516300 301400
rect 516500 301200 516700 301400
rect 511700 300800 511900 301000
rect 512100 300800 512300 301000
rect 512500 300800 512700 301000
rect 512900 300800 513100 301000
rect 513300 300800 513500 301000
rect 513700 300800 513900 301000
rect 514100 300800 514300 301000
rect 514500 300800 514700 301000
rect 514900 300800 515100 301000
rect 515300 300800 515500 301000
rect 515700 300800 515900 301000
rect 516100 300800 516300 301000
rect 516500 300800 516700 301000
rect 511700 300400 511900 300600
rect 512100 300400 512300 300600
rect 512500 300400 512700 300600
rect 512900 300400 513100 300600
rect 513300 300400 513500 300600
rect 513700 300400 513900 300600
rect 514100 300400 514300 300600
rect 514500 300400 514700 300600
rect 514900 300400 515100 300600
rect 515300 300400 515500 300600
rect 515700 300400 515900 300600
rect 516100 300400 516300 300600
rect 516500 300400 516700 300600
rect 530639 298862 530739 298992
rect 530899 298862 530999 298992
rect 528300 294200 528500 294400
rect 528700 294200 528900 294400
rect 529100 294200 529300 294400
rect 529500 294200 529700 294400
rect 529900 294200 530100 294400
rect 528300 293900 528500 294100
rect 528700 293900 528900 294100
rect 529100 293900 529300 294100
rect 529500 293900 529700 294100
rect 529900 293900 530100 294100
rect 528300 293500 528500 293700
rect 528700 293500 528900 293700
rect 529100 293500 529300 293700
rect 529500 293500 529700 293700
rect 529900 293500 530100 293700
rect 528300 293100 528500 293300
rect 528700 293100 528900 293300
rect 529100 293100 529300 293300
rect 529500 293100 529700 293300
rect 529900 293100 530100 293300
rect 528300 292700 528500 292900
rect 528700 292700 528900 292900
rect 529100 292700 529300 292900
rect 529500 292700 529700 292900
rect 529900 292700 530100 292900
rect 533197 298857 536541 298921
rect 536997 298857 540341 298921
rect 540797 298857 544141 298921
rect 544597 298857 547941 298921
rect 550129 298862 550239 298992
rect 550389 298862 550499 298992
rect 537089 294602 537169 294682
rect 537239 294602 537319 294682
rect 539579 294602 539659 294682
rect 539729 294602 539809 294682
rect 542059 294602 542139 294682
rect 542209 294602 542289 294682
rect 537089 294062 537169 294142
rect 537239 294062 537319 294142
rect 539579 294062 539659 294142
rect 539729 294062 539809 294142
rect 542059 294062 542139 294142
rect 542209 294062 542289 294142
rect 537089 293522 537169 293602
rect 537239 293522 537319 293602
rect 539579 293522 539659 293602
rect 539729 293522 539809 293602
rect 542069 293522 542149 293602
rect 542209 293522 542289 293602
rect 538379 292922 538459 293002
rect 538489 292922 538569 293002
rect 540789 292922 540869 293002
rect 540899 292922 540979 293002
rect 543249 292912 543329 292992
rect 543359 292912 543439 292992
rect 538379 292312 538459 292392
rect 538489 292312 538569 292392
rect 540789 292332 540869 292412
rect 540899 292332 540979 292412
rect 543249 292332 543329 292412
rect 543359 292332 543439 292412
rect 569300 301955 569500 302000
rect 569800 301955 570000 302000
rect 569300 301895 569330 301955
rect 569330 301895 569390 301955
rect 569390 301895 569500 301955
rect 569800 301895 569920 301955
rect 569920 301895 569980 301955
rect 569980 301895 570000 301955
rect 569300 301800 569500 301895
rect 569800 301800 570000 301895
rect 569300 301565 569500 301600
rect 569800 301565 570000 301600
rect 569300 301505 569330 301565
rect 569330 301505 569390 301565
rect 569390 301505 569500 301565
rect 569800 301505 569920 301565
rect 569920 301505 569980 301565
rect 569980 301505 570000 301565
rect 569300 301400 569500 301505
rect 569800 301400 570000 301505
rect 569300 301185 569500 301200
rect 569800 301185 570000 301200
rect 569300 301125 569330 301185
rect 569330 301125 569390 301185
rect 569390 301125 569500 301185
rect 569800 301125 569920 301185
rect 569920 301125 569980 301185
rect 569980 301125 570000 301185
rect 569300 301000 569500 301125
rect 569800 301000 570000 301125
rect 569300 300775 569330 300800
rect 569330 300775 569390 300800
rect 569390 300775 569500 300800
rect 569800 300775 569920 300800
rect 569920 300775 569980 300800
rect 569980 300775 570000 300800
rect 569300 300645 569500 300775
rect 569800 300645 570000 300775
rect 569300 300600 569330 300645
rect 569330 300600 569390 300645
rect 569390 300600 569500 300645
rect 569800 300600 569920 300645
rect 569920 300600 569980 300645
rect 569980 300600 570000 300645
rect 569300 300330 569500 300400
rect 569800 300330 570000 300400
rect 569300 300270 569330 300330
rect 569330 300270 569390 300330
rect 569390 300270 569500 300330
rect 569800 300270 569920 300330
rect 569920 300270 569980 300330
rect 569980 300270 570000 300330
rect 569300 300200 569500 300270
rect 569800 300200 570000 300270
rect 538379 291752 538459 291832
rect 538489 291752 538569 291832
rect 540789 291752 540869 291832
rect 540899 291752 540979 291832
rect 543249 291752 543329 291832
rect 543359 291752 543439 291832
rect 534869 291542 534959 291652
rect 535029 291542 535119 291652
rect 544799 291522 544879 291602
rect 544969 291522 545049 291602
rect 545900 291142 546100 291200
rect 546200 291142 546400 291200
rect 545900 291062 546069 291142
rect 546069 291062 546100 291142
rect 546200 291062 546229 291142
rect 546229 291062 546319 291142
rect 546319 291062 546400 291142
rect 545900 291000 546100 291062
rect 546200 291000 546400 291062
rect 546500 291000 546700 291200
rect 546800 291000 547000 291200
rect 547200 291100 547400 291300
rect 547200 290800 547400 291000
rect 547200 290500 547400 290700
rect 547200 290200 547400 290400
rect 545800 289900 546000 290100
rect 546100 290062 546300 290100
rect 546100 289982 546159 290062
rect 546159 289982 546229 290062
rect 546229 289982 546300 290062
rect 546100 289900 546300 289982
rect 546400 289900 546600 290100
rect 546800 289900 547000 290100
rect 538379 289052 538459 289132
rect 538489 289052 538569 289132
rect 540789 289052 540869 289132
rect 540899 289052 540979 289132
rect 543249 289062 543329 289142
rect 543359 289062 543439 289142
rect 511700 288600 511900 288800
rect 512100 288600 512300 288800
rect 512500 288600 512700 288800
rect 512900 288600 513100 288800
rect 513300 288600 513500 288800
rect 513700 288600 513900 288800
rect 514100 288600 514300 288800
rect 514500 288600 514700 288800
rect 514900 288600 515100 288800
rect 515300 288600 515500 288800
rect 515700 288600 515900 288800
rect 516100 288600 516300 288800
rect 516500 288600 516700 288800
rect 572800 288564 573100 288700
rect 573300 288564 573600 288700
rect 573800 288564 574100 288700
rect 574300 288694 574540 288700
rect 574540 288694 574600 288700
rect 574300 288564 574600 288694
rect 511700 288200 511900 288400
rect 512100 288200 512300 288400
rect 512500 288200 512700 288400
rect 512900 288200 513100 288400
rect 513300 288200 513500 288400
rect 513700 288200 513900 288400
rect 514100 288200 514300 288400
rect 514500 288200 514700 288400
rect 514900 288200 515100 288400
rect 515300 288200 515500 288400
rect 515700 288200 515900 288400
rect 516100 288200 516300 288400
rect 516500 288200 516700 288400
rect 537089 288292 537169 288372
rect 537239 288292 537319 288372
rect 539579 288312 539659 288392
rect 539729 288312 539809 288392
rect 542059 288312 542139 288392
rect 542199 288312 542279 288392
rect 511700 287800 511900 288000
rect 512100 287800 512300 288000
rect 512500 287800 512700 288000
rect 512900 287800 513100 288000
rect 513300 287800 513500 288000
rect 513700 287800 513900 288000
rect 514100 287800 514300 288000
rect 514500 287800 514700 288000
rect 514900 287800 515100 288000
rect 515300 287800 515500 288000
rect 515700 287800 515900 288000
rect 516100 287800 516300 288000
rect 516500 287800 516700 288000
rect 511700 287400 511900 287600
rect 512100 287400 512300 287600
rect 512500 287400 512700 287600
rect 512900 287400 513100 287600
rect 513300 287400 513500 287600
rect 513700 287400 513900 287600
rect 514100 287400 514300 287600
rect 514500 287400 514700 287600
rect 514900 287400 515100 287600
rect 515300 287400 515500 287600
rect 515700 287400 515900 287600
rect 516100 287400 516300 287600
rect 516500 287400 516700 287600
rect 572800 288504 572810 288564
rect 572810 288504 572890 288564
rect 572890 288504 572950 288564
rect 572950 288504 573065 288564
rect 573065 288504 573100 288564
rect 573300 288504 573315 288564
rect 573315 288504 573415 288564
rect 573415 288504 573475 288564
rect 573475 288504 573600 288564
rect 573800 288504 573805 288564
rect 573805 288504 573865 288564
rect 573865 288504 573985 288564
rect 573985 288504 574045 288564
rect 574045 288504 574100 288564
rect 574300 288504 574375 288564
rect 574375 288504 574435 288564
rect 574435 288504 574540 288564
rect 574540 288504 574600 288564
rect 572800 288400 573100 288504
rect 573300 288400 573600 288504
rect 573800 288400 574100 288504
rect 574300 288400 574600 288504
rect 572800 288174 573100 288200
rect 573300 288174 573600 288200
rect 573800 288174 574100 288200
rect 574300 288174 574600 288200
rect 572800 288114 572810 288174
rect 572810 288114 572890 288174
rect 572890 288114 572950 288174
rect 572950 288114 573065 288174
rect 573065 288114 573100 288174
rect 573300 288114 573315 288174
rect 573315 288114 573415 288174
rect 573415 288114 573475 288174
rect 573475 288114 573600 288174
rect 573800 288114 573805 288174
rect 573805 288114 573865 288174
rect 573865 288114 573985 288174
rect 573985 288114 574045 288174
rect 574045 288114 574100 288174
rect 574300 288114 574375 288174
rect 574375 288114 574435 288174
rect 574435 288114 574540 288174
rect 574540 288114 574600 288174
rect 572800 287974 573100 288114
rect 573300 287974 573600 288114
rect 573800 287974 574100 288114
rect 574300 287974 574600 288114
rect 572800 287914 572810 287974
rect 572810 287914 572890 287974
rect 572890 287914 572950 287974
rect 572950 287914 573065 287974
rect 573065 287914 573100 287974
rect 573300 287914 573315 287974
rect 573315 287914 573415 287974
rect 573415 287914 573475 287974
rect 573475 287914 573600 287974
rect 573800 287914 573805 287974
rect 573805 287914 573865 287974
rect 573865 287914 573985 287974
rect 573985 287914 574045 287974
rect 574045 287914 574100 287974
rect 574300 287914 574375 287974
rect 574375 287914 574435 287974
rect 574435 287914 574540 287974
rect 574540 287914 574600 287974
rect 572800 287900 573100 287914
rect 573300 287900 573600 287914
rect 573800 287900 574100 287914
rect 574300 287900 574600 287914
rect 511700 287000 511900 287200
rect 512100 287000 512300 287200
rect 512500 287000 512700 287200
rect 512900 287000 513100 287200
rect 513300 287000 513500 287200
rect 513700 287000 513900 287200
rect 514100 287000 514300 287200
rect 514500 287000 514700 287200
rect 514900 287000 515100 287200
rect 515300 287000 515500 287200
rect 515700 287000 515900 287200
rect 516100 287000 516300 287200
rect 516500 287000 516700 287200
rect 511700 286600 511900 286800
rect 512100 286600 512300 286800
rect 512500 286600 512700 286800
rect 512900 286600 513100 286800
rect 513300 286600 513500 286800
rect 513700 286600 513900 286800
rect 514100 286600 514300 286800
rect 514500 286600 514700 286800
rect 514900 286600 515100 286800
rect 515300 286600 515500 286800
rect 515700 286600 515900 286800
rect 516100 286600 516300 286800
rect 516500 286600 516700 286800
rect 542389 286342 542509 286442
rect 545800 285200 546000 285400
rect 546200 285200 546400 285400
rect 546600 285200 546800 285400
rect 547000 285200 547200 285400
rect 547400 285200 547600 285400
rect 547800 285200 548000 285400
rect 548200 285200 548400 285400
rect 548600 285200 548800 285400
rect 545800 284800 546000 285000
rect 546200 284800 546400 285000
rect 546600 284800 546800 285000
rect 547000 284800 547200 285000
rect 547400 284800 547600 285000
rect 547800 284800 548000 285000
rect 548200 284800 548400 285000
rect 548600 284800 548800 285000
rect 511900 283000 512100 283200
rect 512300 283000 512500 283200
rect 512700 283000 512900 283200
rect 513100 283000 513300 283200
rect 513500 283000 513700 283200
rect 513900 283000 514100 283200
rect 514300 283000 514500 283200
rect 514700 283000 514900 283200
rect 515100 283000 515300 283200
rect 515500 283000 515700 283200
rect 515900 283000 516100 283200
rect 516300 283000 516500 283200
rect 516700 283000 516900 283200
rect 511900 282600 512100 282800
rect 512300 282600 512500 282800
rect 512700 282600 512900 282800
rect 513100 282600 513300 282800
rect 513500 282600 513700 282800
rect 513900 282600 514100 282800
rect 514300 282600 514500 282800
rect 514700 282600 514900 282800
rect 515100 282600 515300 282800
rect 515500 282600 515700 282800
rect 515900 282600 516100 282800
rect 516300 282600 516500 282800
rect 516700 282600 516900 282800
rect 511900 282200 512100 282400
rect 512300 282200 512500 282400
rect 512700 282200 512900 282400
rect 513100 282200 513300 282400
rect 513500 282200 513700 282400
rect 513900 282200 514100 282400
rect 514300 282200 514500 282400
rect 514700 282200 514900 282400
rect 515100 282200 515300 282400
rect 515500 282200 515700 282400
rect 515900 282200 516100 282400
rect 516300 282200 516500 282400
rect 516700 282200 516900 282400
rect 511900 281800 512100 282000
rect 512300 281800 512500 282000
rect 512700 281800 512900 282000
rect 513100 281800 513300 282000
rect 513500 281800 513700 282000
rect 513900 281800 514100 282000
rect 514300 281800 514500 282000
rect 514700 281800 514900 282000
rect 515100 281800 515300 282000
rect 515500 281800 515700 282000
rect 515900 281800 516100 282000
rect 516300 281800 516500 282000
rect 516700 281800 516900 282000
rect 511900 281400 512100 281600
rect 512300 281400 512500 281600
rect 512700 281400 512900 281600
rect 513100 281400 513300 281600
rect 513500 281400 513700 281600
rect 513900 281400 514100 281600
rect 514300 281400 514500 281600
rect 514700 281400 514900 281600
rect 515100 281400 515300 281600
rect 515500 281400 515700 281600
rect 515900 281400 516100 281600
rect 516300 281400 516500 281600
rect 516700 281400 516900 281600
rect 511900 281000 512100 281200
rect 512300 281000 512500 281200
rect 512700 281000 512900 281200
rect 513100 281000 513300 281200
rect 513500 281000 513700 281200
rect 513900 281000 514100 281200
rect 514300 281000 514500 281200
rect 514700 281000 514900 281200
rect 515100 281000 515300 281200
rect 515500 281000 515700 281200
rect 515900 281000 516100 281200
rect 516300 281000 516500 281200
rect 516700 281000 516900 281200
rect 511900 280600 512100 280800
rect 512300 280600 512500 280800
rect 512700 280600 512900 280800
rect 513100 280600 513300 280800
rect 513500 280600 513700 280800
rect 513900 280600 514100 280800
rect 514300 280600 514500 280800
rect 514700 280600 514900 280800
rect 515100 280600 515300 280800
rect 515500 280600 515700 280800
rect 515900 280600 516100 280800
rect 516300 280600 516500 280800
rect 516700 280600 516900 280800
rect 546000 248400 546200 248600
rect 546400 248400 546600 248600
rect 546800 248400 547000 248600
rect 547200 248400 547400 248600
rect 547600 248400 547800 248600
rect 548000 248400 548200 248600
rect 548400 248400 548600 248600
rect 548800 248400 549000 248600
rect 546000 248000 546200 248200
rect 546400 248000 546600 248200
rect 546800 248000 547000 248200
rect 547200 248000 547400 248200
rect 547600 248000 547800 248200
rect 548000 248000 548200 248200
rect 548400 248000 548600 248200
rect 548800 248000 549000 248200
rect 546000 247600 546200 247800
rect 546400 247600 546600 247800
rect 546800 247600 547000 247800
rect 547200 247600 547400 247800
rect 547600 247600 547800 247800
rect 548000 247600 548200 247800
rect 548400 247600 548600 247800
rect 548800 247600 549000 247800
rect 546000 247200 546200 247400
rect 546400 247200 546600 247400
rect 546800 247200 547000 247400
rect 547200 247200 547400 247400
rect 547600 247200 547800 247400
rect 548000 247200 548200 247400
rect 548400 247200 548600 247400
rect 548800 247200 549000 247400
rect 546000 246800 546200 247000
rect 546400 246800 546600 247000
rect 546800 246800 547000 247000
rect 547200 246800 547400 247000
rect 547600 246800 547800 247000
rect 548000 246800 548200 247000
rect 548400 246800 548600 247000
rect 548800 246800 549000 247000
rect 546000 246400 546200 246600
rect 546400 246400 546600 246600
rect 546800 246400 547000 246600
rect 547200 246400 547400 246600
rect 547600 246400 547800 246600
rect 548000 246400 548200 246600
rect 548400 246400 548600 246600
rect 548800 246400 549000 246600
rect 546000 246000 546200 246200
rect 546400 246000 546600 246200
rect 546800 246000 547000 246200
rect 547200 246000 547400 246200
rect 547600 246000 547800 246200
rect 548000 246000 548200 246200
rect 548400 246000 548600 246200
rect 548800 246000 549000 246200
rect 546000 245600 546200 245800
rect 546400 245600 546600 245800
rect 546800 245600 547000 245800
rect 547200 245600 547400 245800
rect 547600 245600 547800 245800
rect 548000 245600 548200 245800
rect 548400 245600 548600 245800
rect 548800 245600 549000 245800
rect 546000 245200 546200 245400
rect 546400 245200 546600 245400
rect 546800 245200 547000 245400
rect 547200 245200 547400 245400
rect 547600 245200 547800 245400
rect 548000 245200 548200 245400
rect 548400 245200 548600 245400
rect 548800 245200 549000 245400
rect 546000 244800 546200 245000
rect 546400 244800 546600 245000
rect 546800 244800 547000 245000
rect 547200 244800 547400 245000
rect 547600 244800 547800 245000
rect 548000 244800 548200 245000
rect 548400 244800 548600 245000
rect 548800 244800 549000 245000
rect 546000 244400 546200 244600
rect 546400 244400 546600 244600
rect 546800 244400 547000 244600
rect 547200 244400 547400 244600
rect 547600 244400 547800 244600
rect 548000 244400 548200 244600
rect 548400 244400 548600 244600
rect 548800 244400 549000 244600
rect 546000 244000 546200 244200
rect 546400 244000 546600 244200
rect 546800 244000 547000 244200
rect 547200 244000 547400 244200
rect 547600 244000 547800 244200
rect 548000 244000 548200 244200
rect 548400 244000 548600 244200
rect 548800 244000 549000 244200
rect 546000 243600 546200 243800
rect 546400 243600 546600 243800
rect 546800 243600 547000 243800
rect 547200 243600 547400 243800
rect 547600 243600 547800 243800
rect 548000 243600 548200 243800
rect 548400 243600 548600 243800
rect 548800 243600 549000 243800
rect 546000 243200 546200 243400
rect 546400 243200 546600 243400
rect 546800 243200 547000 243400
rect 547200 243200 547400 243400
rect 547600 243200 547800 243400
rect 548000 243200 548200 243400
rect 548400 243200 548600 243400
rect 548800 243200 549000 243400
rect 546000 242800 546200 243000
rect 546400 242800 546600 243000
rect 546800 242800 547000 243000
rect 547200 242800 547400 243000
rect 547600 242800 547800 243000
rect 548000 242800 548200 243000
rect 548400 242800 548600 243000
rect 548800 242800 549000 243000
rect 546000 242400 546200 242600
rect 546400 242400 546600 242600
rect 546800 242400 547000 242600
rect 547200 242400 547400 242600
rect 547600 242400 547800 242600
rect 548000 242400 548200 242600
rect 548400 242400 548600 242600
rect 548800 242400 549000 242600
rect 546000 242000 546200 242200
rect 546400 242000 546600 242200
rect 546800 242000 547000 242200
rect 547200 242000 547400 242200
rect 547600 242000 547800 242200
rect 548000 242000 548200 242200
rect 548400 242000 548600 242200
rect 548800 242000 549000 242200
rect 546000 241600 546200 241800
rect 546400 241600 546600 241800
rect 546800 241600 547000 241800
rect 547200 241600 547400 241800
rect 547600 241600 547800 241800
rect 548000 241600 548200 241800
rect 548400 241600 548600 241800
rect 548800 241600 549000 241800
rect 546000 241200 546200 241400
rect 546400 241200 546600 241400
rect 546800 241200 547000 241400
rect 547200 241200 547400 241400
rect 547600 241200 547800 241400
rect 548000 241200 548200 241400
rect 548400 241200 548600 241400
rect 548800 241200 549000 241400
rect 546000 240800 546200 241000
rect 546400 240800 546600 241000
rect 546800 240800 547000 241000
rect 547200 240800 547400 241000
rect 547600 240800 547800 241000
rect 548000 240800 548200 241000
rect 548400 240800 548600 241000
rect 548800 240800 549000 241000
rect 546000 240400 546200 240600
rect 546400 240400 546600 240600
rect 546800 240400 547000 240600
rect 547200 240400 547400 240600
rect 547600 240400 547800 240600
rect 548000 240400 548200 240600
rect 548400 240400 548600 240600
rect 548800 240400 549000 240600
rect 546000 240000 546200 240200
rect 546400 240000 546600 240200
rect 546800 240000 547000 240200
rect 547200 240000 547400 240200
rect 547600 240000 547800 240200
rect 548000 240000 548200 240200
rect 548400 240000 548600 240200
rect 548800 240000 549000 240200
rect 546000 239600 546200 239800
rect 546400 239600 546600 239800
rect 546800 239600 547000 239800
rect 547200 239600 547400 239800
rect 547600 239600 547800 239800
rect 548000 239600 548200 239800
rect 548400 239600 548600 239800
rect 548800 239600 549000 239800
rect 546000 239200 546200 239400
rect 546400 239200 546600 239400
rect 546800 239200 547000 239400
rect 547200 239200 547400 239400
rect 547600 239200 547800 239400
rect 548000 239200 548200 239400
rect 548400 239200 548600 239400
rect 548800 239200 549000 239400
rect 546000 238800 546200 239000
rect 546400 238800 546600 239000
rect 546800 238800 547000 239000
rect 547200 238800 547400 239000
rect 547600 238800 547800 239000
rect 548000 238800 548200 239000
rect 548400 238800 548600 239000
rect 548800 238800 549000 239000
rect 546000 238400 546200 238600
rect 546400 238400 546600 238600
rect 546800 238400 547000 238600
rect 547200 238400 547400 238600
rect 547600 238400 547800 238600
rect 548000 238400 548200 238600
rect 548400 238400 548600 238600
rect 548800 238400 549000 238600
rect 546000 238000 546200 238200
rect 546400 238000 546600 238200
rect 546800 238000 547000 238200
rect 547200 238000 547400 238200
rect 547600 238000 547800 238200
rect 548000 238000 548200 238200
rect 548400 238000 548600 238200
rect 548800 238000 549000 238200
rect 546000 237600 546200 237800
rect 546400 237600 546600 237800
rect 546800 237600 547000 237800
rect 547200 237600 547400 237800
rect 547600 237600 547800 237800
rect 548000 237600 548200 237800
rect 548400 237600 548600 237800
rect 548800 237600 549000 237800
rect 546000 237200 546200 237400
rect 546400 237200 546600 237400
rect 546800 237200 547000 237400
rect 547200 237200 547400 237400
rect 547600 237200 547800 237400
rect 548000 237200 548200 237400
rect 548400 237200 548600 237400
rect 548800 237200 549000 237400
rect 546000 236800 546200 237000
rect 546400 236800 546600 237000
rect 546800 236800 547000 237000
rect 547200 236800 547400 237000
rect 547600 236800 547800 237000
rect 548000 236800 548200 237000
rect 548400 236800 548600 237000
rect 548800 236800 549000 237000
rect 546000 236400 546200 236600
rect 546400 236400 546600 236600
rect 546800 236400 547000 236600
rect 547200 236400 547400 236600
rect 547600 236400 547800 236600
rect 548000 236400 548200 236600
rect 548400 236400 548600 236600
rect 548800 236400 549000 236600
rect 546000 236000 546200 236200
rect 546400 236000 546600 236200
rect 546800 236000 547000 236200
rect 547200 236000 547400 236200
rect 547600 236000 547800 236200
rect 548000 236000 548200 236200
rect 548400 236000 548600 236200
rect 548800 236000 549000 236200
rect 546000 235600 546200 235800
rect 546400 235600 546600 235800
rect 546800 235600 547000 235800
rect 547200 235600 547400 235800
rect 547600 235600 547800 235800
rect 548000 235600 548200 235800
rect 548400 235600 548600 235800
rect 548800 235600 549000 235800
rect 546000 235200 546200 235400
rect 546400 235200 546600 235400
rect 546800 235200 547000 235400
rect 547200 235200 547400 235400
rect 547600 235200 547800 235400
rect 548000 235200 548200 235400
rect 548400 235200 548600 235400
rect 548800 235200 549000 235400
rect 546000 234800 546200 235000
rect 546400 234800 546600 235000
rect 546800 234800 547000 235000
rect 547200 234800 547400 235000
rect 547600 234800 547800 235000
rect 548000 234800 548200 235000
rect 548400 234800 548600 235000
rect 548800 234800 549000 235000
rect 546000 234500 546200 234700
rect 546400 234500 546600 234700
rect 546800 234500 547000 234700
rect 547200 234500 547400 234700
rect 547600 234500 547800 234700
rect 548000 234500 548200 234700
rect 548400 234500 548600 234700
rect 548800 234500 549000 234700
rect 546000 234200 546200 234400
rect 546400 234200 546600 234400
rect 546800 234200 547000 234400
rect 547200 234200 547400 234400
rect 547600 234200 547800 234400
rect 548000 234200 548200 234400
rect 548400 234200 548600 234400
rect 548800 234200 549000 234400
rect 546000 233800 546200 234000
rect 546400 233800 546600 234000
rect 546800 233800 547000 234000
rect 547200 233800 547400 234000
rect 547600 233800 547800 234000
rect 548000 233800 548200 234000
rect 548400 233800 548600 234000
rect 548800 233800 549000 234000
rect 512000 195200 512400 195600
rect 512800 195200 513200 195600
rect 513600 195200 514000 195600
rect 514400 195200 514800 195600
rect 515200 195200 515600 195600
rect 516000 195200 516400 195600
rect 512000 194400 512400 194800
rect 512800 194400 513200 194800
rect 513600 194400 514000 194800
rect 514400 194400 514800 194800
rect 515200 194400 515600 194800
rect 516000 194400 516400 194800
rect 512000 193600 512400 194000
rect 512800 193600 513200 194000
rect 513600 193600 514000 194000
rect 514400 193600 514800 194000
rect 515200 193600 515600 194000
rect 516000 193600 516400 194000
rect 512000 192800 512400 193200
rect 512800 192800 513200 193200
rect 513600 192800 514000 193200
rect 514400 192800 514800 193200
rect 515200 192800 515600 193200
rect 516000 192800 516400 193200
rect 512000 192000 512400 192400
rect 512800 192000 513200 192400
rect 513600 192000 514000 192400
rect 514400 192000 514800 192400
rect 515200 192000 515600 192400
rect 516000 192000 516400 192400
rect 512000 191200 512400 191600
rect 512800 191200 513200 191600
rect 513600 191200 514000 191600
rect 514400 191200 514800 191600
rect 515200 191200 515600 191600
rect 516000 191200 516400 191600
rect 512000 190400 512400 190800
rect 512800 190400 513200 190800
rect 513600 190400 514000 190800
rect 514400 190400 514800 190800
rect 515200 190400 515600 190800
rect 516000 190400 516400 190800
rect 512000 189600 512400 190000
rect 512800 189600 513200 190000
rect 513600 189600 514000 190000
rect 514400 189600 514800 190000
rect 515200 189600 515600 190000
rect 516000 189600 516400 190000
rect 512000 188800 512400 189200
rect 512800 188800 513200 189200
rect 513600 188800 514000 189200
rect 514400 188800 514800 189200
rect 515200 188800 515600 189200
rect 516000 188800 516400 189200
rect 512000 188000 512400 188400
rect 512800 188000 513200 188400
rect 513600 188000 514000 188400
rect 514400 188000 514800 188400
rect 515200 188000 515600 188400
rect 516000 188000 516400 188400
rect 512000 187200 512400 187600
rect 512800 187200 513200 187600
rect 513600 187200 514000 187600
rect 514400 187200 514800 187600
rect 515200 187200 515600 187600
rect 516000 187200 516400 187600
rect 512000 186400 512400 186800
rect 512800 186400 513200 186800
rect 513600 186400 514000 186800
rect 514400 186400 514800 186800
rect 515200 186400 515600 186800
rect 516000 186400 516400 186800
rect 512000 185600 512400 186000
rect 512800 185600 513200 186000
rect 513600 185600 514000 186000
rect 514400 185600 514800 186000
rect 515200 185600 515600 186000
rect 516000 185600 516400 186000
rect 512000 184800 512400 185200
rect 512800 184800 513200 185200
rect 513600 184800 514000 185200
rect 514400 184800 514800 185200
rect 515200 184800 515600 185200
rect 516000 184800 516400 185200
rect 512000 184000 512400 184400
rect 512800 184000 513200 184400
rect 513600 184000 514000 184400
rect 514400 184000 514800 184400
rect 515200 184000 515600 184400
rect 516000 184000 516400 184400
rect 512000 183200 512400 183600
rect 512800 183200 513200 183600
rect 513600 183200 514000 183600
rect 514400 183200 514800 183600
rect 515200 183200 515600 183600
rect 516000 183200 516400 183600
rect 512000 182400 512400 182800
rect 512800 182400 513200 182800
rect 513600 182400 514000 182800
rect 514400 182400 514800 182800
rect 515200 182400 515600 182800
rect 516000 182400 516400 182800
rect 512000 181600 512400 182000
rect 512800 181600 513200 182000
rect 513600 181600 514000 182000
rect 514400 181600 514800 182000
rect 515200 181600 515600 182000
rect 516000 181600 516400 182000
<< mimcap >>
rect 533269 298702 536469 298742
rect 533269 295582 533309 298702
rect 536429 295582 536469 298702
rect 533269 295542 536469 295582
rect 537069 298702 540269 298742
rect 537069 295582 537109 298702
rect 540229 295582 540269 298702
rect 537069 295542 540269 295582
rect 540869 298702 544069 298742
rect 540869 295582 540909 298702
rect 544029 295582 544069 298702
rect 540869 295542 544069 295582
rect 544669 298702 547869 298742
rect 544669 295582 544709 298702
rect 547829 295582 547869 298702
rect 544669 295542 547869 295582
rect 7070 279910 10270 279950
rect 7070 276790 7110 279910
rect 10230 276790 10270 279910
rect 7070 276750 10270 276790
rect 7070 276110 10270 276150
rect 7070 272990 7110 276110
rect 10230 272990 10270 276110
rect 7070 272950 10270 272990
rect 7070 272310 10270 272350
rect 7070 269190 7110 272310
rect 10230 269190 10270 272310
rect 7070 269150 10270 269190
rect 7070 268510 10270 268550
rect 7070 265390 7110 268510
rect 10230 265390 10270 268510
rect 7070 265350 10270 265390
<< mimcapcontact >>
rect 533309 295582 536429 298702
rect 537109 295582 540229 298702
rect 540909 295582 544029 298702
rect 544709 295582 547829 298702
rect 7110 276790 10230 279910
rect 7110 272990 10230 276110
rect 7110 269190 10230 272310
rect 7110 265390 10230 268510
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 16200 702200 24340 702300
rect 16200 702000 16400 702200
rect 16600 702000 16800 702200
rect 17000 702000 17200 702200
rect 17400 702000 17600 702200
rect 17800 702000 18000 702200
rect 18200 702000 18400 702200
rect 18600 702000 18800 702200
rect 19000 702000 19200 702200
rect 19400 702000 19600 702200
rect 19800 702000 20000 702200
rect 20200 702000 20400 702200
rect 20600 702000 20800 702200
rect 21000 702180 24340 702200
rect 21000 702060 23400 702180
rect 23520 702060 23600 702180
rect 23720 702060 23800 702180
rect 23920 702060 24000 702180
rect 24120 702060 24200 702180
rect 24320 702060 24340 702180
rect 21000 702000 24340 702060
rect 65040 702260 73200 702300
rect 65040 702080 65060 702260
rect 65240 702080 65400 702260
rect 65580 702080 65740 702260
rect 65920 702200 73200 702260
rect 65920 702080 68400 702200
rect 65040 702040 68400 702080
rect 16200 701940 24340 702000
rect 68200 702000 68400 702040
rect 68600 702000 68800 702200
rect 69000 702000 69200 702200
rect 69400 702000 69600 702200
rect 69800 702000 70000 702200
rect 70200 702000 70400 702200
rect 70600 702000 70800 702200
rect 71000 702000 71200 702200
rect 71400 702000 71600 702200
rect 71800 702000 72000 702200
rect 72200 702000 72400 702200
rect 72600 702000 72800 702200
rect 73000 702000 73200 702200
rect 16200 701800 21200 701940
rect 16200 701600 16400 701800
rect 16600 701600 16800 701800
rect 17000 701600 17200 701800
rect 17400 701600 17600 701800
rect 17800 701600 18000 701800
rect 18200 701600 18400 701800
rect 18600 701600 18800 701800
rect 19000 701600 19200 701800
rect 19400 701600 19600 701800
rect 19800 701600 20000 701800
rect 20200 701600 20400 701800
rect 20600 701600 20800 701800
rect 21000 701600 21200 701800
rect 16200 701400 21200 701600
rect 16200 701200 16400 701400
rect 16600 701200 16800 701400
rect 17000 701200 17200 701400
rect 17400 701200 17600 701400
rect 17800 701200 18000 701400
rect 18200 701200 18400 701400
rect 18600 701200 18800 701400
rect 19000 701200 19200 701400
rect 19400 701200 19600 701400
rect 19800 701200 20000 701400
rect 20200 701200 20400 701400
rect 20600 701200 20800 701400
rect 21000 701200 21200 701400
rect 16200 701000 21200 701200
rect 16200 700800 16400 701000
rect 16600 700800 16800 701000
rect 17000 700800 17200 701000
rect 17400 700800 17600 701000
rect 17800 700800 18000 701000
rect 18200 700800 18400 701000
rect 18600 700800 18800 701000
rect 19000 700800 19200 701000
rect 19400 700800 19600 701000
rect 19800 700800 20000 701000
rect 20200 700800 20400 701000
rect 20600 700800 20800 701000
rect 21000 700800 21200 701000
rect 16200 700600 21200 700800
rect 16200 700400 16400 700600
rect 16600 700400 16800 700600
rect 17000 700400 17200 700600
rect 17400 700400 17600 700600
rect 17800 700400 18000 700600
rect 18200 700400 18400 700600
rect 18600 700400 18800 700600
rect 19000 700400 19200 700600
rect 19400 700400 19600 700600
rect 19800 700400 20000 700600
rect 20200 700400 20400 700600
rect 20600 700400 20800 700600
rect 21000 700400 21200 700600
rect 16200 700200 21200 700400
rect 16200 700000 16400 700200
rect 16600 700000 16800 700200
rect 17000 700000 17200 700200
rect 17400 700000 17600 700200
rect 17800 700000 18000 700200
rect 18200 700000 18400 700200
rect 18600 700000 18800 700200
rect 19000 700000 19200 700200
rect 19400 700000 19600 700200
rect 19800 700000 20000 700200
rect 20200 700000 20400 700200
rect 20600 700000 20800 700200
rect 21000 700000 21200 700200
rect 16200 698400 21200 700000
rect 68200 701800 73200 702000
rect 68200 701600 68400 701800
rect 68600 701600 68800 701800
rect 69000 701600 69200 701800
rect 69400 701600 69600 701800
rect 69800 701600 70000 701800
rect 70200 701600 70400 701800
rect 70600 701600 70800 701800
rect 71000 701600 71200 701800
rect 71400 701600 71600 701800
rect 71800 701600 72000 701800
rect 72200 701600 72400 701800
rect 72600 701600 72800 701800
rect 73000 701600 73200 701800
rect 68200 701400 73200 701600
rect 68200 701200 68400 701400
rect 68600 701200 68800 701400
rect 69000 701200 69200 701400
rect 69400 701200 69600 701400
rect 69800 701200 70000 701400
rect 70200 701200 70400 701400
rect 70600 701200 70800 701400
rect 71000 701200 71200 701400
rect 71400 701200 71600 701400
rect 71800 701200 72000 701400
rect 72200 701200 72400 701400
rect 72600 701200 72800 701400
rect 73000 701200 73200 701400
rect 68200 701000 73200 701200
rect 68200 700800 68400 701000
rect 68600 700800 68800 701000
rect 69000 700800 69200 701000
rect 69400 700800 69600 701000
rect 69800 700800 70000 701000
rect 70200 700800 70400 701000
rect 70600 700800 70800 701000
rect 71000 700800 71200 701000
rect 71400 700800 71600 701000
rect 71800 700800 72000 701000
rect 72200 700800 72400 701000
rect 72600 700800 72800 701000
rect 73000 700800 73200 701000
rect 68200 700600 73200 700800
rect 68200 700400 68400 700600
rect 68600 700400 68800 700600
rect 69000 700400 69200 700600
rect 69400 700400 69600 700600
rect 69800 700400 70000 700600
rect 70200 700400 70400 700600
rect 70600 700400 70800 700600
rect 71000 700400 71200 700600
rect 71400 700400 71600 700600
rect 71800 700400 72000 700600
rect 72200 700400 72400 700600
rect 72600 700400 72800 700600
rect 73000 700400 73200 700600
rect 68200 700200 73200 700400
rect 68200 700000 68400 700200
rect 68600 700000 68800 700200
rect 69000 700000 69200 700200
rect 69400 700000 69600 700200
rect 69800 700000 70000 700200
rect 70200 700000 70400 700200
rect 70600 700000 70800 700200
rect 71000 700000 71200 700200
rect 71400 700000 71600 700200
rect 71800 700000 72000 700200
rect 72200 700000 72400 700200
rect 72600 700000 72800 700200
rect 73000 700000 73200 700200
rect 68200 698400 73200 700000
rect 515500 701600 521000 701800
rect 515500 701400 515700 701600
rect 515900 701400 516100 701600
rect 516300 701400 516500 701600
rect 516700 701400 516900 701600
rect 517100 701400 517300 701600
rect 517500 701400 517700 701600
rect 517900 701400 518100 701600
rect 518300 701400 518500 701600
rect 518700 701400 518900 701600
rect 519100 701400 519300 701600
rect 519500 701400 519700 701600
rect 519900 701400 520100 701600
rect 520300 701400 520500 701600
rect 520700 701400 521000 701600
rect 515500 701200 521000 701400
rect 515500 701000 515700 701200
rect 515900 701000 516100 701200
rect 516300 701000 516500 701200
rect 516700 701000 516900 701200
rect 517100 701000 517300 701200
rect 517500 701000 517700 701200
rect 517900 701000 518100 701200
rect 518300 701000 518500 701200
rect 518700 701000 518900 701200
rect 519100 701000 519300 701200
rect 519500 701000 519700 701200
rect 519900 701000 520100 701200
rect 520300 701000 520500 701200
rect 520700 701000 521000 701200
rect 515500 700800 521000 701000
rect 515500 700600 515700 700800
rect 515900 700600 516100 700800
rect 516300 700600 516500 700800
rect 516700 700600 516900 700800
rect 517100 700600 517300 700800
rect 517500 700600 517700 700800
rect 517900 700600 518100 700800
rect 518300 700600 518500 700800
rect 518700 700600 518900 700800
rect 519100 700600 519300 700800
rect 519500 700600 519700 700800
rect 519900 700600 520100 700800
rect 520300 700600 520500 700800
rect 520700 700600 521000 700800
rect 515500 700400 521000 700600
rect 515500 700200 515700 700400
rect 515900 700200 516100 700400
rect 516300 700200 516500 700400
rect 516700 700200 516900 700400
rect 517100 700200 517300 700400
rect 517500 700200 517700 700400
rect 517900 700200 518100 700400
rect 518300 700200 518500 700400
rect 518700 700200 518900 700400
rect 519100 700200 519300 700400
rect 519500 700200 519700 700400
rect 519900 700200 520100 700400
rect 520300 700200 520500 700400
rect 520700 700200 521000 700400
rect 515500 700000 521000 700200
rect 515500 699800 515700 700000
rect 515900 699800 516100 700000
rect 516300 699800 516500 700000
rect 516700 699800 516900 700000
rect 517100 699800 517300 700000
rect 517500 699800 517700 700000
rect 517900 699800 518100 700000
rect 518300 699800 518500 700000
rect 518700 699800 518900 700000
rect 519100 699800 519300 700000
rect 519500 699800 519700 700000
rect 519900 699800 520100 700000
rect 520300 699800 520500 700000
rect 520700 699800 521000 700000
rect 515500 699600 521000 699800
rect 515500 699400 515700 699600
rect 515900 699400 516100 699600
rect 516300 699400 516500 699600
rect 516700 699400 516900 699600
rect 517100 699400 517300 699600
rect 517500 699400 517700 699600
rect 517900 699400 518100 699600
rect 518300 699400 518500 699600
rect 518700 699400 518900 699600
rect 519100 699400 519300 699600
rect 519500 699400 519700 699600
rect 519900 699400 520100 699600
rect 520300 699400 520500 699600
rect 520700 699400 521000 699600
rect 515500 699200 521000 699400
rect 515500 699000 515700 699200
rect 515900 699000 516100 699200
rect 516300 699000 516500 699200
rect 516700 699000 516900 699200
rect 517100 699000 517300 699200
rect 517500 699000 517700 699200
rect 517900 699000 518100 699200
rect 518300 699000 518500 699200
rect 518700 699000 518900 699200
rect 519100 699000 519300 699200
rect 519500 699000 519700 699200
rect 519900 699000 520100 699200
rect 520300 699000 520500 699200
rect 520700 699000 521000 699200
rect 515500 698500 521000 699000
rect 12800 698200 21200 698400
rect 12800 698000 13000 698200
rect 13200 698000 13600 698200
rect 13800 698000 21200 698200
rect 12800 697800 21200 698000
rect 12800 697600 13000 697800
rect 13200 697600 13600 697800
rect 13800 697600 21200 697800
rect 12800 697200 21200 697600
rect 12800 697000 13000 697200
rect 13200 697000 13600 697200
rect 13800 697000 21200 697200
rect 12800 696800 21200 697000
rect 12800 696600 13000 696800
rect 13200 696600 13600 696800
rect 13800 696600 21200 696800
rect 12800 696400 21200 696600
rect 12800 691900 14120 691980
rect 12800 691700 12900 691900
rect 13100 691700 13200 691900
rect 13400 691700 13500 691900
rect 13700 691700 13800 691900
rect 14000 691700 14120 691900
rect 12800 674100 14120 691700
rect 16200 688700 21200 696400
rect 16200 688500 16400 688700
rect 16600 688500 16800 688700
rect 17000 688500 17200 688700
rect 17400 688500 17600 688700
rect 17800 688500 18000 688700
rect 18200 688500 18400 688700
rect 18600 688500 18800 688700
rect 19000 688500 19200 688700
rect 19400 688500 19600 688700
rect 19800 688500 20000 688700
rect 20200 688500 20400 688700
rect 20600 688500 20800 688700
rect 21000 688500 21200 688700
rect 16200 688300 21200 688500
rect 16200 688100 16400 688300
rect 16600 688100 16800 688300
rect 17000 688100 17200 688300
rect 17400 688100 17600 688300
rect 17800 688100 18000 688300
rect 18200 688100 18400 688300
rect 18600 688100 18800 688300
rect 19000 688100 19200 688300
rect 19400 688100 19600 688300
rect 19800 688100 20000 688300
rect 20200 688100 20400 688300
rect 20600 688100 20800 688300
rect 21000 688100 21200 688300
rect 16200 688000 21200 688100
rect 23200 698200 24600 698400
rect 23200 698000 23400 698200
rect 23600 698000 23800 698200
rect 24000 698000 24200 698200
rect 24400 698000 24600 698200
rect 23200 697800 24600 698000
rect 23200 697600 23400 697800
rect 23600 697600 23800 697800
rect 24000 697600 24200 697800
rect 24400 697600 24600 697800
rect 23200 697400 24600 697600
rect 23200 697200 23400 697400
rect 23600 697200 23800 697400
rect 24000 697200 24200 697400
rect 24400 697200 24600 697400
rect 23200 697000 24600 697200
rect 23200 696800 23400 697000
rect 23600 696800 23800 697000
rect 24000 696800 24200 697000
rect 24400 696800 24600 697000
rect 23200 696600 24600 696800
rect 23200 696400 23400 696600
rect 23600 696400 23800 696600
rect 24000 696400 24200 696600
rect 24400 696400 24600 696600
rect 12800 673800 12900 674100
rect 13200 673800 13700 674100
rect 14000 673800 14120 674100
rect 12800 673600 14120 673800
rect 12800 673300 12900 673600
rect 13200 673300 13700 673600
rect 14000 673300 14120 673600
rect 12800 673100 14120 673300
rect 12800 672800 12900 673100
rect 13200 672800 13700 673100
rect 14000 672800 14120 673100
rect 12800 672700 14120 672800
rect 2499 648600 2801 648601
rect 2499 648300 2500 648600
rect 2800 648300 2801 648600
rect 2499 648299 2801 648300
rect 2999 648600 3301 648601
rect 2999 648300 3000 648600
rect 3300 648300 3301 648600
rect 2999 648299 3301 648300
rect 3499 648600 3801 648601
rect 3499 648300 3500 648600
rect 3800 648300 3801 648600
rect 3499 648299 3801 648300
rect 23200 648500 24600 696400
rect 57800 698200 66000 698400
rect 57800 698000 65000 698200
rect 65200 698000 65600 698200
rect 65800 698000 66000 698200
rect 57800 697800 66000 698000
rect 57800 697600 65000 697800
rect 65200 697600 65600 697800
rect 65800 697600 66000 697800
rect 57800 697400 66000 697600
rect 57800 697200 65000 697400
rect 65200 697200 65600 697400
rect 65800 697200 66000 697400
rect 57800 697000 66000 697200
rect 57800 696800 65000 697000
rect 65200 696800 65600 697000
rect 65800 696800 66000 697000
rect 57800 696600 66000 696800
rect 57800 696400 65000 696600
rect 65200 696400 65600 696600
rect 65800 696400 66000 696600
rect 57800 696200 66000 696400
rect 68200 698200 76400 698400
rect 68200 698000 75400 698200
rect 75600 698000 76000 698200
rect 76200 698000 76400 698200
rect 68200 697800 76400 698000
rect 68200 697600 75400 697800
rect 75600 697600 76000 697800
rect 76200 697600 76400 697800
rect 68200 697400 76400 697600
rect 68200 697200 75400 697400
rect 75600 697200 76000 697400
rect 76200 697200 76400 697400
rect 68200 697000 76400 697200
rect 68200 696800 75400 697000
rect 75600 696800 76000 697000
rect 76200 696800 76400 697000
rect 68200 696600 76400 696800
rect 68200 696400 75400 696600
rect 75600 696400 76000 696600
rect 76200 696400 76400 696600
rect 68200 696200 76400 696400
rect 515500 697400 521000 697940
rect 515500 697200 515700 697400
rect 515900 697200 516100 697400
rect 516300 697200 516500 697400
rect 516700 697200 516900 697400
rect 517100 697200 517300 697400
rect 517500 697200 517700 697400
rect 517900 697200 518100 697400
rect 518300 697200 518500 697400
rect 518700 697200 518900 697400
rect 519100 697200 519300 697400
rect 519500 697200 519700 697400
rect 519900 697200 520100 697400
rect 520300 697200 520500 697400
rect 520700 697200 521000 697400
rect 515500 697000 521000 697200
rect 515500 696800 515700 697000
rect 515900 696800 516100 697000
rect 516300 696800 516500 697000
rect 516700 696800 516900 697000
rect 517100 696800 517300 697000
rect 517500 696800 517700 697000
rect 517900 696800 518100 697000
rect 518300 696800 518500 697000
rect 518700 696800 518900 697000
rect 519100 696800 519300 697000
rect 519500 696800 519700 697000
rect 519900 696800 520100 697000
rect 520300 696800 520500 697000
rect 520700 696800 521000 697000
rect 515500 696600 521000 696800
rect 515500 696400 515700 696600
rect 515900 696400 516100 696600
rect 516300 696400 516500 696600
rect 516700 696400 516900 696600
rect 517100 696400 517300 696600
rect 517500 696400 517700 696600
rect 517900 696400 518100 696600
rect 518300 696400 518500 696600
rect 518700 696400 518900 696600
rect 519100 696400 519300 696600
rect 519500 696400 519700 696600
rect 519900 696400 520100 696600
rect 520300 696400 520500 696600
rect 520700 696400 521000 696600
rect 38699 693000 38861 693001
rect 38699 692840 38700 693000
rect 38860 692840 38861 693000
rect 38699 692839 38861 692840
rect 39119 693000 39281 693001
rect 39119 692840 39120 693000
rect 39280 692840 39281 693000
rect 49959 693000 50101 693001
rect 49959 692860 49960 693000
rect 50100 692860 50101 693000
rect 49959 692859 50101 692860
rect 50179 693000 50321 693001
rect 50179 692860 50180 693000
rect 50320 692860 50321 693000
rect 50179 692859 50321 692860
rect 50399 693000 50541 693001
rect 50399 692860 50400 693000
rect 50540 692860 50541 693000
rect 50399 692859 50541 692860
rect 39119 692839 39281 692840
rect 49959 692800 50101 692801
rect 38699 692780 38861 692781
rect 38699 692620 38700 692780
rect 38860 692620 38861 692780
rect 38699 692619 38861 692620
rect 39119 692780 39281 692781
rect 39119 692620 39120 692780
rect 39280 692620 39281 692780
rect 49959 692660 49960 692800
rect 50100 692660 50101 692800
rect 49959 692659 50101 692660
rect 50179 692800 50321 692801
rect 50179 692660 50180 692800
rect 50320 692660 50321 692800
rect 50179 692659 50321 692660
rect 50399 692800 50541 692801
rect 50399 692660 50400 692800
rect 50540 692660 50541 692800
rect 50399 692659 50541 692660
rect 39119 692619 39281 692620
rect 38699 692560 38861 692561
rect 38699 692400 38700 692560
rect 38860 692400 38861 692560
rect 38699 692399 38861 692400
rect 39119 692560 39281 692561
rect 39119 692400 39120 692560
rect 39280 692400 39281 692560
rect 39119 692399 39281 692400
rect 38699 692340 38861 692341
rect 38699 692180 38700 692340
rect 38860 692180 38861 692340
rect 38699 692179 38861 692180
rect 39119 692340 39281 692341
rect 39119 692180 39120 692340
rect 39280 692180 39281 692340
rect 39119 692179 39281 692180
rect 57800 691900 62200 696200
rect 57800 691700 58000 691900
rect 58200 691700 58400 691900
rect 58600 691700 58800 691900
rect 59000 691700 59200 691900
rect 59400 691700 59600 691900
rect 59800 691700 60000 691900
rect 60200 691700 60400 691900
rect 60600 691700 60800 691900
rect 61000 691700 61200 691900
rect 61400 691700 61600 691900
rect 61800 691700 62200 691900
rect 36600 687300 38400 687400
rect 36600 687100 36800 687300
rect 37000 687100 37200 687300
rect 37400 687100 37600 687300
rect 37800 687100 38000 687300
rect 38200 687100 38400 687300
rect 36600 685300 38400 687100
rect 36600 685100 36800 685300
rect 37000 685100 37200 685300
rect 37400 685100 37600 685300
rect 37800 685100 38000 685300
rect 38200 685100 38400 685300
rect 36600 684900 38400 685100
rect 36600 684700 36800 684900
rect 37000 684700 37200 684900
rect 37400 684700 37600 684900
rect 37800 684700 38000 684900
rect 38200 684700 38400 684900
rect 36600 684500 38400 684700
rect 36600 684300 36800 684500
rect 37000 684300 37200 684500
rect 37400 684300 37600 684500
rect 37800 684300 38000 684500
rect 38200 684300 38400 684500
rect 36600 684100 38400 684300
rect 36600 683900 36800 684100
rect 37000 683900 37200 684100
rect 37400 683900 37600 684100
rect 37800 683900 38000 684100
rect 38200 683900 38400 684100
rect 36600 683700 38400 683900
rect 36600 683500 36800 683700
rect 37000 683500 37200 683700
rect 37400 683500 37600 683700
rect 37800 683500 38000 683700
rect 38200 683500 38400 683700
rect 36600 683300 38400 683500
rect 36600 683100 36800 683300
rect 37000 683100 37200 683300
rect 37400 683100 37600 683300
rect 37800 683100 38000 683300
rect 38200 683100 38400 683300
rect 36600 682900 38400 683100
rect 36600 682700 36800 682900
rect 37000 682700 37200 682900
rect 37400 682700 37600 682900
rect 37800 682700 38000 682900
rect 38200 682700 38400 682900
rect 36600 682500 38400 682700
rect 36600 682300 36800 682500
rect 37000 682300 37200 682500
rect 37400 682300 37600 682500
rect 37800 682300 38000 682500
rect 38200 682300 38400 682500
rect 36600 682100 38400 682300
rect 36600 681900 36800 682100
rect 37000 681900 37200 682100
rect 37400 681900 37600 682100
rect 37800 681900 38000 682100
rect 38200 681900 38400 682100
rect 36600 681700 38400 681900
rect 36600 681500 36800 681700
rect 37000 681500 37200 681700
rect 37400 681500 37600 681700
rect 37800 681500 38000 681700
rect 38200 681500 38400 681700
rect 36600 681300 38400 681500
rect 36600 681100 36800 681300
rect 37000 681100 37200 681300
rect 37400 681100 37600 681300
rect 37800 681100 38000 681300
rect 38200 681100 38400 681300
rect 36600 680900 38400 681100
rect 36600 680700 36800 680900
rect 37000 680700 37200 680900
rect 37400 680700 37600 680900
rect 37800 680700 38000 680900
rect 38200 680700 38400 680900
rect 36600 680500 38400 680700
rect 36600 680300 36800 680500
rect 37000 680300 37200 680500
rect 37400 680300 37600 680500
rect 37800 680300 38000 680500
rect 38200 680300 38400 680500
rect 36600 680200 38400 680300
rect 38670 675000 39330 686050
rect 23200 648200 23400 648500
rect 23700 648200 24100 648500
rect 24400 648200 24600 648500
rect 2499 648100 2801 648101
rect 2499 647800 2500 648100
rect 2800 647800 2801 648100
rect 2499 647799 2801 647800
rect 2999 648100 3301 648101
rect 2999 647800 3000 648100
rect 3300 647800 3301 648100
rect 2999 647799 3301 647800
rect 3499 648100 3801 648101
rect 3499 647800 3500 648100
rect 3800 647800 3801 648100
rect 3499 647799 3801 647800
rect 23200 647900 24600 648200
rect 2499 647600 2801 647601
rect 2499 647300 2500 647600
rect 2800 647300 2801 647600
rect 2499 647299 2801 647300
rect 2999 647600 3301 647601
rect 2999 647300 3000 647600
rect 3300 647300 3301 647600
rect 2999 647299 3301 647300
rect 3499 647600 3801 647601
rect 3499 647300 3500 647600
rect 3800 647300 3801 647600
rect 3499 647299 3801 647300
rect 23200 647600 23400 647900
rect 23700 647600 24100 647900
rect 24400 647600 24600 647900
rect 23200 647300 24600 647600
rect 2499 647100 2801 647101
rect 2499 646800 2500 647100
rect 2800 646800 2801 647100
rect 2499 646799 2801 646800
rect 2999 647100 3301 647101
rect 2999 646800 3000 647100
rect 3300 646800 3301 647100
rect 2999 646799 3301 646800
rect 3499 647100 3801 647101
rect 3499 646800 3500 647100
rect 3800 646800 3801 647100
rect 3499 646799 3801 646800
rect 23200 647000 23400 647300
rect 23700 647000 24100 647300
rect 24400 647000 24600 647300
rect 2499 646600 2801 646601
rect 2499 646300 2500 646600
rect 2800 646300 2801 646600
rect 2499 646299 2801 646300
rect 2999 646600 3301 646601
rect 2999 646300 3000 646600
rect 3300 646300 3301 646600
rect 2999 646299 3301 646300
rect 3499 646600 3801 646601
rect 3499 646300 3500 646600
rect 3800 646300 3801 646600
rect 3499 646299 3801 646300
rect 23200 646600 24600 647000
rect 23200 646300 23400 646600
rect 23700 646300 24100 646600
rect 24400 646300 24600 646600
rect 2499 646100 2801 646101
rect 2499 645800 2500 646100
rect 2800 645800 2801 646100
rect 2499 645799 2801 645800
rect 2999 646100 3301 646101
rect 2999 645800 3000 646100
rect 3300 645800 3301 646100
rect 2999 645799 3301 645800
rect 3499 646100 3801 646101
rect 3499 645800 3500 646100
rect 3800 645800 3801 646100
rect 3499 645799 3801 645800
rect 23200 646000 24600 646300
rect 23200 645700 23400 646000
rect 23700 645700 24100 646000
rect 24400 645700 24600 646000
rect 2499 645600 2801 645601
rect 2499 645300 2500 645600
rect 2800 645300 2801 645600
rect 2499 645299 2801 645300
rect 2999 645600 3301 645601
rect 2999 645300 3000 645600
rect 3300 645300 3301 645600
rect 2999 645299 3301 645300
rect 3499 645600 3801 645601
rect 3499 645300 3500 645600
rect 3800 645300 3801 645600
rect 3499 645299 3801 645300
rect 23200 645400 24600 645700
rect 2499 645100 2801 645101
rect 2499 644800 2500 645100
rect 2800 644800 2801 645100
rect 2499 644799 2801 644800
rect 2999 645100 3301 645101
rect 2999 644800 3000 645100
rect 3300 644800 3301 645100
rect 2999 644799 3301 644800
rect 3499 645100 3801 645101
rect 3499 644800 3500 645100
rect 3800 644800 3801 645100
rect 3499 644799 3801 644800
rect 23200 645100 23400 645400
rect 23700 645100 24100 645400
rect 24400 645100 24600 645400
rect 23200 644800 24600 645100
rect 2499 644600 2801 644601
rect 2499 644300 2500 644600
rect 2800 644300 2801 644600
rect 2499 644299 2801 644300
rect 2999 644600 3301 644601
rect 2999 644300 3000 644600
rect 3300 644300 3301 644600
rect 2999 644299 3301 644300
rect 3499 644600 3801 644601
rect 3499 644300 3500 644600
rect 3800 644300 3801 644600
rect 3499 644299 3801 644300
rect 23200 644500 23400 644800
rect 23700 644500 24100 644800
rect 24400 644500 24600 644800
rect 23200 644200 24600 644500
rect 2499 644100 2801 644101
rect 2499 643800 2500 644100
rect 2800 643800 2801 644100
rect 2499 643799 2801 643800
rect 2999 644100 3301 644101
rect 2999 643800 3000 644100
rect 3300 643800 3301 644100
rect 2999 643799 3301 643800
rect 3499 644100 3801 644101
rect 3499 643800 3500 644100
rect 3800 643800 3801 644100
rect 3499 643799 3801 643800
rect 23200 643900 23400 644200
rect 23700 643900 24100 644200
rect 24400 643900 24600 644200
rect 2499 643600 2801 643601
rect 2499 643300 2500 643600
rect 2800 643300 2801 643600
rect 2499 643299 2801 643300
rect 2999 643600 3301 643601
rect 2999 643300 3000 643600
rect 3300 643300 3301 643600
rect 2999 643299 3301 643300
rect 3499 643600 3801 643601
rect 3499 643300 3500 643600
rect 3800 643300 3801 643600
rect 3499 643299 3801 643300
rect 23200 643600 24600 643900
rect 23200 643300 23400 643600
rect 23700 643300 24100 643600
rect 24400 643300 24600 643600
rect 2499 643100 2801 643101
rect 2499 642800 2500 643100
rect 2800 642800 2801 643100
rect 2499 642799 2801 642800
rect 2999 643100 3301 643101
rect 2999 642800 3000 643100
rect 3300 642800 3301 643100
rect 2999 642799 3301 642800
rect 3499 643100 3801 643101
rect 3499 642800 3500 643100
rect 3800 642800 3801 643100
rect 3499 642799 3801 642800
rect 23200 642900 24600 643300
rect 2499 642600 2801 642601
rect 2499 642300 2500 642600
rect 2800 642300 2801 642600
rect 2499 642299 2801 642300
rect 2999 642600 3301 642601
rect 2999 642300 3000 642600
rect 3300 642300 3301 642600
rect 2999 642299 3301 642300
rect 3499 642600 3801 642601
rect 3499 642300 3500 642600
rect 3800 642300 3801 642600
rect 3499 642299 3801 642300
rect 23200 642600 23400 642900
rect 23700 642600 24100 642900
rect 24400 642600 24600 642900
rect 23200 642300 24600 642600
rect 2499 642100 2801 642101
rect 2499 641800 2500 642100
rect 2800 641800 2801 642100
rect 2499 641799 2801 641800
rect 2999 642100 3301 642101
rect 2999 641800 3000 642100
rect 3300 641800 3301 642100
rect 2999 641799 3301 641800
rect 3499 642100 3801 642101
rect 3499 641800 3500 642100
rect 3800 641800 3801 642100
rect 3499 641799 3801 641800
rect 23200 642000 23400 642300
rect 23700 642000 24100 642300
rect 24400 642000 24600 642300
rect 23200 641700 24600 642000
rect 2499 641600 2801 641601
rect 2499 641300 2500 641600
rect 2800 641300 2801 641600
rect 2499 641299 2801 641300
rect 2999 641600 3301 641601
rect 2999 641300 3000 641600
rect 3300 641300 3301 641600
rect 2999 641299 3301 641300
rect 3499 641600 3801 641601
rect 3499 641300 3500 641600
rect 3800 641300 3801 641600
rect 3499 641299 3801 641300
rect 23200 641400 23400 641700
rect 23700 641400 24100 641700
rect 24400 641400 24600 641700
rect 2499 641100 2801 641101
rect 2499 640800 2500 641100
rect 2800 640800 2801 641100
rect 2499 640799 2801 640800
rect 2999 641100 3301 641101
rect 2999 640800 3000 641100
rect 3300 640800 3301 641100
rect 2999 640799 3301 640800
rect 3499 641100 3801 641101
rect 3499 640800 3500 641100
rect 3800 640800 3801 641100
rect 3499 640799 3801 640800
rect 23200 641100 24600 641400
rect 23200 640800 23400 641100
rect 23700 640800 24100 641100
rect 24400 640800 24600 641100
rect 2499 640600 2801 640601
rect 2499 640300 2500 640600
rect 2800 640300 2801 640600
rect 2499 640299 2801 640300
rect 2999 640600 3301 640601
rect 2999 640300 3000 640600
rect 3300 640300 3301 640600
rect 2999 640299 3301 640300
rect 3499 640600 3801 640601
rect 3499 640300 3500 640600
rect 3800 640300 3801 640600
rect 3499 640299 3801 640300
rect 23200 640500 24600 640800
rect 23200 640200 23400 640500
rect 23700 640200 24100 640500
rect 24400 640200 24600 640500
rect 2499 640100 2801 640101
rect 2499 639800 2500 640100
rect 2800 639800 2801 640100
rect 2499 639799 2801 639800
rect 2999 640100 3301 640101
rect 2999 639800 3000 640100
rect 3300 639800 3301 640100
rect 2999 639799 3301 639800
rect 3499 640100 3801 640101
rect 3499 639800 3500 640100
rect 3800 639800 3801 640100
rect 3499 639799 3801 639800
rect 23200 639900 24600 640200
rect 2499 639600 2801 639601
rect 2499 639300 2500 639600
rect 2800 639300 2801 639600
rect 2499 639299 2801 639300
rect 2999 639600 3301 639601
rect 2999 639300 3000 639600
rect 3300 639300 3301 639600
rect 2999 639299 3301 639300
rect 3499 639600 3801 639601
rect 3499 639300 3500 639600
rect 3800 639300 3801 639600
rect 3499 639299 3801 639300
rect 23200 639600 23400 639900
rect 23700 639600 24100 639900
rect 24400 639600 24600 639900
rect 23200 639300 24600 639600
rect 2499 639100 2801 639101
rect 2499 638800 2500 639100
rect 2800 638800 2801 639100
rect 2499 638799 2801 638800
rect 2999 639100 3301 639101
rect 2999 638800 3000 639100
rect 3300 638800 3301 639100
rect 2999 638799 3301 638800
rect 3499 639100 3801 639101
rect 3499 638800 3500 639100
rect 3800 638800 3801 639100
rect 3499 638799 3801 638800
rect 23200 639000 23400 639300
rect 23700 639000 24100 639300
rect 24400 639000 24600 639300
rect 23200 638700 24600 639000
rect 2499 638600 2801 638601
rect 2499 638300 2500 638600
rect 2800 638300 2801 638600
rect 2499 638299 2801 638300
rect 2999 638600 3301 638601
rect 2999 638300 3000 638600
rect 3300 638300 3301 638600
rect 2999 638299 3301 638300
rect 3499 638600 3801 638601
rect 3499 638300 3500 638600
rect 3800 638300 3801 638600
rect 3499 638299 3801 638300
rect 23200 638400 23400 638700
rect 23700 638400 24100 638700
rect 24400 638400 24600 638700
rect 2499 638100 2801 638101
rect 2499 637800 2500 638100
rect 2800 637800 2801 638100
rect 2499 637799 2801 637800
rect 2999 638100 3301 638101
rect 2999 637800 3000 638100
rect 3300 637800 3301 638100
rect 2999 637799 3301 637800
rect 3499 638100 3801 638101
rect 3499 637800 3500 638100
rect 3800 637800 3801 638100
rect 3499 637799 3801 637800
rect 23200 638100 24600 638400
rect 23200 637800 23400 638100
rect 23700 637800 24100 638100
rect 24400 637800 24600 638100
rect 2499 637600 2801 637601
rect 2499 637300 2500 637600
rect 2800 637300 2801 637600
rect 2499 637299 2801 637300
rect 2999 637600 3301 637601
rect 2999 637300 3000 637600
rect 3300 637300 3301 637600
rect 2999 637299 3301 637300
rect 3499 637600 3801 637601
rect 3499 637300 3500 637600
rect 3800 637300 3801 637600
rect 3499 637299 3801 637300
rect 23200 637400 24600 637800
rect 2499 637100 2801 637101
rect 2499 636800 2500 637100
rect 2800 636800 2801 637100
rect 2499 636799 2801 636800
rect 2999 637100 3301 637101
rect 2999 636800 3000 637100
rect 3300 636800 3301 637100
rect 2999 636799 3301 636800
rect 3499 637100 3801 637101
rect 3499 636800 3500 637100
rect 3800 636800 3801 637100
rect 3499 636799 3801 636800
rect 23200 637100 23400 637400
rect 23700 637100 24100 637400
rect 24400 637100 24600 637400
rect 23200 636700 24600 637100
rect 2499 636600 2801 636601
rect 2499 636300 2500 636600
rect 2800 636300 2801 636600
rect 2499 636299 2801 636300
rect 2999 636600 3301 636601
rect 2999 636300 3000 636600
rect 3300 636300 3301 636600
rect 2999 636299 3301 636300
rect 3499 636600 3801 636601
rect 3499 636300 3500 636600
rect 3800 636300 3801 636600
rect 3499 636299 3801 636300
rect 23200 636400 23400 636700
rect 23700 636400 24100 636700
rect 24400 636400 24600 636700
rect 2499 636100 2801 636101
rect 2499 635800 2500 636100
rect 2800 635800 2801 636100
rect 2499 635799 2801 635800
rect 2999 636100 3301 636101
rect 2999 635800 3000 636100
rect 3300 635800 3301 636100
rect 2999 635799 3301 635800
rect 3499 636100 3801 636101
rect 3499 635800 3500 636100
rect 3800 635800 3801 636100
rect 3499 635799 3801 635800
rect 23200 636000 24600 636400
rect 23200 635700 23400 636000
rect 23700 635700 24100 636000
rect 24400 635700 24600 636000
rect 2499 635600 2801 635601
rect 2499 635300 2500 635600
rect 2800 635300 2801 635600
rect 2499 635299 2801 635300
rect 2999 635600 3301 635601
rect 2999 635300 3000 635600
rect 3300 635300 3301 635600
rect 2999 635299 3301 635300
rect 3499 635600 3801 635601
rect 3499 635300 3500 635600
rect 3800 635300 3801 635600
rect 3499 635299 3801 635300
rect 23200 635200 24600 635700
rect 2499 635100 2801 635101
rect 2499 634800 2500 635100
rect 2800 634800 2801 635100
rect 2499 634799 2801 634800
rect 2999 635100 3301 635101
rect 2999 634800 3000 635100
rect 3300 634800 3301 635100
rect 2999 634799 3301 634800
rect 3499 635100 3801 635101
rect 3499 634800 3500 635100
rect 3800 634800 3801 635100
rect 3499 634799 3801 634800
rect 23200 634900 23400 635200
rect 23700 634900 24100 635200
rect 24400 634900 24600 635200
rect 2499 634600 2801 634601
rect 2499 634300 2500 634600
rect 2800 634300 2801 634600
rect 2499 634299 2801 634300
rect 2999 634600 3301 634601
rect 2999 634300 3000 634600
rect 3300 634300 3301 634600
rect 2999 634299 3301 634300
rect 3499 634600 3801 634601
rect 3499 634300 3500 634600
rect 3800 634300 3801 634600
rect 3499 634299 3801 634300
rect 23200 634500 24600 634900
rect 23200 634200 23400 634500
rect 23700 634200 24100 634500
rect 24400 634200 24600 634500
rect 23200 633800 24600 634200
rect 32600 674000 40800 675000
rect 32600 673700 32800 674000
rect 33100 673700 33300 674000
rect 33600 673700 33800 674000
rect 34100 673700 34300 674000
rect 34600 673700 34800 674000
rect 35100 673700 35300 674000
rect 35600 673700 35800 674000
rect 36100 673700 36300 674000
rect 36600 673700 36800 674000
rect 37100 673700 37300 674000
rect 37600 673700 37800 674000
rect 38100 673700 38300 674000
rect 38600 673700 38800 674000
rect 39100 673700 39300 674000
rect 39600 673700 39800 674000
rect 40100 673700 40300 674000
rect 40600 673700 40800 674000
rect 32600 673200 40800 673700
rect 32600 672900 32800 673200
rect 33100 672900 33300 673200
rect 33600 672900 33800 673200
rect 34100 672900 34300 673200
rect 34600 672900 34800 673200
rect 35100 672900 35300 673200
rect 35600 672900 35800 673200
rect 36100 672900 36300 673200
rect 36600 672900 36800 673200
rect 37100 672900 37300 673200
rect 37600 672900 37800 673200
rect 38100 672900 38300 673200
rect 38600 672900 38800 673200
rect 39100 672900 39300 673200
rect 39600 672900 39800 673200
rect 40100 672900 40300 673200
rect 40600 672900 40800 673200
rect 32600 670700 40800 672900
rect 49920 674000 50580 686100
rect 49920 673700 50100 674000
rect 50400 673700 50580 674000
rect 49920 673600 50580 673700
rect 49920 673300 50100 673600
rect 50400 673300 50580 673600
rect 49920 673200 50580 673300
rect 49920 672900 50100 673200
rect 50400 672900 50580 673200
rect 49920 672700 50580 672900
rect 57800 682200 62200 691700
rect 68200 690200 73200 696200
rect 68200 690000 68400 690200
rect 68600 690000 68800 690200
rect 69000 690000 69200 690200
rect 69400 690000 69600 690200
rect 69800 690000 70000 690200
rect 70200 690000 70400 690200
rect 70600 690000 70800 690200
rect 71000 690000 71200 690200
rect 71400 690000 71600 690200
rect 71800 690000 72000 690200
rect 72200 690000 72400 690200
rect 72600 690000 72800 690200
rect 73000 690000 73200 690200
rect 68200 689800 73200 690000
rect 68200 689600 68400 689800
rect 68600 689600 68800 689800
rect 69000 689600 69200 689800
rect 69400 689600 69600 689800
rect 69800 689600 70000 689800
rect 70200 689600 70400 689800
rect 70600 689600 70800 689800
rect 71000 689600 71200 689800
rect 71400 689600 71600 689800
rect 71800 689600 72000 689800
rect 72200 689600 72400 689800
rect 72600 689600 72800 689800
rect 73000 689600 73200 689800
rect 68200 689400 73200 689600
rect 57800 682000 58000 682200
rect 58200 682000 58400 682200
rect 58600 682000 58800 682200
rect 59000 682000 59200 682200
rect 59400 682000 59600 682200
rect 59800 682000 60000 682200
rect 60200 682000 60400 682200
rect 60600 682000 60800 682200
rect 61000 682000 61200 682200
rect 61400 682000 61600 682200
rect 61800 682000 62200 682200
rect 32600 670400 32800 670700
rect 33100 670400 33300 670700
rect 33600 670400 33800 670700
rect 34100 670400 34300 670700
rect 34600 670400 34800 670700
rect 35100 670400 35300 670700
rect 35600 670400 35800 670700
rect 36100 670400 36300 670700
rect 36600 670400 36800 670700
rect 37100 670400 37300 670700
rect 37600 670400 37800 670700
rect 38100 670400 38300 670700
rect 38600 670400 38800 670700
rect 39100 670400 39300 670700
rect 39600 670400 39800 670700
rect 40100 670400 40300 670700
rect 40600 670400 40800 670700
rect 32600 670000 40800 670400
rect 32600 669700 32800 670000
rect 33100 669700 33300 670000
rect 33600 669700 33800 670000
rect 34100 669700 34300 670000
rect 34600 669700 34800 670000
rect 35100 669700 35300 670000
rect 35600 669700 35800 670000
rect 36100 669700 36300 670000
rect 36600 669700 36800 670000
rect 37100 669700 37300 670000
rect 37600 669700 37800 670000
rect 38100 669700 38300 670000
rect 38600 669700 38800 670000
rect 39100 669700 39300 670000
rect 39600 669700 39800 670000
rect 40100 669700 40300 670000
rect 40600 669700 40800 670000
rect 32600 667400 40800 669700
rect 32600 667100 32800 667400
rect 33100 667100 33300 667400
rect 33600 667100 33800 667400
rect 34100 667100 34300 667400
rect 34600 667100 34800 667400
rect 35100 667100 35300 667400
rect 35600 667100 35800 667400
rect 36100 667100 36300 667400
rect 36600 667100 36800 667400
rect 37100 667100 37300 667400
rect 37600 667100 37800 667400
rect 38100 667100 38300 667400
rect 38600 667100 38800 667400
rect 39100 667100 39300 667400
rect 39600 667100 39800 667400
rect 40100 667100 40300 667400
rect 40600 667100 40800 667400
rect 32600 666700 40800 667100
rect 32600 666400 32800 666700
rect 33100 666400 33300 666700
rect 33600 666400 33800 666700
rect 34100 666400 34300 666700
rect 34600 666400 34800 666700
rect 35100 666400 35300 666700
rect 35600 666400 35800 666700
rect 36100 666400 36300 666700
rect 36600 666400 36800 666700
rect 37100 666400 37300 666700
rect 37600 666400 37800 666700
rect 38100 666400 38300 666700
rect 38600 666400 38800 666700
rect 39100 666400 39300 666700
rect 39600 666400 39800 666700
rect 40100 666400 40300 666700
rect 40600 666400 40800 666700
rect 32600 663300 40800 666400
rect 32600 663000 32800 663300
rect 33100 663000 33300 663300
rect 33600 663000 33800 663300
rect 34100 663000 34300 663300
rect 34600 663000 34800 663300
rect 35100 663000 35300 663300
rect 35600 663000 35800 663300
rect 36100 663000 36300 663300
rect 36600 663000 36800 663300
rect 37100 663000 37300 663300
rect 37600 663000 37800 663300
rect 38100 663000 38300 663300
rect 38600 663000 38800 663300
rect 39100 663000 39300 663300
rect 39600 663000 39800 663300
rect 40100 663000 40300 663300
rect 40600 663000 40800 663300
rect 32600 564100 40800 663000
rect 57800 648600 62200 682000
rect 515500 684800 521000 696400
rect 573100 698000 574220 698200
rect 573100 697800 573300 698000
rect 573500 697800 573800 698000
rect 574000 697800 574220 698000
rect 573100 697600 574220 697800
rect 573100 697400 573300 697600
rect 573500 697400 573800 697600
rect 574000 697400 574220 697600
rect 573100 697200 574220 697400
rect 573100 697000 573300 697200
rect 573500 697000 573800 697200
rect 574000 697000 574220 697200
rect 573100 696800 574220 697000
rect 573100 696600 573300 696800
rect 573500 696600 573800 696800
rect 574000 696600 574220 696800
rect 573100 696400 574220 696600
rect 573100 696200 573300 696400
rect 573500 696200 573800 696400
rect 574000 696200 574220 696400
rect 532200 690400 539200 690500
rect 532200 690200 532300 690400
rect 532500 690200 532700 690400
rect 532900 690200 533100 690400
rect 533300 690200 533500 690400
rect 533700 690200 533900 690400
rect 534100 690200 539200 690400
rect 532200 690100 539200 690200
rect 532200 689900 532300 690100
rect 532500 689900 532700 690100
rect 532900 689900 533100 690100
rect 533300 689900 533500 690100
rect 533700 689900 533900 690100
rect 534100 689900 539200 690100
rect 532200 689700 539200 689900
rect 532200 689500 532300 689700
rect 532500 689500 532700 689700
rect 532900 689500 533100 689700
rect 533300 689500 533500 689700
rect 533700 689500 533900 689700
rect 534100 689500 539200 689700
rect 532200 689300 539200 689500
rect 532200 689100 532300 689300
rect 532500 689100 532700 689300
rect 532900 689100 533100 689300
rect 533300 689100 533500 689300
rect 533700 689100 533900 689300
rect 534100 689100 539200 689300
rect 532200 688900 539200 689100
rect 532200 688700 532300 688900
rect 532500 688700 532700 688900
rect 532900 688700 533100 688900
rect 533300 688700 533500 688900
rect 533700 688700 533900 688900
rect 534100 688700 539200 688900
rect 532200 688600 539200 688700
rect 515500 684600 515700 684800
rect 515900 684600 516100 684800
rect 516300 684600 516500 684800
rect 516700 684600 516900 684800
rect 517100 684600 517300 684800
rect 517500 684600 517700 684800
rect 517900 684600 518100 684800
rect 518300 684600 518500 684800
rect 518700 684600 518900 684800
rect 519100 684600 519300 684800
rect 519500 684600 519700 684800
rect 519900 684600 520100 684800
rect 520300 684600 520500 684800
rect 520700 684600 521000 684800
rect 515500 684400 521000 684600
rect 515500 684200 515700 684400
rect 515900 684200 516100 684400
rect 516300 684200 516500 684400
rect 516700 684200 516900 684400
rect 517100 684200 517300 684400
rect 517500 684200 517700 684400
rect 517900 684200 518100 684400
rect 518300 684200 518500 684400
rect 518700 684200 518900 684400
rect 519100 684200 519300 684400
rect 519500 684200 519700 684400
rect 519900 684200 520100 684400
rect 520300 684200 520500 684400
rect 520700 684200 521000 684400
rect 515500 684000 521000 684200
rect 515500 683800 515700 684000
rect 515900 683800 516100 684000
rect 516300 683800 516500 684000
rect 516700 683800 516900 684000
rect 517100 683800 517300 684000
rect 517500 683800 517700 684000
rect 517900 683800 518100 684000
rect 518300 683800 518500 684000
rect 518700 683800 518900 684000
rect 519100 683800 519300 684000
rect 519500 683800 519700 684000
rect 519900 683800 520100 684000
rect 520300 683800 520500 684000
rect 520700 683800 521000 684000
rect 515500 683600 521000 683800
rect 515500 683400 515700 683600
rect 515900 683400 516100 683600
rect 516300 683400 516500 683600
rect 516700 683400 516900 683600
rect 517100 683400 517300 683600
rect 517500 683400 517700 683600
rect 517900 683400 518100 683600
rect 518300 683400 518500 683600
rect 518700 683400 518900 683600
rect 519100 683400 519300 683600
rect 519500 683400 519700 683600
rect 519900 683400 520100 683600
rect 520300 683400 520500 683600
rect 520700 683400 521000 683600
rect 515500 683200 521000 683400
rect 515500 683000 515700 683200
rect 515900 683000 516100 683200
rect 516300 683000 516500 683200
rect 516700 683000 516900 683200
rect 517100 683000 517300 683200
rect 517500 683000 517700 683200
rect 517900 683000 518100 683200
rect 518300 683000 518500 683200
rect 518700 683000 518900 683200
rect 519100 683000 519300 683200
rect 519500 683000 519700 683200
rect 519900 683000 520100 683200
rect 520300 683000 520500 683200
rect 520700 683000 521000 683200
rect 515500 682800 521000 683000
rect 515500 682600 515700 682800
rect 515900 682600 516100 682800
rect 516300 682600 516500 682800
rect 516700 682600 516900 682800
rect 517100 682600 517300 682800
rect 517500 682600 517700 682800
rect 517900 682600 518100 682800
rect 518300 682600 518500 682800
rect 518700 682600 518900 682800
rect 519100 682600 519300 682800
rect 519500 682600 519700 682800
rect 519900 682600 520100 682800
rect 520300 682600 520500 682800
rect 520700 682600 521000 682800
rect 515500 679200 521000 682600
rect 515500 679000 515900 679200
rect 516100 679000 516300 679200
rect 516500 679000 516700 679200
rect 516900 679000 517100 679200
rect 517300 679000 517500 679200
rect 517700 679000 517900 679200
rect 518100 679000 518300 679200
rect 518500 679000 518700 679200
rect 518900 679000 519100 679200
rect 519300 679000 519500 679200
rect 519700 679000 519900 679200
rect 520100 679000 520300 679200
rect 520500 679000 520700 679200
rect 520900 679000 521000 679200
rect 515500 678800 521000 679000
rect 515500 678600 515900 678800
rect 516100 678600 516300 678800
rect 516500 678600 516700 678800
rect 516900 678600 517100 678800
rect 517300 678600 517500 678800
rect 517700 678600 517900 678800
rect 518100 678600 518300 678800
rect 518500 678600 518700 678800
rect 518900 678600 519100 678800
rect 519300 678600 519500 678800
rect 519700 678600 519900 678800
rect 520100 678600 520300 678800
rect 520500 678600 520700 678800
rect 520900 678600 521000 678800
rect 515500 678400 521000 678600
rect 515500 678200 515900 678400
rect 516100 678200 516300 678400
rect 516500 678200 516700 678400
rect 516900 678200 517100 678400
rect 517300 678200 517500 678400
rect 517700 678200 517900 678400
rect 518100 678200 518300 678400
rect 518500 678200 518700 678400
rect 518900 678200 519100 678400
rect 519300 678200 519500 678400
rect 519700 678200 519900 678400
rect 520100 678200 520300 678400
rect 520500 678200 520700 678400
rect 520900 678200 521000 678400
rect 515500 678000 521000 678200
rect 515500 677800 515900 678000
rect 516100 677800 516300 678000
rect 516500 677800 516700 678000
rect 516900 677800 517100 678000
rect 517300 677800 517500 678000
rect 517700 677800 517900 678000
rect 518100 677800 518300 678000
rect 518500 677800 518700 678000
rect 518900 677800 519100 678000
rect 519300 677800 519500 678000
rect 519700 677800 519900 678000
rect 520100 677800 520300 678000
rect 520500 677800 520700 678000
rect 520900 677800 521000 678000
rect 515500 677600 521000 677800
rect 515500 677400 515900 677600
rect 516100 677400 516300 677600
rect 516500 677400 516700 677600
rect 516900 677400 517100 677600
rect 517300 677400 517500 677600
rect 517700 677400 517900 677600
rect 518100 677400 518300 677600
rect 518500 677400 518700 677600
rect 518900 677400 519100 677600
rect 519300 677400 519500 677600
rect 519700 677400 519900 677600
rect 520100 677400 520300 677600
rect 520500 677400 520700 677600
rect 520900 677400 521000 677600
rect 515500 677200 521000 677400
rect 515500 677000 515900 677200
rect 516100 677000 516300 677200
rect 516500 677000 516700 677200
rect 516900 677000 517100 677200
rect 517300 677000 517500 677200
rect 517700 677000 517900 677200
rect 518100 677000 518300 677200
rect 518500 677000 518700 677200
rect 518900 677000 519100 677200
rect 519300 677000 519500 677200
rect 519700 677000 519900 677200
rect 520100 677000 520300 677200
rect 520500 677000 520700 677200
rect 520900 677000 521000 677200
rect 515500 676800 521000 677000
rect 515500 676600 515900 676800
rect 516100 676600 516300 676800
rect 516500 676600 516700 676800
rect 516900 676600 517100 676800
rect 517300 676600 517500 676800
rect 517700 676600 517900 676800
rect 518100 676600 518300 676800
rect 518500 676600 518700 676800
rect 518900 676600 519100 676800
rect 519300 676600 519500 676800
rect 519700 676600 519900 676800
rect 520100 676600 520300 676800
rect 520500 676600 520700 676800
rect 520900 676600 521000 676800
rect 515500 676460 521000 676600
rect 549700 687300 553100 687400
rect 549700 687200 551200 687300
rect 549700 687000 549900 687200
rect 550100 687000 550200 687200
rect 550400 687000 550500 687200
rect 550700 687000 550800 687200
rect 551000 687100 551200 687200
rect 551400 687100 553100 687300
rect 551000 687000 553100 687100
rect 549700 686800 551200 687000
rect 551400 686800 553100 687000
rect 549700 686700 553100 686800
rect 549700 686500 551200 686700
rect 551400 686500 553100 686700
rect 549700 686400 553100 686500
rect 549700 686200 551200 686400
rect 551400 686200 553100 686400
rect 549700 686100 553100 686200
rect 549700 685900 549800 686100
rect 550000 685900 550100 686100
rect 550300 685900 550400 686100
rect 550600 685900 550800 686100
rect 551000 685900 553100 686100
rect 549700 684900 553100 685900
rect 549700 684600 549900 684900
rect 550200 684600 550400 684900
rect 550700 684600 550900 684900
rect 551200 684600 551400 684900
rect 551700 684600 551900 684900
rect 552200 684600 552400 684900
rect 552700 684600 553100 684900
rect 549700 684400 553100 684600
rect 549700 684100 549900 684400
rect 550200 684100 550400 684400
rect 550700 684100 550900 684400
rect 551200 684100 551400 684400
rect 551700 684100 551900 684400
rect 552200 684100 552400 684400
rect 552700 684100 553100 684400
rect 549700 683900 553100 684100
rect 549700 683600 549900 683900
rect 550200 683600 550400 683900
rect 550700 683600 550900 683900
rect 551200 683600 551400 683900
rect 551700 683600 551900 683900
rect 552200 683600 552400 683900
rect 552700 683600 553100 683900
rect 549700 681400 553100 683600
rect 573100 684900 574220 696200
rect 573100 684600 573200 684900
rect 573500 684600 573800 684900
rect 574100 684600 574220 684900
rect 573100 684400 574220 684600
rect 573100 684100 573200 684400
rect 573500 684100 573800 684400
rect 574100 684100 574220 684400
rect 576799 684700 577101 684701
rect 576799 684400 576800 684700
rect 577100 684400 577101 684700
rect 576799 684399 577101 684400
rect 577299 684700 577601 684701
rect 577299 684400 577300 684700
rect 577600 684400 577601 684700
rect 577299 684399 577601 684400
rect 577799 684700 578101 684701
rect 577799 684400 577800 684700
rect 578100 684400 578101 684700
rect 577799 684399 578101 684400
rect 578299 684700 578601 684701
rect 578299 684400 578300 684700
rect 578600 684400 578601 684700
rect 578299 684399 578601 684400
rect 573100 683900 574220 684100
rect 573100 683600 573200 683900
rect 573500 683600 573800 683900
rect 574100 683600 574220 683900
rect 576799 684200 577101 684201
rect 576799 683900 576800 684200
rect 577100 683900 577101 684200
rect 576799 683899 577101 683900
rect 577299 684200 577601 684201
rect 577299 683900 577300 684200
rect 577600 683900 577601 684200
rect 577299 683899 577601 683900
rect 577799 684200 578101 684201
rect 577799 683900 577800 684200
rect 578100 683900 578101 684200
rect 577799 683899 578101 683900
rect 578299 684200 578601 684201
rect 578299 683900 578300 684200
rect 578600 683900 578601 684200
rect 578299 683899 578601 683900
rect 573100 683400 574220 683600
rect 549700 681200 549800 681400
rect 550000 681200 550200 681400
rect 550400 681200 550600 681400
rect 550800 681200 551000 681400
rect 551200 681200 551400 681400
rect 551600 681200 551800 681400
rect 552000 681200 552200 681400
rect 552400 681200 552600 681400
rect 552800 681200 553100 681400
rect 549700 681000 553100 681200
rect 549700 680800 549800 681000
rect 550000 680800 550200 681000
rect 550400 680800 550600 681000
rect 550800 680800 551000 681000
rect 551200 680800 551400 681000
rect 551600 680800 551800 681000
rect 552000 680800 552200 681000
rect 552400 680800 552600 681000
rect 552800 680800 553100 681000
rect 57800 648300 58000 648600
rect 58300 648300 58500 648600
rect 58800 648300 59000 648600
rect 59300 648300 59500 648600
rect 59800 648300 60000 648600
rect 60300 648300 60500 648600
rect 60800 648300 61000 648600
rect 61300 648300 61500 648600
rect 61800 648300 62200 648600
rect 57800 648100 62200 648300
rect 57800 647800 58000 648100
rect 58300 647800 58500 648100
rect 58800 647800 59000 648100
rect 59300 647800 59500 648100
rect 59800 647800 60000 648100
rect 60300 647800 60500 648100
rect 60800 647800 61000 648100
rect 61300 647800 61500 648100
rect 61800 647800 62200 648100
rect 57800 647600 62200 647800
rect 57800 647300 58000 647600
rect 58300 647300 58500 647600
rect 58800 647300 59000 647600
rect 59300 647300 59500 647600
rect 59800 647300 60000 647600
rect 60300 647300 60500 647600
rect 60800 647300 61000 647600
rect 61300 647300 61500 647600
rect 61800 647300 62200 647600
rect 57800 647100 62200 647300
rect 57800 646800 58000 647100
rect 58300 646800 58500 647100
rect 58800 646800 59000 647100
rect 59300 646800 59500 647100
rect 59800 646800 60000 647100
rect 60300 646800 60500 647100
rect 60800 646800 61000 647100
rect 61300 646800 61500 647100
rect 61800 646800 62200 647100
rect 57800 646600 62200 646800
rect 57800 646300 58000 646600
rect 58300 646300 58500 646600
rect 58800 646300 59000 646600
rect 59300 646300 59500 646600
rect 59800 646300 60000 646600
rect 60300 646300 60500 646600
rect 60800 646300 61000 646600
rect 61300 646300 61500 646600
rect 61800 646300 62200 646600
rect 57800 646100 62200 646300
rect 57800 645800 58000 646100
rect 58300 645800 58500 646100
rect 58800 645800 59000 646100
rect 59300 645800 59500 646100
rect 59800 645800 60000 646100
rect 60300 645800 60500 646100
rect 60800 645800 61000 646100
rect 61300 645800 61500 646100
rect 61800 645800 62200 646100
rect 57800 645600 62200 645800
rect 57800 645300 58000 645600
rect 58300 645300 58500 645600
rect 58800 645300 59000 645600
rect 59300 645300 59500 645600
rect 59800 645300 60000 645600
rect 60300 645300 60500 645600
rect 60800 645300 61000 645600
rect 61300 645300 61500 645600
rect 61800 645300 62200 645600
rect 57800 645100 62200 645300
rect 57800 644800 58000 645100
rect 58300 644800 58500 645100
rect 58800 644800 59000 645100
rect 59300 644800 59500 645100
rect 59800 644800 60000 645100
rect 60300 644800 60500 645100
rect 60800 644800 61000 645100
rect 61300 644800 61500 645100
rect 61800 644800 62200 645100
rect 57800 644600 62200 644800
rect 57800 644300 58000 644600
rect 58300 644300 58500 644600
rect 58800 644300 59000 644600
rect 59300 644300 59500 644600
rect 59800 644300 60000 644600
rect 60300 644300 60500 644600
rect 60800 644300 61000 644600
rect 61300 644300 61500 644600
rect 61800 644300 62200 644600
rect 57800 644100 62200 644300
rect 57800 643800 58000 644100
rect 58300 643800 58500 644100
rect 58800 643800 59000 644100
rect 59300 643800 59500 644100
rect 59800 643800 60000 644100
rect 60300 643800 60500 644100
rect 60800 643800 61000 644100
rect 61300 643800 61500 644100
rect 61800 643800 62200 644100
rect 57800 643600 62200 643800
rect 57800 643300 58000 643600
rect 58300 643300 58500 643600
rect 58800 643300 59000 643600
rect 59300 643300 59500 643600
rect 59800 643300 60000 643600
rect 60300 643300 60500 643600
rect 60800 643300 61000 643600
rect 61300 643300 61500 643600
rect 61800 643300 62200 643600
rect 57800 643100 62200 643300
rect 57800 642800 58000 643100
rect 58300 642800 58500 643100
rect 58800 642800 59000 643100
rect 59300 642800 59500 643100
rect 59800 642800 60000 643100
rect 60300 642800 60500 643100
rect 60800 642800 61000 643100
rect 61300 642800 61500 643100
rect 61800 642800 62200 643100
rect 57800 642600 62200 642800
rect 57800 642300 58000 642600
rect 58300 642300 58500 642600
rect 58800 642300 59000 642600
rect 59300 642300 59500 642600
rect 59800 642300 60000 642600
rect 60300 642300 60500 642600
rect 60800 642300 61000 642600
rect 61300 642300 61500 642600
rect 61800 642300 62200 642600
rect 57800 642100 62200 642300
rect 57800 641800 58000 642100
rect 58300 641800 58500 642100
rect 58800 641800 59000 642100
rect 59300 641800 59500 642100
rect 59800 641800 60000 642100
rect 60300 641800 60500 642100
rect 60800 641800 61000 642100
rect 61300 641800 61500 642100
rect 61800 641800 62200 642100
rect 57800 641600 62200 641800
rect 57800 641300 58000 641600
rect 58300 641300 58500 641600
rect 58800 641300 59000 641600
rect 59300 641300 59500 641600
rect 59800 641300 60000 641600
rect 60300 641300 60500 641600
rect 60800 641300 61000 641600
rect 61300 641300 61500 641600
rect 61800 641300 62200 641600
rect 57800 641100 62200 641300
rect 57800 640800 58000 641100
rect 58300 640800 58500 641100
rect 58800 640800 59000 641100
rect 59300 640800 59500 641100
rect 59800 640800 60000 641100
rect 60300 640800 60500 641100
rect 60800 640800 61000 641100
rect 61300 640800 61500 641100
rect 61800 640800 62200 641100
rect 57800 640600 62200 640800
rect 57800 640300 58000 640600
rect 58300 640300 58500 640600
rect 58800 640300 59000 640600
rect 59300 640300 59500 640600
rect 59800 640300 60000 640600
rect 60300 640300 60500 640600
rect 60800 640300 61000 640600
rect 61300 640300 61500 640600
rect 61800 640300 62200 640600
rect 57800 640100 62200 640300
rect 57800 639800 58000 640100
rect 58300 639800 58500 640100
rect 58800 639800 59000 640100
rect 59300 639800 59500 640100
rect 59800 639800 60000 640100
rect 60300 639800 60500 640100
rect 60800 639800 61000 640100
rect 61300 639800 61500 640100
rect 61800 639800 62200 640100
rect 57800 639600 62200 639800
rect 57800 639300 58000 639600
rect 58300 639300 58500 639600
rect 58800 639300 59000 639600
rect 59300 639300 59500 639600
rect 59800 639300 60000 639600
rect 60300 639300 60500 639600
rect 60800 639300 61000 639600
rect 61300 639300 61500 639600
rect 61800 639300 62200 639600
rect 57800 639100 62200 639300
rect 57800 638800 58000 639100
rect 58300 638800 58500 639100
rect 58800 638800 59000 639100
rect 59300 638800 59500 639100
rect 59800 638800 60000 639100
rect 60300 638800 60500 639100
rect 60800 638800 61000 639100
rect 61300 638800 61500 639100
rect 61800 638800 62200 639100
rect 57800 638600 62200 638800
rect 57800 638300 58000 638600
rect 58300 638300 58500 638600
rect 58800 638300 59000 638600
rect 59300 638300 59500 638600
rect 59800 638300 60000 638600
rect 60300 638300 60500 638600
rect 60800 638300 61000 638600
rect 61300 638300 61500 638600
rect 61800 638300 62200 638600
rect 57800 638100 62200 638300
rect 57800 637800 58000 638100
rect 58300 637800 58500 638100
rect 58800 637800 59000 638100
rect 59300 637800 59500 638100
rect 59800 637800 60000 638100
rect 60300 637800 60500 638100
rect 60800 637800 61000 638100
rect 61300 637800 61500 638100
rect 61800 637800 62200 638100
rect 57800 637600 62200 637800
rect 57800 637300 58000 637600
rect 58300 637300 58500 637600
rect 58800 637300 59000 637600
rect 59300 637300 59500 637600
rect 59800 637300 60000 637600
rect 60300 637300 60500 637600
rect 60800 637300 61000 637600
rect 61300 637300 61500 637600
rect 61800 637300 62200 637600
rect 57800 637100 62200 637300
rect 57800 636800 58000 637100
rect 58300 636800 58500 637100
rect 58800 636800 59000 637100
rect 59300 636800 59500 637100
rect 59800 636800 60000 637100
rect 60300 636800 60500 637100
rect 60800 636800 61000 637100
rect 61300 636800 61500 637100
rect 61800 636800 62200 637100
rect 57800 636600 62200 636800
rect 57800 636300 58000 636600
rect 58300 636300 58500 636600
rect 58800 636300 59000 636600
rect 59300 636300 59500 636600
rect 59800 636300 60000 636600
rect 60300 636300 60500 636600
rect 60800 636300 61000 636600
rect 61300 636300 61500 636600
rect 61800 636300 62200 636600
rect 57800 636100 62200 636300
rect 57800 635800 58000 636100
rect 58300 635800 58500 636100
rect 58800 635800 59000 636100
rect 59300 635800 59500 636100
rect 59800 635800 60000 636100
rect 60300 635800 60500 636100
rect 60800 635800 61000 636100
rect 61300 635800 61500 636100
rect 61800 635800 62200 636100
rect 57800 635600 62200 635800
rect 57800 635300 58000 635600
rect 58300 635300 58500 635600
rect 58800 635300 59000 635600
rect 59300 635300 59500 635600
rect 59800 635300 60000 635600
rect 60300 635300 60500 635600
rect 60800 635300 61000 635600
rect 61300 635300 61500 635600
rect 61800 635300 62200 635600
rect 57800 635100 62200 635300
rect 57800 634800 58000 635100
rect 58300 634800 58500 635100
rect 58800 634800 59000 635100
rect 59300 634800 59500 635100
rect 59800 634800 60000 635100
rect 60300 634800 60500 635100
rect 60800 634800 61000 635100
rect 61300 634800 61500 635100
rect 61800 634800 62200 635100
rect 57800 634600 62200 634800
rect 57800 634300 58000 634600
rect 58300 634300 58500 634600
rect 58800 634300 59000 634600
rect 59300 634300 59500 634600
rect 59800 634300 60000 634600
rect 60300 634300 60500 634600
rect 60800 634300 61000 634600
rect 61300 634300 61500 634600
rect 61800 634300 62200 634600
rect 57800 633800 62200 634300
rect 549700 644600 553100 680800
rect 549700 644400 550000 644600
rect 550200 644400 550400 644600
rect 550600 644400 550800 644600
rect 551000 644400 551200 644600
rect 551400 644400 551600 644600
rect 551800 644400 552000 644600
rect 552200 644400 552400 644600
rect 552600 644400 552800 644600
rect 553000 644400 553100 644600
rect 549700 644200 553100 644400
rect 549700 644000 550000 644200
rect 550200 644000 550400 644200
rect 550600 644000 550800 644200
rect 551000 644000 551200 644200
rect 551400 644000 551600 644200
rect 551800 644000 552000 644200
rect 552200 644000 552400 644200
rect 552600 644000 552800 644200
rect 553000 644000 553100 644200
rect 549700 643800 553100 644000
rect 549700 643600 550000 643800
rect 550200 643600 550400 643800
rect 550600 643600 550800 643800
rect 551000 643600 551200 643800
rect 551400 643600 551600 643800
rect 551800 643600 552000 643800
rect 552200 643600 552400 643800
rect 552600 643600 552800 643800
rect 553000 643600 553100 643800
rect 549700 643400 553100 643600
rect 549700 643200 550000 643400
rect 550200 643200 550400 643400
rect 550600 643200 550800 643400
rect 551000 643200 551200 643400
rect 551400 643200 551600 643400
rect 551800 643200 552000 643400
rect 552200 643200 552400 643400
rect 552600 643200 552800 643400
rect 553000 643200 553100 643400
rect 549700 643000 553100 643200
rect 549700 642800 550000 643000
rect 550200 642800 550400 643000
rect 550600 642800 550800 643000
rect 551000 642800 551200 643000
rect 551400 642800 551600 643000
rect 551800 642800 552000 643000
rect 552200 642800 552400 643000
rect 552600 642800 552800 643000
rect 553000 642800 553100 643000
rect 549700 642600 553100 642800
rect 549700 642400 550000 642600
rect 550200 642400 550400 642600
rect 550600 642400 550800 642600
rect 551000 642400 551200 642600
rect 551400 642400 551600 642600
rect 551800 642400 552000 642600
rect 552200 642400 552400 642600
rect 552600 642400 552800 642600
rect 553000 642400 553100 642600
rect 549700 642200 553100 642400
rect 549700 642000 550000 642200
rect 550200 642000 550400 642200
rect 550600 642000 550800 642200
rect 551000 642000 551200 642200
rect 551400 642000 551600 642200
rect 551800 642000 552000 642200
rect 552200 642000 552400 642200
rect 552600 642000 552800 642200
rect 553000 642000 553100 642200
rect 549700 641800 553100 642000
rect 549700 641600 550000 641800
rect 550200 641600 550400 641800
rect 550600 641600 550800 641800
rect 551000 641600 551200 641800
rect 551400 641600 551600 641800
rect 551800 641600 552000 641800
rect 552200 641600 552400 641800
rect 552600 641600 552800 641800
rect 553000 641600 553100 641800
rect 549700 641400 553100 641600
rect 549700 641200 550000 641400
rect 550200 641200 550400 641400
rect 550600 641200 550800 641400
rect 551000 641200 551200 641400
rect 551400 641200 551600 641400
rect 551800 641200 552000 641400
rect 552200 641200 552400 641400
rect 552600 641200 552800 641400
rect 553000 641200 553100 641400
rect 549700 641000 553100 641200
rect 549700 640800 550000 641000
rect 550200 640800 550400 641000
rect 550600 640800 550800 641000
rect 551000 640800 551200 641000
rect 551400 640800 551600 641000
rect 551800 640800 552000 641000
rect 552200 640800 552400 641000
rect 552600 640800 552800 641000
rect 553000 640800 553100 641000
rect 549700 640600 553100 640800
rect 549700 640400 550000 640600
rect 550200 640400 550400 640600
rect 550600 640400 550800 640600
rect 551000 640400 551200 640600
rect 551400 640400 551600 640600
rect 551800 640400 552000 640600
rect 552200 640400 552400 640600
rect 552600 640400 552800 640600
rect 553000 640400 553100 640600
rect 549700 640200 553100 640400
rect 549700 640000 550000 640200
rect 550200 640000 550400 640200
rect 550600 640000 550800 640200
rect 551000 640000 551200 640200
rect 551400 640000 551600 640200
rect 551800 640000 552000 640200
rect 552200 640000 552400 640200
rect 552600 640000 552800 640200
rect 553000 640000 553100 640200
rect 549700 639800 553100 640000
rect 549700 639600 550000 639800
rect 550200 639600 550400 639800
rect 550600 639600 550800 639800
rect 551000 639600 551200 639800
rect 551400 639600 551600 639800
rect 551800 639600 552000 639800
rect 552200 639600 552400 639800
rect 552600 639600 552800 639800
rect 553000 639600 553100 639800
rect 549700 639400 553100 639600
rect 549700 639200 550000 639400
rect 550200 639200 550400 639400
rect 550600 639200 550800 639400
rect 551000 639200 551200 639400
rect 551400 639200 551600 639400
rect 551800 639200 552000 639400
rect 552200 639200 552400 639400
rect 552600 639200 552800 639400
rect 553000 639200 553100 639400
rect 549700 639000 553100 639200
rect 549700 638800 550000 639000
rect 550200 638800 550400 639000
rect 550600 638800 550800 639000
rect 551000 638800 551200 639000
rect 551400 638800 551600 639000
rect 551800 638800 552000 639000
rect 552200 638800 552400 639000
rect 552600 638800 552800 639000
rect 553000 638800 553100 639000
rect 549700 638600 553100 638800
rect 549700 638400 550000 638600
rect 550200 638400 550400 638600
rect 550600 638400 550800 638600
rect 551000 638400 551200 638600
rect 551400 638400 551600 638600
rect 551800 638400 552000 638600
rect 552200 638400 552400 638600
rect 552600 638400 552800 638600
rect 553000 638400 553100 638600
rect 549700 638200 553100 638400
rect 549700 638000 550000 638200
rect 550200 638000 550400 638200
rect 550600 638000 550800 638200
rect 551000 638000 551200 638200
rect 551400 638000 551600 638200
rect 551800 638000 552000 638200
rect 552200 638000 552400 638200
rect 552600 638000 552800 638200
rect 553000 638000 553100 638200
rect 549700 637800 553100 638000
rect 549700 637600 550000 637800
rect 550200 637600 550400 637800
rect 550600 637600 550800 637800
rect 551000 637600 551200 637800
rect 551400 637600 551600 637800
rect 551800 637600 552000 637800
rect 552200 637600 552400 637800
rect 552600 637600 552800 637800
rect 553000 637600 553100 637800
rect 549700 637400 553100 637600
rect 549700 637200 550000 637400
rect 550200 637200 550400 637400
rect 550600 637200 550800 637400
rect 551000 637200 551200 637400
rect 551400 637200 551600 637400
rect 551800 637200 552000 637400
rect 552200 637200 552400 637400
rect 552600 637200 552800 637400
rect 553000 637200 553100 637400
rect 549700 637000 553100 637200
rect 549700 636800 550000 637000
rect 550200 636800 550400 637000
rect 550600 636800 550800 637000
rect 551000 636800 551200 637000
rect 551400 636800 551600 637000
rect 551800 636800 552000 637000
rect 552200 636800 552400 637000
rect 552600 636800 552800 637000
rect 553000 636800 553100 637000
rect 549700 636600 553100 636800
rect 549700 636400 550000 636600
rect 550200 636400 550400 636600
rect 550600 636400 550800 636600
rect 551000 636400 551200 636600
rect 551400 636400 551600 636600
rect 551800 636400 552000 636600
rect 552200 636400 552400 636600
rect 552600 636400 552800 636600
rect 553000 636400 553100 636600
rect 549700 636200 553100 636400
rect 549700 636000 550000 636200
rect 550200 636000 550400 636200
rect 550600 636000 550800 636200
rect 551000 636000 551200 636200
rect 551400 636000 551600 636200
rect 551800 636000 552000 636200
rect 552200 636000 552400 636200
rect 552600 636000 552800 636200
rect 553000 636000 553100 636200
rect 549700 635800 553100 636000
rect 549700 635600 550000 635800
rect 550200 635600 550400 635800
rect 550600 635600 550800 635800
rect 551000 635600 551200 635800
rect 551400 635600 551600 635800
rect 551800 635600 552000 635800
rect 552200 635600 552400 635800
rect 552600 635600 552800 635800
rect 553000 635600 553100 635800
rect 549700 635400 553100 635600
rect 549700 635200 550000 635400
rect 550200 635200 550400 635400
rect 550600 635200 550800 635400
rect 551000 635200 551200 635400
rect 551400 635200 551600 635400
rect 551800 635200 552000 635400
rect 552200 635200 552400 635400
rect 552600 635200 552800 635400
rect 553000 635200 553100 635400
rect 549700 635000 553100 635200
rect 549700 634800 550000 635000
rect 550200 634800 550400 635000
rect 550600 634800 550800 635000
rect 551000 634800 551200 635000
rect 551400 634800 551600 635000
rect 551800 634800 552000 635000
rect 552200 634800 552400 635000
rect 552600 634800 552800 635000
rect 553000 634800 553100 635000
rect 549700 634600 553100 634800
rect 549700 634400 550000 634600
rect 550200 634400 550400 634600
rect 550600 634400 550800 634600
rect 551000 634400 551200 634600
rect 551400 634400 551600 634600
rect 551800 634400 552000 634600
rect 552200 634400 552400 634600
rect 552600 634400 552800 634600
rect 553000 634400 553100 634600
rect 549700 634200 553100 634400
rect 549700 634000 550000 634200
rect 550200 634000 550400 634200
rect 550600 634000 550800 634200
rect 551000 634000 551200 634200
rect 551400 634000 551600 634200
rect 551800 634000 552000 634200
rect 552200 634000 552400 634200
rect 552600 634000 552800 634200
rect 553000 634000 553100 634200
rect 549700 633800 553100 634000
rect 549700 633600 550000 633800
rect 550200 633600 550400 633800
rect 550600 633600 550800 633800
rect 551000 633600 551200 633800
rect 551400 633600 551600 633800
rect 551800 633600 552000 633800
rect 552200 633600 552400 633800
rect 552600 633600 552800 633800
rect 553000 633600 553100 633800
rect 549700 633400 553100 633600
rect 549700 633200 550000 633400
rect 550200 633200 550400 633400
rect 550600 633200 550800 633400
rect 551000 633200 551200 633400
rect 551400 633200 551600 633400
rect 551800 633200 552000 633400
rect 552200 633200 552400 633400
rect 552600 633200 552800 633400
rect 553000 633200 553100 633400
rect 549700 633000 553100 633200
rect 549700 632800 550000 633000
rect 550200 632800 550400 633000
rect 550600 632800 550800 633000
rect 551000 632800 551200 633000
rect 551400 632800 551600 633000
rect 551800 632800 552000 633000
rect 552200 632800 552400 633000
rect 552600 632800 552800 633000
rect 553000 632800 553100 633000
rect 549700 632600 553100 632800
rect 549700 632400 550000 632600
rect 550200 632400 550400 632600
rect 550600 632400 550800 632600
rect 551000 632400 551200 632600
rect 551400 632400 551600 632600
rect 551800 632400 552000 632600
rect 552200 632400 552400 632600
rect 552600 632400 552800 632600
rect 553000 632400 553100 632600
rect 549700 632200 553100 632400
rect 549700 632000 550000 632200
rect 550200 632000 550400 632200
rect 550600 632000 550800 632200
rect 551000 632000 551200 632200
rect 551400 632000 551600 632200
rect 551800 632000 552000 632200
rect 552200 632000 552400 632200
rect 552600 632000 552800 632200
rect 553000 632000 553100 632200
rect 549700 631800 553100 632000
rect 549700 631600 550000 631800
rect 550200 631600 550400 631800
rect 550600 631600 550800 631800
rect 551000 631600 551200 631800
rect 551400 631600 551600 631800
rect 551800 631600 552000 631800
rect 552200 631600 552400 631800
rect 552600 631600 552800 631800
rect 553000 631600 553100 631800
rect 549700 631400 553100 631600
rect 549700 631200 550000 631400
rect 550200 631200 550400 631400
rect 550600 631200 550800 631400
rect 551000 631200 551200 631400
rect 551400 631200 551600 631400
rect 551800 631200 552000 631400
rect 552200 631200 552400 631400
rect 552600 631200 552800 631400
rect 553000 631200 553100 631400
rect 549700 631000 553100 631200
rect 549700 630800 550000 631000
rect 550200 630800 550400 631000
rect 550600 630800 550800 631000
rect 551000 630800 551200 631000
rect 551400 630800 551600 631000
rect 551800 630800 552000 631000
rect 552200 630800 552400 631000
rect 552600 630800 552800 631000
rect 553000 630800 553100 631000
rect 549700 630700 553100 630800
rect 549700 630500 550000 630700
rect 550200 630500 550400 630700
rect 550600 630500 550800 630700
rect 551000 630500 551200 630700
rect 551400 630500 551600 630700
rect 551800 630500 552000 630700
rect 552200 630500 552400 630700
rect 552600 630500 552800 630700
rect 553000 630500 553100 630700
rect 549700 630400 553100 630500
rect 549700 630200 550000 630400
rect 550200 630200 550400 630400
rect 550600 630200 550800 630400
rect 551000 630200 551200 630400
rect 551400 630200 551600 630400
rect 551800 630200 552000 630400
rect 552200 630200 552400 630400
rect 552600 630200 552800 630400
rect 553000 630200 553100 630400
rect 549700 630000 553100 630200
rect 549700 629800 550000 630000
rect 550200 629800 550400 630000
rect 550600 629800 550800 630000
rect 551000 629800 551200 630000
rect 551400 629800 551600 630000
rect 551800 629800 552000 630000
rect 552200 629800 552400 630000
rect 552600 629800 552800 630000
rect 553000 629800 553100 630000
rect 549700 629700 553100 629800
rect 32600 563900 32800 564100
rect 33000 563900 33200 564100
rect 33400 563900 33600 564100
rect 33800 563900 34000 564100
rect 34200 563900 34400 564100
rect 34600 563900 34800 564100
rect 35000 563900 35200 564100
rect 35400 563900 35600 564100
rect 35800 563900 36000 564100
rect 36200 563900 36400 564100
rect 36600 563900 36800 564100
rect 37000 563900 37200 564100
rect 37400 563900 37600 564100
rect 37800 563900 38000 564100
rect 38200 563900 38400 564100
rect 38600 563900 38800 564100
rect 39000 563900 39200 564100
rect 39400 563900 39600 564100
rect 39800 563900 40000 564100
rect 40200 563900 40400 564100
rect 40600 563900 40800 564100
rect 32600 563700 40800 563900
rect 32600 563500 32800 563700
rect 33000 563500 33200 563700
rect 33400 563500 33600 563700
rect 33800 563500 34000 563700
rect 34200 563500 34400 563700
rect 34600 563500 34800 563700
rect 35000 563500 35200 563700
rect 35400 563500 35600 563700
rect 35800 563500 36000 563700
rect 36200 563500 36400 563700
rect 36600 563500 36800 563700
rect 37000 563500 37200 563700
rect 37400 563500 37600 563700
rect 37800 563500 38000 563700
rect 38200 563500 38400 563700
rect 38600 563500 38800 563700
rect 39000 563500 39200 563700
rect 39400 563500 39600 563700
rect 39800 563500 40000 563700
rect 40200 563500 40400 563700
rect 40600 563500 40800 563700
rect 32600 563300 40800 563500
rect 32600 563100 32800 563300
rect 33000 563100 33200 563300
rect 33400 563100 33600 563300
rect 33800 563100 34000 563300
rect 34200 563100 34400 563300
rect 34600 563100 34800 563300
rect 35000 563100 35200 563300
rect 35400 563100 35600 563300
rect 35800 563100 36000 563300
rect 36200 563100 36400 563300
rect 36600 563100 36800 563300
rect 37000 563100 37200 563300
rect 37400 563100 37600 563300
rect 37800 563100 38000 563300
rect 38200 563100 38400 563300
rect 38600 563100 38800 563300
rect 39000 563100 39200 563300
rect 39400 563100 39600 563300
rect 39800 563100 40000 563300
rect 40200 563100 40400 563300
rect 40600 563100 40800 563300
rect 32600 562900 40800 563100
rect 32600 562700 32800 562900
rect 33000 562700 33200 562900
rect 33400 562700 33600 562900
rect 33800 562700 34000 562900
rect 34200 562700 34400 562900
rect 34600 562700 34800 562900
rect 35000 562700 35200 562900
rect 35400 562700 35600 562900
rect 35800 562700 36000 562900
rect 36200 562700 36400 562900
rect 36600 562700 36800 562900
rect 37000 562700 37200 562900
rect 37400 562700 37600 562900
rect 37800 562700 38000 562900
rect 38200 562700 38400 562900
rect 38600 562700 38800 562900
rect 39000 562700 39200 562900
rect 39400 562700 39600 562900
rect 39800 562700 40000 562900
rect 40200 562700 40400 562900
rect 40600 562700 40800 562900
rect 32600 562500 40800 562700
rect 32600 562300 32800 562500
rect 33000 562300 33200 562500
rect 33400 562300 33600 562500
rect 33800 562300 34000 562500
rect 34200 562300 34400 562500
rect 34600 562300 34800 562500
rect 35000 562300 35200 562500
rect 35400 562300 35600 562500
rect 35800 562300 36000 562500
rect 36200 562300 36400 562500
rect 36600 562300 36800 562500
rect 37000 562300 37200 562500
rect 37400 562300 37600 562500
rect 37800 562300 38000 562500
rect 38200 562300 38400 562500
rect 38600 562300 38800 562500
rect 39000 562300 39200 562500
rect 39400 562300 39600 562500
rect 39800 562300 40000 562500
rect 40200 562300 40400 562500
rect 40600 562300 40800 562500
rect 32600 562100 40800 562300
rect 32600 561900 32800 562100
rect 33000 561900 33200 562100
rect 33400 561900 33600 562100
rect 33800 561900 34000 562100
rect 34200 561900 34400 562100
rect 34600 561900 34800 562100
rect 35000 561900 35200 562100
rect 35400 561900 35600 562100
rect 35800 561900 36000 562100
rect 36200 561900 36400 562100
rect 36600 561900 36800 562100
rect 37000 561900 37200 562100
rect 37400 561900 37600 562100
rect 37800 561900 38000 562100
rect 38200 561900 38400 562100
rect 38600 561900 38800 562100
rect 39000 561900 39200 562100
rect 39400 561900 39600 562100
rect 39800 561900 40000 562100
rect 40200 561900 40400 562100
rect 40600 561900 40800 562100
rect 32600 561700 40800 561900
rect 32600 561500 32800 561700
rect 33000 561500 33200 561700
rect 33400 561500 33600 561700
rect 33800 561500 34000 561700
rect 34200 561500 34400 561700
rect 34600 561500 34800 561700
rect 35000 561500 35200 561700
rect 35400 561500 35600 561700
rect 35800 561500 36000 561700
rect 36200 561500 36400 561700
rect 36600 561500 36800 561700
rect 37000 561500 37200 561700
rect 37400 561500 37600 561700
rect 37800 561500 38000 561700
rect 38200 561500 38400 561700
rect 38600 561500 38800 561700
rect 39000 561500 39200 561700
rect 39400 561500 39600 561700
rect 39800 561500 40000 561700
rect 40200 561500 40400 561700
rect 40600 561500 40800 561700
rect 32600 561300 40800 561500
rect 32600 561100 32800 561300
rect 33000 561100 33200 561300
rect 33400 561100 33600 561300
rect 33800 561100 34000 561300
rect 34200 561100 34400 561300
rect 34600 561100 34800 561300
rect 35000 561100 35200 561300
rect 35400 561100 35600 561300
rect 35800 561100 36000 561300
rect 36200 561100 36400 561300
rect 36600 561100 36800 561300
rect 37000 561100 37200 561300
rect 37400 561100 37600 561300
rect 37800 561100 38000 561300
rect 38200 561100 38400 561300
rect 38600 561100 38800 561300
rect 39000 561100 39200 561300
rect 39400 561100 39600 561300
rect 39800 561100 40000 561300
rect 40200 561100 40400 561300
rect 40600 561100 40800 561300
rect 32600 560900 40800 561100
rect 32600 560700 32800 560900
rect 33000 560700 33200 560900
rect 33400 560700 33600 560900
rect 33800 560700 34000 560900
rect 34200 560700 34400 560900
rect 34600 560700 34800 560900
rect 35000 560700 35200 560900
rect 35400 560700 35600 560900
rect 35800 560700 36000 560900
rect 36200 560700 36400 560900
rect 36600 560700 36800 560900
rect 37000 560700 37200 560900
rect 37400 560700 37600 560900
rect 37800 560700 38000 560900
rect 38200 560700 38400 560900
rect 38600 560700 38800 560900
rect 39000 560700 39200 560900
rect 39400 560700 39600 560900
rect 39800 560700 40000 560900
rect 40200 560700 40400 560900
rect 40600 560700 40800 560900
rect 32600 560500 40800 560700
rect 32600 560300 32800 560500
rect 33000 560300 33200 560500
rect 33400 560300 33600 560500
rect 33800 560300 34000 560500
rect 34200 560300 34400 560500
rect 34600 560300 34800 560500
rect 35000 560300 35200 560500
rect 35400 560300 35600 560500
rect 35800 560300 36000 560500
rect 36200 560300 36400 560500
rect 36600 560300 36800 560500
rect 37000 560300 37200 560500
rect 37400 560300 37600 560500
rect 37800 560300 38000 560500
rect 38200 560300 38400 560500
rect 38600 560300 38800 560500
rect 39000 560300 39200 560500
rect 39400 560300 39600 560500
rect 39800 560300 40000 560500
rect 40200 560300 40400 560500
rect 40600 560300 40800 560500
rect 32600 560100 40800 560300
rect 32600 559900 32800 560100
rect 33000 559900 33200 560100
rect 33400 559900 33600 560100
rect 33800 559900 34000 560100
rect 34200 559900 34400 560100
rect 34600 559900 34800 560100
rect 35000 559900 35200 560100
rect 35400 559900 35600 560100
rect 35800 559900 36000 560100
rect 36200 559900 36400 560100
rect 36600 559900 36800 560100
rect 37000 559900 37200 560100
rect 37400 559900 37600 560100
rect 37800 559900 38000 560100
rect 38200 559900 38400 560100
rect 38600 559900 38800 560100
rect 39000 559900 39200 560100
rect 39400 559900 39600 560100
rect 39800 559900 40000 560100
rect 40200 559900 40400 560100
rect 40600 559900 40800 560100
rect 32600 559700 40800 559900
rect 32600 559500 32800 559700
rect 33000 559500 33200 559700
rect 33400 559500 33600 559700
rect 33800 559500 34000 559700
rect 34200 559500 34400 559700
rect 34600 559500 34800 559700
rect 35000 559500 35200 559700
rect 35400 559500 35600 559700
rect 35800 559500 36000 559700
rect 36200 559500 36400 559700
rect 36600 559500 36800 559700
rect 37000 559500 37200 559700
rect 37400 559500 37600 559700
rect 37800 559500 38000 559700
rect 38200 559500 38400 559700
rect 38600 559500 38800 559700
rect 39000 559500 39200 559700
rect 39400 559500 39600 559700
rect 39800 559500 40000 559700
rect 40200 559500 40400 559700
rect 40600 559500 40800 559700
rect 32600 559300 40800 559500
rect 32600 559100 32800 559300
rect 33000 559100 33200 559300
rect 33400 559100 33600 559300
rect 33800 559100 34000 559300
rect 34200 559100 34400 559300
rect 34600 559100 34800 559300
rect 35000 559100 35200 559300
rect 35400 559100 35600 559300
rect 35800 559100 36000 559300
rect 36200 559100 36400 559300
rect 36600 559100 36800 559300
rect 37000 559100 37200 559300
rect 37400 559100 37600 559300
rect 37800 559100 38000 559300
rect 38200 559100 38400 559300
rect 38600 559100 38800 559300
rect 39000 559100 39200 559300
rect 39400 559100 39600 559300
rect 39800 559100 40000 559300
rect 40200 559100 40400 559300
rect 40600 559100 40800 559300
rect 32600 558900 40800 559100
rect 32600 558700 32800 558900
rect 33000 558700 33200 558900
rect 33400 558700 33600 558900
rect 33800 558700 34000 558900
rect 34200 558700 34400 558900
rect 34600 558700 34800 558900
rect 35000 558700 35200 558900
rect 35400 558700 35600 558900
rect 35800 558700 36000 558900
rect 36200 558700 36400 558900
rect 36600 558700 36800 558900
rect 37000 558700 37200 558900
rect 37400 558700 37600 558900
rect 37800 558700 38000 558900
rect 38200 558700 38400 558900
rect 38600 558700 38800 558900
rect 39000 558700 39200 558900
rect 39400 558700 39600 558900
rect 39800 558700 40000 558900
rect 40200 558700 40400 558900
rect 40600 558700 40800 558900
rect 32600 558500 40800 558700
rect 32600 558300 32800 558500
rect 33000 558300 33200 558500
rect 33400 558300 33600 558500
rect 33800 558300 34000 558500
rect 34200 558300 34400 558500
rect 34600 558300 34800 558500
rect 35000 558300 35200 558500
rect 35400 558300 35600 558500
rect 35800 558300 36000 558500
rect 36200 558300 36400 558500
rect 36600 558300 36800 558500
rect 37000 558300 37200 558500
rect 37400 558300 37600 558500
rect 37800 558300 38000 558500
rect 38200 558300 38400 558500
rect 38600 558300 38800 558500
rect 39000 558300 39200 558500
rect 39400 558300 39600 558500
rect 39800 558300 40000 558500
rect 40200 558300 40400 558500
rect 40600 558300 40800 558500
rect 32600 558100 40800 558300
rect 32600 557900 32800 558100
rect 33000 557900 33200 558100
rect 33400 557900 33600 558100
rect 33800 557900 34000 558100
rect 34200 557900 34400 558100
rect 34600 557900 34800 558100
rect 35000 557900 35200 558100
rect 35400 557900 35600 558100
rect 35800 557900 36000 558100
rect 36200 557900 36400 558100
rect 36600 557900 36800 558100
rect 37000 557900 37200 558100
rect 37400 557900 37600 558100
rect 37800 557900 38000 558100
rect 38200 557900 38400 558100
rect 38600 557900 38800 558100
rect 39000 557900 39200 558100
rect 39400 557900 39600 558100
rect 39800 557900 40000 558100
rect 40200 557900 40400 558100
rect 40600 557900 40800 558100
rect 32600 557700 40800 557900
rect 32600 557500 32800 557700
rect 33000 557500 33200 557700
rect 33400 557500 33600 557700
rect 33800 557500 34000 557700
rect 34200 557500 34400 557700
rect 34600 557500 34800 557700
rect 35000 557500 35200 557700
rect 35400 557500 35600 557700
rect 35800 557500 36000 557700
rect 36200 557500 36400 557700
rect 36600 557500 36800 557700
rect 37000 557500 37200 557700
rect 37400 557500 37600 557700
rect 37800 557500 38000 557700
rect 38200 557500 38400 557700
rect 38600 557500 38800 557700
rect 39000 557500 39200 557700
rect 39400 557500 39600 557700
rect 39800 557500 40000 557700
rect 40200 557500 40400 557700
rect 40600 557500 40800 557700
rect 32600 557300 40800 557500
rect 32600 557100 32800 557300
rect 33000 557100 33200 557300
rect 33400 557100 33600 557300
rect 33800 557100 34000 557300
rect 34200 557100 34400 557300
rect 34600 557100 34800 557300
rect 35000 557100 35200 557300
rect 35400 557100 35600 557300
rect 35800 557100 36000 557300
rect 36200 557100 36400 557300
rect 36600 557100 36800 557300
rect 37000 557100 37200 557300
rect 37400 557100 37600 557300
rect 37800 557100 38000 557300
rect 38200 557100 38400 557300
rect 38600 557100 38800 557300
rect 39000 557100 39200 557300
rect 39400 557100 39600 557300
rect 39800 557100 40000 557300
rect 40200 557100 40400 557300
rect 40600 557100 40800 557300
rect 32600 556900 40800 557100
rect 32600 556700 32800 556900
rect 33000 556700 33200 556900
rect 33400 556700 33600 556900
rect 33800 556700 34000 556900
rect 34200 556700 34400 556900
rect 34600 556700 34800 556900
rect 35000 556700 35200 556900
rect 35400 556700 35600 556900
rect 35800 556700 36000 556900
rect 36200 556700 36400 556900
rect 36600 556700 36800 556900
rect 37000 556700 37200 556900
rect 37400 556700 37600 556900
rect 37800 556700 38000 556900
rect 38200 556700 38400 556900
rect 38600 556700 38800 556900
rect 39000 556700 39200 556900
rect 39400 556700 39600 556900
rect 39800 556700 40000 556900
rect 40200 556700 40400 556900
rect 40600 556700 40800 556900
rect 32600 556500 40800 556700
rect 32600 556300 32800 556500
rect 33000 556300 33200 556500
rect 33400 556300 33600 556500
rect 33800 556300 34000 556500
rect 34200 556300 34400 556500
rect 34600 556300 34800 556500
rect 35000 556300 35200 556500
rect 35400 556300 35600 556500
rect 35800 556300 36000 556500
rect 36200 556300 36400 556500
rect 36600 556300 36800 556500
rect 37000 556300 37200 556500
rect 37400 556300 37600 556500
rect 37800 556300 38000 556500
rect 38200 556300 38400 556500
rect 38600 556300 38800 556500
rect 39000 556300 39200 556500
rect 39400 556300 39600 556500
rect 39800 556300 40000 556500
rect 40200 556300 40400 556500
rect 40600 556300 40800 556500
rect 32600 556100 40800 556300
rect 32600 555900 32800 556100
rect 33000 555900 33200 556100
rect 33400 555900 33600 556100
rect 33800 555900 34000 556100
rect 34200 555900 34400 556100
rect 34600 555900 34800 556100
rect 35000 555900 35200 556100
rect 35400 555900 35600 556100
rect 35800 555900 36000 556100
rect 36200 555900 36400 556100
rect 36600 555900 36800 556100
rect 37000 555900 37200 556100
rect 37400 555900 37600 556100
rect 37800 555900 38000 556100
rect 38200 555900 38400 556100
rect 38600 555900 38800 556100
rect 39000 555900 39200 556100
rect 39400 555900 39600 556100
rect 39800 555900 40000 556100
rect 40200 555900 40400 556100
rect 40600 555900 40800 556100
rect 32600 555700 40800 555900
rect 32600 555500 32800 555700
rect 33000 555500 33200 555700
rect 33400 555500 33600 555700
rect 33800 555500 34000 555700
rect 34200 555500 34400 555700
rect 34600 555500 34800 555700
rect 35000 555500 35200 555700
rect 35400 555500 35600 555700
rect 35800 555500 36000 555700
rect 36200 555500 36400 555700
rect 36600 555500 36800 555700
rect 37000 555500 37200 555700
rect 37400 555500 37600 555700
rect 37800 555500 38000 555700
rect 38200 555500 38400 555700
rect 38600 555500 38800 555700
rect 39000 555500 39200 555700
rect 39400 555500 39600 555700
rect 39800 555500 40000 555700
rect 40200 555500 40400 555700
rect 40600 555500 40800 555700
rect 32600 555300 40800 555500
rect 32600 555100 32800 555300
rect 33000 555100 33200 555300
rect 33400 555100 33600 555300
rect 33800 555100 34000 555300
rect 34200 555100 34400 555300
rect 34600 555100 34800 555300
rect 35000 555100 35200 555300
rect 35400 555100 35600 555300
rect 35800 555100 36000 555300
rect 36200 555100 36400 555300
rect 36600 555100 36800 555300
rect 37000 555100 37200 555300
rect 37400 555100 37600 555300
rect 37800 555100 38000 555300
rect 38200 555100 38400 555300
rect 38600 555100 38800 555300
rect 39000 555100 39200 555300
rect 39400 555100 39600 555300
rect 39800 555100 40000 555300
rect 40200 555100 40400 555300
rect 40600 555100 40800 555300
rect 32600 554900 40800 555100
rect 32600 554700 32800 554900
rect 33000 554700 33200 554900
rect 33400 554700 33600 554900
rect 33800 554700 34000 554900
rect 34200 554700 34400 554900
rect 34600 554700 34800 554900
rect 35000 554700 35200 554900
rect 35400 554700 35600 554900
rect 35800 554700 36000 554900
rect 36200 554700 36400 554900
rect 36600 554700 36800 554900
rect 37000 554700 37200 554900
rect 37400 554700 37600 554900
rect 37800 554700 38000 554900
rect 38200 554700 38400 554900
rect 38600 554700 38800 554900
rect 39000 554700 39200 554900
rect 39400 554700 39600 554900
rect 39800 554700 40000 554900
rect 40200 554700 40400 554900
rect 40600 554700 40800 554900
rect 32600 554500 40800 554700
rect 32600 554300 32800 554500
rect 33000 554300 33200 554500
rect 33400 554300 33600 554500
rect 33800 554300 34000 554500
rect 34200 554300 34400 554500
rect 34600 554300 34800 554500
rect 35000 554300 35200 554500
rect 35400 554300 35600 554500
rect 35800 554300 36000 554500
rect 36200 554300 36400 554500
rect 36600 554300 36800 554500
rect 37000 554300 37200 554500
rect 37400 554300 37600 554500
rect 37800 554300 38000 554500
rect 38200 554300 38400 554500
rect 38600 554300 38800 554500
rect 39000 554300 39200 554500
rect 39400 554300 39600 554500
rect 39800 554300 40000 554500
rect 40200 554300 40400 554500
rect 40600 554300 40800 554500
rect 32600 554100 40800 554300
rect 32600 553900 32800 554100
rect 33000 553900 33200 554100
rect 33400 553900 33600 554100
rect 33800 553900 34000 554100
rect 34200 553900 34400 554100
rect 34600 553900 34800 554100
rect 35000 553900 35200 554100
rect 35400 553900 35600 554100
rect 35800 553900 36000 554100
rect 36200 553900 36400 554100
rect 36600 553900 36800 554100
rect 37000 553900 37200 554100
rect 37400 553900 37600 554100
rect 37800 553900 38000 554100
rect 38200 553900 38400 554100
rect 38600 553900 38800 554100
rect 39000 553900 39200 554100
rect 39400 553900 39600 554100
rect 39800 553900 40000 554100
rect 40200 553900 40400 554100
rect 40600 553900 40800 554100
rect 32600 553700 40800 553900
rect 32600 553500 32800 553700
rect 33000 553500 33200 553700
rect 33400 553500 33600 553700
rect 33800 553500 34000 553700
rect 34200 553500 34400 553700
rect 34600 553500 34800 553700
rect 35000 553500 35200 553700
rect 35400 553500 35600 553700
rect 35800 553500 36000 553700
rect 36200 553500 36400 553700
rect 36600 553500 36800 553700
rect 37000 553500 37200 553700
rect 37400 553500 37600 553700
rect 37800 553500 38000 553700
rect 38200 553500 38400 553700
rect 38600 553500 38800 553700
rect 39000 553500 39200 553700
rect 39400 553500 39600 553700
rect 39800 553500 40000 553700
rect 40200 553500 40400 553700
rect 40600 553500 40800 553700
rect 32600 553300 40800 553500
rect 32600 553100 32800 553300
rect 33000 553100 33200 553300
rect 33400 553100 33600 553300
rect 33800 553100 34000 553300
rect 34200 553100 34400 553300
rect 34600 553100 34800 553300
rect 35000 553100 35200 553300
rect 35400 553100 35600 553300
rect 35800 553100 36000 553300
rect 36200 553100 36400 553300
rect 36600 553100 36800 553300
rect 37000 553100 37200 553300
rect 37400 553100 37600 553300
rect 37800 553100 38000 553300
rect 38200 553100 38400 553300
rect 38600 553100 38800 553300
rect 39000 553100 39200 553300
rect 39400 553100 39600 553300
rect 39800 553100 40000 553300
rect 40200 553100 40400 553300
rect 40600 553100 40800 553300
rect 32600 552900 40800 553100
rect 32600 552700 32800 552900
rect 33000 552700 33200 552900
rect 33400 552700 33600 552900
rect 33800 552700 34000 552900
rect 34200 552700 34400 552900
rect 34600 552700 34800 552900
rect 35000 552700 35200 552900
rect 35400 552700 35600 552900
rect 35800 552700 36000 552900
rect 36200 552700 36400 552900
rect 36600 552700 36800 552900
rect 37000 552700 37200 552900
rect 37400 552700 37600 552900
rect 37800 552700 38000 552900
rect 38200 552700 38400 552900
rect 38600 552700 38800 552900
rect 39000 552700 39200 552900
rect 39400 552700 39600 552900
rect 39800 552700 40000 552900
rect 40200 552700 40400 552900
rect 40600 552700 40800 552900
rect 32600 552500 40800 552700
rect 32600 552300 32800 552500
rect 33000 552300 33200 552500
rect 33400 552300 33600 552500
rect 33800 552300 34000 552500
rect 34200 552300 34400 552500
rect 34600 552300 34800 552500
rect 35000 552300 35200 552500
rect 35400 552300 35600 552500
rect 35800 552300 36000 552500
rect 36200 552300 36400 552500
rect 36600 552300 36800 552500
rect 37000 552300 37200 552500
rect 37400 552300 37600 552500
rect 37800 552300 38000 552500
rect 38200 552300 38400 552500
rect 38600 552300 38800 552500
rect 39000 552300 39200 552500
rect 39400 552300 39600 552500
rect 39800 552300 40000 552500
rect 40200 552300 40400 552500
rect 40600 552300 40800 552500
rect 32600 552100 40800 552300
rect 32600 551900 32800 552100
rect 33000 551900 33200 552100
rect 33400 551900 33600 552100
rect 33800 551900 34000 552100
rect 34200 551900 34400 552100
rect 34600 551900 34800 552100
rect 35000 551900 35200 552100
rect 35400 551900 35600 552100
rect 35800 551900 36000 552100
rect 36200 551900 36400 552100
rect 36600 551900 36800 552100
rect 37000 551900 37200 552100
rect 37400 551900 37600 552100
rect 37800 551900 38000 552100
rect 38200 551900 38400 552100
rect 38600 551900 38800 552100
rect 39000 551900 39200 552100
rect 39400 551900 39600 552100
rect 39800 551900 40000 552100
rect 40200 551900 40400 552100
rect 40600 551900 40800 552100
rect 32600 551700 40800 551900
rect 32600 551500 32800 551700
rect 33000 551500 33200 551700
rect 33400 551500 33600 551700
rect 33800 551500 34000 551700
rect 34200 551500 34400 551700
rect 34600 551500 34800 551700
rect 35000 551500 35200 551700
rect 35400 551500 35600 551700
rect 35800 551500 36000 551700
rect 36200 551500 36400 551700
rect 36600 551500 36800 551700
rect 37000 551500 37200 551700
rect 37400 551500 37600 551700
rect 37800 551500 38000 551700
rect 38200 551500 38400 551700
rect 38600 551500 38800 551700
rect 39000 551500 39200 551700
rect 39400 551500 39600 551700
rect 39800 551500 40000 551700
rect 40200 551500 40400 551700
rect 40600 551500 40800 551700
rect 32600 551300 40800 551500
rect 32600 551100 32800 551300
rect 33000 551100 33200 551300
rect 33400 551100 33600 551300
rect 33800 551100 34000 551300
rect 34200 551100 34400 551300
rect 34600 551100 34800 551300
rect 35000 551100 35200 551300
rect 35400 551100 35600 551300
rect 35800 551100 36000 551300
rect 36200 551100 36400 551300
rect 36600 551100 36800 551300
rect 37000 551100 37200 551300
rect 37400 551100 37600 551300
rect 37800 551100 38000 551300
rect 38200 551100 38400 551300
rect 38600 551100 38800 551300
rect 39000 551100 39200 551300
rect 39400 551100 39600 551300
rect 39800 551100 40000 551300
rect 40200 551100 40400 551300
rect 40600 551100 40800 551300
rect 32600 550900 40800 551100
rect 32600 550700 32800 550900
rect 33000 550700 33200 550900
rect 33400 550700 33600 550900
rect 33800 550700 34000 550900
rect 34200 550700 34400 550900
rect 34600 550700 34800 550900
rect 35000 550700 35200 550900
rect 35400 550700 35600 550900
rect 35800 550700 36000 550900
rect 36200 550700 36400 550900
rect 36600 550700 36800 550900
rect 37000 550700 37200 550900
rect 37400 550700 37600 550900
rect 37800 550700 38000 550900
rect 38200 550700 38400 550900
rect 38600 550700 38800 550900
rect 39000 550700 39200 550900
rect 39400 550700 39600 550900
rect 39800 550700 40000 550900
rect 40200 550700 40400 550900
rect 40600 550700 40800 550900
rect 32600 550500 40800 550700
rect 32600 550300 32800 550500
rect 33000 550300 33200 550500
rect 33400 550300 33600 550500
rect 33800 550300 34000 550500
rect 34200 550300 34400 550500
rect 34600 550300 34800 550500
rect 35000 550300 35200 550500
rect 35400 550300 35600 550500
rect 35800 550300 36000 550500
rect 36200 550300 36400 550500
rect 36600 550300 36800 550500
rect 37000 550300 37200 550500
rect 37400 550300 37600 550500
rect 37800 550300 38000 550500
rect 38200 550300 38400 550500
rect 38600 550300 38800 550500
rect 39000 550300 39200 550500
rect 39400 550300 39600 550500
rect 39800 550300 40000 550500
rect 40200 550300 40400 550500
rect 40600 550300 40800 550500
rect 32600 550100 40800 550300
rect 32600 549900 32800 550100
rect 33000 549900 33200 550100
rect 33400 549900 33600 550100
rect 33800 549900 34000 550100
rect 34200 549900 34400 550100
rect 34600 549900 34800 550100
rect 35000 549900 35200 550100
rect 35400 549900 35600 550100
rect 35800 549900 36000 550100
rect 36200 549900 36400 550100
rect 36600 549900 36800 550100
rect 37000 549900 37200 550100
rect 37400 549900 37600 550100
rect 37800 549900 38000 550100
rect 38200 549900 38400 550100
rect 38600 549900 38800 550100
rect 39000 549900 39200 550100
rect 39400 549900 39600 550100
rect 39800 549900 40000 550100
rect 40200 549900 40400 550100
rect 40600 549900 40800 550100
rect 32600 549700 40800 549900
rect 32600 549500 32800 549700
rect 33000 549500 33200 549700
rect 33400 549500 33600 549700
rect 33800 549500 34000 549700
rect 34200 549500 34400 549700
rect 34600 549500 34800 549700
rect 35000 549500 35200 549700
rect 35400 549500 35600 549700
rect 35800 549500 36000 549700
rect 36200 549500 36400 549700
rect 36600 549500 36800 549700
rect 37000 549500 37200 549700
rect 37400 549500 37600 549700
rect 37800 549500 38000 549700
rect 38200 549500 38400 549700
rect 38600 549500 38800 549700
rect 39000 549500 39200 549700
rect 39400 549500 39600 549700
rect 39800 549500 40000 549700
rect 40200 549500 40400 549700
rect 40600 549500 40800 549700
rect 32600 549400 40800 549500
rect 282000 583800 284000 584200
rect 282000 583400 282400 583800
rect 282800 583400 283200 583800
rect 283600 583400 284000 583800
rect 282000 583000 284000 583400
rect 282000 582600 282400 583000
rect 282800 582600 283200 583000
rect 283600 582600 284000 583000
rect 282000 582200 284000 582600
rect 282000 581800 282400 582200
rect 282800 581800 283200 582200
rect 283600 581800 284000 582200
rect 282000 581400 284000 581800
rect 282000 581000 282400 581400
rect 282800 581000 283200 581400
rect 283600 581000 284000 581400
rect 282000 580600 284000 581000
rect 282000 580200 282400 580600
rect 282800 580200 283200 580600
rect 283600 580200 284000 580600
rect 282000 579800 284000 580200
rect 282000 579400 282400 579800
rect 282800 579400 283200 579800
rect 283600 579400 284000 579800
rect 282000 354300 284000 579400
rect 285000 494200 287000 494600
rect 285000 493800 285400 494200
rect 285800 493800 286200 494200
rect 286600 493800 287000 494200
rect 285000 493400 287000 493800
rect 285000 493000 285400 493400
rect 285800 493000 286200 493400
rect 286600 493000 287000 493400
rect 285000 492600 287000 493000
rect 285000 492200 285400 492600
rect 285800 492200 286200 492600
rect 286600 492200 287000 492600
rect 285000 491800 287000 492200
rect 285000 491400 285400 491800
rect 285800 491400 286200 491800
rect 286600 491400 287000 491800
rect 285000 491000 287000 491400
rect 285000 490600 285400 491000
rect 285800 490600 286200 491000
rect 286600 490600 287000 491000
rect 285000 490200 287000 490600
rect 285000 489800 285400 490200
rect 285800 489800 286200 490200
rect 286600 489800 287000 490200
rect 285000 354900 287000 489800
rect 288000 449800 290000 450100
rect 288000 449400 288400 449800
rect 288800 449400 289200 449800
rect 289600 449400 290000 449800
rect 288000 449000 290000 449400
rect 288000 448600 288400 449000
rect 288800 448600 289200 449000
rect 289600 448600 290000 449000
rect 288000 448200 290000 448600
rect 288000 447800 288400 448200
rect 288800 447800 289200 448200
rect 289600 447800 290000 448200
rect 288000 447400 290000 447800
rect 288000 447000 288400 447400
rect 288800 447000 289200 447400
rect 289600 447000 290000 447400
rect 288000 446600 290000 447000
rect 288000 446200 288400 446600
rect 288800 446200 289200 446600
rect 289600 446200 290000 446600
rect 288000 445800 290000 446200
rect 288000 445400 288400 445800
rect 288800 445400 289200 445800
rect 289600 445400 290000 445800
rect 288000 354900 290000 445400
rect 285000 354600 287467 354900
rect 282000 354000 287067 354300
rect 286847 353870 287067 354000
rect 287247 353890 287467 354600
rect 287647 354810 290000 354900
rect 291100 405400 293100 405700
rect 291100 405000 291400 405400
rect 291800 405000 292200 405400
rect 292600 405000 293100 405400
rect 291100 404600 293100 405000
rect 291100 404200 291400 404600
rect 291800 404200 292200 404600
rect 292600 404200 293100 404600
rect 291100 403800 293100 404200
rect 291100 403400 291400 403800
rect 291800 403400 292200 403800
rect 292600 403400 293100 403800
rect 291100 403000 293100 403400
rect 291100 402600 291400 403000
rect 291800 402600 292200 403000
rect 292600 402600 293100 403000
rect 291100 402200 293100 402600
rect 291100 401800 291400 402200
rect 291800 401800 292200 402200
rect 292600 401800 293100 402200
rect 291100 401400 293100 401800
rect 291100 401000 291400 401400
rect 291800 401000 292200 401400
rect 292600 401000 293100 401400
rect 287647 354590 290010 354810
rect 287647 353700 287867 354590
rect 291100 354300 293100 401000
rect 288047 354000 293100 354300
rect 294000 359000 296000 359400
rect 294000 358600 294400 359000
rect 294800 358600 295200 359000
rect 295600 358600 296000 359000
rect 294000 358200 296000 358600
rect 294000 357800 294400 358200
rect 294800 357800 295200 358200
rect 295600 357800 296000 358200
rect 294000 357400 296000 357800
rect 294000 357000 294400 357400
rect 294800 357000 295200 357400
rect 295600 357000 296000 357400
rect 294000 356600 296000 357000
rect 294000 356200 294400 356600
rect 294800 356200 295200 356600
rect 295600 356200 296000 356600
rect 294000 355800 296000 356200
rect 294000 355400 294400 355800
rect 294800 355400 295200 355800
rect 295600 355400 296000 355800
rect 294000 355000 296000 355400
rect 294000 354600 294400 355000
rect 294800 354600 295200 355000
rect 295600 354600 296000 355000
rect 288047 353700 288267 354000
rect 294000 353500 296000 354600
rect 294173 351766 294641 353500
rect 297000 344300 306000 344600
rect 294799 344200 295101 344201
rect 294799 343900 294800 344200
rect 295100 343900 295101 344200
rect 294799 343899 295101 343900
rect 297000 343900 299000 344300
rect 299400 343900 299600 344300
rect 300000 343900 300200 344300
rect 300600 343900 300800 344300
rect 301200 343900 301400 344300
rect 301800 343900 302000 344300
rect 302400 343900 302600 344300
rect 303000 343900 303200 344300
rect 303600 343900 306000 344300
rect 297000 343700 306000 343900
rect 297000 343300 299000 343700
rect 299400 343300 299600 343700
rect 300000 343300 300200 343700
rect 300600 343300 300800 343700
rect 301200 343300 301400 343700
rect 301800 343300 302000 343700
rect 302400 343300 302600 343700
rect 303000 343300 303200 343700
rect 303600 343300 306000 343700
rect 288299 340800 288601 340801
rect 288299 340500 288300 340800
rect 288600 340500 288601 340800
rect 288299 340499 288601 340500
rect 9600 304200 11800 304400
rect 9600 304000 9800 304200
rect 10000 304000 10200 304200
rect 10400 304000 10600 304200
rect 10800 304000 11000 304200
rect 11200 304000 11400 304200
rect 11600 304000 11800 304200
rect 9600 303600 11800 304000
rect 9600 303400 9800 303600
rect 10000 303400 10200 303600
rect 10400 303400 10600 303600
rect 10800 303400 11000 303600
rect 11200 303400 11400 303600
rect 11600 303400 11800 303600
rect 9600 301200 11800 303400
rect 5700 301000 18600 301200
rect 5700 300800 5800 301000
rect 6000 300800 6200 301000
rect 6400 300800 6600 301000
rect 6800 300800 7000 301000
rect 7200 300800 7400 301000
rect 7600 300800 7800 301000
rect 8000 300800 17800 301000
rect 18000 300800 18200 301000
rect 18400 300800 18600 301000
rect 5700 300600 18600 300800
rect 5700 300400 5800 300600
rect 6000 300400 6200 300600
rect 6400 300400 6600 300600
rect 6800 300400 7000 300600
rect 7200 300400 7400 300600
rect 7600 300400 7800 300600
rect 8000 300400 17800 300600
rect 18000 300400 18200 300600
rect 18400 300400 18600 300600
rect 5700 300200 18600 300400
rect 5700 300000 5800 300200
rect 6000 300000 6200 300200
rect 6400 300000 6600 300200
rect 6800 300000 7000 300200
rect 7200 300000 7400 300200
rect 7600 300000 7800 300200
rect 8000 300000 17800 300200
rect 18000 300000 18200 300200
rect 18400 300000 18600 300200
rect 5700 299800 18600 300000
rect 5700 299600 5800 299800
rect 6000 299600 6200 299800
rect 6400 299600 6600 299800
rect 6800 299600 7000 299800
rect 7200 299600 7400 299800
rect 7600 299600 7800 299800
rect 8000 299600 17800 299800
rect 18000 299600 18200 299800
rect 18400 299600 18600 299800
rect 5700 299400 18600 299600
rect 5700 299200 5800 299400
rect 6000 299200 6200 299400
rect 6400 299200 6600 299400
rect 6800 299200 7000 299400
rect 7200 299200 7400 299400
rect 7600 299200 7800 299400
rect 8000 299200 17800 299400
rect 18000 299200 18200 299400
rect 18400 299200 18600 299400
rect 5700 299000 18600 299200
rect 5700 298800 5800 299000
rect 6000 298800 6200 299000
rect 6400 298800 6600 299000
rect 6800 298800 7000 299000
rect 7200 298800 7400 299000
rect 7600 298800 7800 299000
rect 8000 298800 17800 299000
rect 18000 298800 18200 299000
rect 18400 298800 18600 299000
rect 5700 298600 18600 298800
rect 5700 298400 5800 298600
rect 6000 298400 6200 298600
rect 6400 298400 6600 298600
rect 6800 298400 7000 298600
rect 7200 298400 7400 298600
rect 7600 298400 7800 298600
rect 8000 298400 17800 298600
rect 18000 298400 18200 298600
rect 18400 298400 18600 298600
rect 5700 298200 18600 298400
rect 5700 298000 5800 298200
rect 6000 298000 6200 298200
rect 6400 298000 6600 298200
rect 6800 298000 7000 298200
rect 7200 298000 7400 298200
rect 7600 298000 7800 298200
rect 8000 298000 17800 298200
rect 18000 298000 18200 298200
rect 18400 298000 18600 298200
rect 5700 297800 18600 298000
rect 5700 297600 5800 297800
rect 6000 297600 6200 297800
rect 6400 297600 6600 297800
rect 6800 297600 7000 297800
rect 7200 297600 7400 297800
rect 7600 297600 7800 297800
rect 8000 297600 17800 297800
rect 18000 297600 18200 297800
rect 18400 297600 18600 297800
rect 5700 297400 18600 297600
rect 5700 297200 5800 297400
rect 6000 297200 6200 297400
rect 6400 297200 6600 297400
rect 6800 297200 7000 297400
rect 7200 297200 7400 297400
rect 7600 297200 7800 297400
rect 8000 297200 17800 297400
rect 18000 297200 18200 297400
rect 18400 297200 18600 297400
rect 5700 297000 18600 297200
rect 5700 296800 5800 297000
rect 6000 296800 6200 297000
rect 6400 296800 6600 297000
rect 6800 296800 7000 297000
rect 7200 296800 7400 297000
rect 7600 296800 7800 297000
rect 8000 296800 17800 297000
rect 18000 296800 18200 297000
rect 18400 296800 18600 297000
rect 5700 296600 18600 296800
rect 5700 296400 5800 296600
rect 6000 296400 6200 296600
rect 6400 296400 6600 296600
rect 6800 296400 7000 296600
rect 7200 296400 7400 296600
rect 7600 296400 7800 296600
rect 8000 296400 17800 296600
rect 18000 296400 18200 296600
rect 18400 296400 18600 296600
rect 5700 296200 18600 296400
rect 5700 293920 5960 296200
rect 5700 293740 5740 293920
rect 5920 293740 5960 293920
rect 5700 293580 5960 293740
rect 5700 293400 5740 293580
rect 5920 293400 5960 293580
rect 5700 293240 5960 293400
rect 5700 293060 5740 293240
rect 5920 293060 5960 293240
rect 5700 293040 5960 293060
rect 9600 293800 11800 294000
rect 9600 293600 9800 293800
rect 10000 293600 10200 293800
rect 10400 293600 10600 293800
rect 10800 293600 11000 293800
rect 11200 293600 11400 293800
rect 11600 293600 11800 293800
rect 9600 293200 11800 293600
rect 9600 293000 9800 293200
rect 10000 293000 10200 293200
rect 10400 293000 10600 293200
rect 10800 293000 11000 293200
rect 11200 293000 11400 293200
rect 11600 293000 11800 293200
rect 9600 290200 11800 293000
rect 9600 289800 74200 290200
rect 9600 289600 16100 289800
rect 16300 289600 25800 289800
rect 26000 289600 59400 289800
rect 9600 289500 59400 289600
rect 59700 289500 59900 289800
rect 60200 289500 60400 289800
rect 60700 289500 60900 289800
rect 61200 289500 61400 289800
rect 61700 289500 61900 289800
rect 62200 289500 62400 289800
rect 62700 289500 62900 289800
rect 63200 289500 63400 289800
rect 63700 289500 63900 289800
rect 64200 289500 64400 289800
rect 64700 289500 64900 289800
rect 65200 289500 65400 289800
rect 65700 289500 65900 289800
rect 66200 289500 66400 289800
rect 66700 289500 66900 289800
rect 67200 289500 67400 289800
rect 67700 289500 67900 289800
rect 68200 289500 68400 289800
rect 68700 289500 68900 289800
rect 69200 289500 69400 289800
rect 69700 289500 69900 289800
rect 70200 289500 70400 289800
rect 70700 289500 70900 289800
rect 71200 289500 71400 289800
rect 71700 289500 71900 289800
rect 72200 289500 72400 289800
rect 72700 289500 72900 289800
rect 73200 289500 73400 289800
rect 73700 289500 74200 289800
rect 9600 289400 74200 289500
rect 9600 289200 16100 289400
rect 16300 289200 25800 289400
rect 26000 289300 74200 289400
rect 26000 289200 59400 289300
rect 9600 289000 59400 289200
rect 59700 289000 59900 289300
rect 60200 289000 60400 289300
rect 60700 289000 60900 289300
rect 61200 289000 61400 289300
rect 61700 289000 61900 289300
rect 62200 289000 62400 289300
rect 62700 289000 62900 289300
rect 63200 289000 63400 289300
rect 63700 289000 63900 289300
rect 64200 289000 64400 289300
rect 64700 289000 64900 289300
rect 65200 289000 65400 289300
rect 65700 289000 65900 289300
rect 66200 289000 66400 289300
rect 66700 289000 66900 289300
rect 67200 289000 67400 289300
rect 67700 289000 67900 289300
rect 68200 289000 68400 289300
rect 68700 289000 68900 289300
rect 69200 289000 69400 289300
rect 69700 289000 69900 289300
rect 70200 289000 70400 289300
rect 70700 289000 70900 289300
rect 71200 289000 71400 289300
rect 71700 289000 71900 289300
rect 72200 289000 72400 289300
rect 72700 289000 72900 289300
rect 73200 289000 73400 289300
rect 73700 289000 74200 289300
rect 9600 288800 16100 289000
rect 16300 288800 25800 289000
rect 26000 288800 74200 289000
rect 9600 288600 59400 288800
rect 9600 288400 16100 288600
rect 16300 288400 25800 288600
rect 26000 288500 59400 288600
rect 59700 288500 59900 288800
rect 60200 288500 60400 288800
rect 60700 288500 60900 288800
rect 61200 288500 61400 288800
rect 61700 288500 61900 288800
rect 62200 288500 62400 288800
rect 62700 288500 62900 288800
rect 63200 288500 63400 288800
rect 63700 288500 63900 288800
rect 64200 288500 64400 288800
rect 64700 288500 64900 288800
rect 65200 288500 65400 288800
rect 65700 288500 65900 288800
rect 66200 288500 66400 288800
rect 66700 288500 66900 288800
rect 67200 288500 67400 288800
rect 67700 288500 67900 288800
rect 68200 288500 68400 288800
rect 68700 288500 68900 288800
rect 69200 288500 69400 288800
rect 69700 288500 69900 288800
rect 70200 288500 70400 288800
rect 70700 288500 70900 288800
rect 71200 288500 71400 288800
rect 71700 288500 71900 288800
rect 72200 288500 72400 288800
rect 72700 288500 72900 288800
rect 73200 288500 73400 288800
rect 73700 288500 74200 288800
rect 26000 288400 74200 288500
rect 9600 288300 74200 288400
rect 9600 288200 59400 288300
rect 9600 288000 16100 288200
rect 16300 288000 25800 288200
rect 26000 288000 59400 288200
rect 59700 288000 59900 288300
rect 60200 288000 60400 288300
rect 60700 288000 60900 288300
rect 61200 288000 61400 288300
rect 61700 288000 61900 288300
rect 62200 288000 62400 288300
rect 62700 288000 62900 288300
rect 63200 288000 63400 288300
rect 63700 288000 63900 288300
rect 64200 288000 64400 288300
rect 64700 288000 64900 288300
rect 65200 288000 65400 288300
rect 65700 288000 65900 288300
rect 66200 288000 66400 288300
rect 66700 288000 66900 288300
rect 67200 288000 67400 288300
rect 67700 288000 67900 288300
rect 68200 288000 68400 288300
rect 68700 288000 68900 288300
rect 69200 288000 69400 288300
rect 69700 288000 69900 288300
rect 70200 288000 70400 288300
rect 70700 288000 70900 288300
rect 71200 288000 71400 288300
rect 71700 288000 71900 288300
rect 72200 288000 72400 288300
rect 72700 288000 72900 288300
rect 73200 288000 73400 288300
rect 73700 288000 74200 288300
rect 9600 287800 74200 288000
rect 9600 287600 16100 287800
rect 16300 287600 25800 287800
rect 26000 287600 59400 287800
rect 9600 287500 59400 287600
rect 59700 287500 59900 287800
rect 60200 287500 60400 287800
rect 60700 287500 60900 287800
rect 61200 287500 61400 287800
rect 61700 287500 61900 287800
rect 62200 287500 62400 287800
rect 62700 287500 62900 287800
rect 63200 287500 63400 287800
rect 63700 287500 63900 287800
rect 64200 287500 64400 287800
rect 64700 287500 64900 287800
rect 65200 287500 65400 287800
rect 65700 287500 65900 287800
rect 66200 287500 66400 287800
rect 66700 287500 66900 287800
rect 67200 287500 67400 287800
rect 67700 287500 67900 287800
rect 68200 287500 68400 287800
rect 68700 287500 68900 287800
rect 69200 287500 69400 287800
rect 69700 287500 69900 287800
rect 70200 287500 70400 287800
rect 70700 287500 70900 287800
rect 71200 287500 71400 287800
rect 71700 287500 71900 287800
rect 72200 287500 72400 287800
rect 72700 287500 72900 287800
rect 73200 287500 73400 287800
rect 73700 287500 74200 287800
rect 9600 287400 74200 287500
rect 9600 287200 16100 287400
rect 16300 287200 25800 287400
rect 26000 287300 74200 287400
rect 26000 287200 59400 287300
rect 9600 287000 59400 287200
rect 59700 287000 59900 287300
rect 60200 287000 60400 287300
rect 60700 287000 60900 287300
rect 61200 287000 61400 287300
rect 61700 287000 61900 287300
rect 62200 287000 62400 287300
rect 62700 287000 62900 287300
rect 63200 287000 63400 287300
rect 63700 287000 63900 287300
rect 64200 287000 64400 287300
rect 64700 287000 64900 287300
rect 65200 287000 65400 287300
rect 65700 287000 65900 287300
rect 66200 287000 66400 287300
rect 66700 287000 66900 287300
rect 67200 287000 67400 287300
rect 67700 287000 67900 287300
rect 68200 287000 68400 287300
rect 68700 287000 68900 287300
rect 69200 287000 69400 287300
rect 69700 287000 69900 287300
rect 70200 287000 70400 287300
rect 70700 287000 70900 287300
rect 71200 287000 71400 287300
rect 71700 287000 71900 287300
rect 72200 287000 72400 287300
rect 72700 287000 72900 287300
rect 73200 287000 73400 287300
rect 73700 287000 74200 287300
rect 9600 286800 16100 287000
rect 16300 286800 25800 287000
rect 26000 286800 74200 287000
rect 9600 286600 59400 286800
rect 9600 286400 16100 286600
rect 16300 286400 25800 286600
rect 26000 286500 59400 286600
rect 59700 286500 59900 286800
rect 60200 286500 60400 286800
rect 60700 286500 60900 286800
rect 61200 286500 61400 286800
rect 61700 286500 61900 286800
rect 62200 286500 62400 286800
rect 62700 286500 62900 286800
rect 63200 286500 63400 286800
rect 63700 286500 63900 286800
rect 64200 286500 64400 286800
rect 64700 286500 64900 286800
rect 65200 286500 65400 286800
rect 65700 286500 65900 286800
rect 66200 286500 66400 286800
rect 66700 286500 66900 286800
rect 67200 286500 67400 286800
rect 67700 286500 67900 286800
rect 68200 286500 68400 286800
rect 68700 286500 68900 286800
rect 69200 286500 69400 286800
rect 69700 286500 69900 286800
rect 70200 286500 70400 286800
rect 70700 286500 70900 286800
rect 71200 286500 71400 286800
rect 71700 286500 71900 286800
rect 72200 286500 72400 286800
rect 72700 286500 72900 286800
rect 73200 286500 73400 286800
rect 73700 286500 74200 286800
rect 26000 286400 74200 286500
rect 9600 286300 74200 286400
rect 9600 286200 59400 286300
rect 9600 286000 16100 286200
rect 16300 286000 25800 286200
rect 26000 286000 59400 286200
rect 59700 286000 59900 286300
rect 60200 286000 60400 286300
rect 60700 286000 60900 286300
rect 61200 286000 61400 286300
rect 61700 286000 61900 286300
rect 62200 286000 62400 286300
rect 62700 286000 62900 286300
rect 63200 286000 63400 286300
rect 63700 286000 63900 286300
rect 64200 286000 64400 286300
rect 64700 286000 64900 286300
rect 65200 286000 65400 286300
rect 65700 286000 65900 286300
rect 66200 286000 66400 286300
rect 66700 286000 66900 286300
rect 67200 286000 67400 286300
rect 67700 286000 67900 286300
rect 68200 286000 68400 286300
rect 68700 286000 68900 286300
rect 69200 286000 69400 286300
rect 69700 286000 69900 286300
rect 70200 286000 70400 286300
rect 70700 286000 70900 286300
rect 71200 286000 71400 286300
rect 71700 286000 71900 286300
rect 72200 286000 72400 286300
rect 72700 286000 72900 286300
rect 73200 286000 73400 286300
rect 73700 286000 74200 286300
rect 9600 285800 74200 286000
rect 6740 280500 13280 280520
rect 6740 280430 13190 280500
rect 13260 280430 13280 280500
rect 6740 280390 13280 280430
rect 6740 280320 13080 280390
rect 13150 280320 13280 280390
rect 6740 280300 13280 280320
rect 6740 280022 6980 280300
rect 6740 276678 6891 280022
rect 6955 276678 6980 280022
rect 7109 279910 10231 279911
rect 7109 276790 7110 279910
rect 10230 276790 10231 279910
rect 14510 278550 35300 278580
rect 14510 278370 14540 278550
rect 14640 278540 21980 278550
rect 14640 278400 15000 278540
rect 15140 278400 15200 278540
rect 15340 278400 21980 278540
rect 14640 278370 21980 278400
rect 14510 278320 21980 278370
rect 14510 278180 15000 278320
rect 15140 278180 15200 278320
rect 15340 278310 21980 278320
rect 22220 278310 22320 278550
rect 22560 278400 35300 278550
rect 22560 278310 34000 278400
rect 15340 278190 34000 278310
rect 15340 278180 21980 278190
rect 14510 278130 21980 278180
rect 14510 277950 14540 278130
rect 14640 278100 21980 278130
rect 14640 277960 15000 278100
rect 15140 277960 15200 278100
rect 15340 277960 21980 278100
rect 14640 277950 21980 277960
rect 22220 277950 22320 278190
rect 22560 278100 34000 278190
rect 34300 278100 34400 278400
rect 34700 278100 34800 278400
rect 35100 278100 35300 278400
rect 22560 277950 35300 278100
rect 14510 277920 35300 277950
rect 7109 276789 10231 276790
rect 6740 276222 6980 276678
rect 6740 272878 6891 276222
rect 6955 272878 6980 276222
rect 8450 276620 8810 276789
rect 8450 276600 14160 276620
rect 8450 276510 14040 276600
rect 14140 276510 14160 276600
rect 8450 276410 14160 276510
rect 8450 276320 14040 276410
rect 14140 276320 14160 276410
rect 8450 276300 14160 276320
rect 8450 276111 8810 276300
rect 34459 276140 34701 276141
rect 7109 276110 10231 276111
rect 7109 272990 7110 276110
rect 10230 272990 10231 276110
rect 34459 275900 34460 276140
rect 34700 275900 34701 276140
rect 34459 275899 34701 275900
rect 37659 276140 37901 276141
rect 37659 275900 37660 276140
rect 37900 275900 37901 276140
rect 37659 275899 37901 275900
rect 40979 276140 41221 276141
rect 40979 275900 40980 276140
rect 41220 275900 41221 276140
rect 40979 275899 41221 275900
rect 12869 275470 13121 275471
rect 12869 275220 12870 275470
rect 13120 275220 13121 275470
rect 12869 275219 13121 275220
rect 14519 274130 14781 274131
rect 14519 273870 14520 274130
rect 14780 273870 14781 274130
rect 14519 273869 14781 273870
rect 16069 274130 16331 274131
rect 16069 273870 16070 274130
rect 16330 273870 16331 274130
rect 16069 273869 16331 273870
rect 22849 274070 23101 274071
rect 22849 273820 22850 274070
rect 23100 273820 23101 274070
rect 22849 273819 23101 273820
rect 21329 273810 21581 273811
rect 12869 273570 13121 273571
rect 12359 273330 12631 273331
rect 12359 273060 12360 273330
rect 12630 273060 12631 273330
rect 12869 273320 12870 273570
rect 13120 273320 13121 273570
rect 21329 273560 21330 273810
rect 21580 273560 21581 273810
rect 21329 273559 21581 273560
rect 24320 273670 26320 273730
rect 24320 273590 25860 273670
rect 25940 273590 26080 273670
rect 26160 273590 26220 273670
rect 26300 273590 26320 273670
rect 24320 273550 26320 273590
rect 15609 273540 15871 273541
rect 12869 273319 13121 273320
rect 13999 273330 14271 273331
rect 12359 273059 12631 273060
rect 13999 273060 14000 273330
rect 14270 273060 14271 273330
rect 15609 273280 15610 273540
rect 15870 273280 15871 273540
rect 24560 273510 26320 273550
rect 15609 273279 15871 273280
rect 13999 273059 14271 273060
rect 7109 272989 10231 272990
rect 6740 272422 6980 272878
rect 6740 269078 6891 272422
rect 6955 269078 6980 272422
rect 8450 272311 8810 272989
rect 14519 272870 14781 272871
rect 14519 272610 14520 272870
rect 14780 272610 14781 272870
rect 14519 272609 14781 272610
rect 16069 272870 16331 272871
rect 16069 272610 16070 272870
rect 16330 272610 16331 272870
rect 27300 273010 41780 273090
rect 27300 272890 27470 273010
rect 27590 272890 33980 273010
rect 16069 272609 16331 272610
rect 18709 272780 18971 272781
rect 18709 272520 18710 272780
rect 18970 272520 18971 272780
rect 18709 272519 18971 272520
rect 20229 272780 20491 272781
rect 20229 272520 20230 272780
rect 20490 272520 20491 272780
rect 21749 272780 22001 272781
rect 21749 272530 21750 272780
rect 22000 272530 22001 272780
rect 21749 272529 22001 272530
rect 23279 272780 23531 272781
rect 23279 272530 23280 272780
rect 23530 272530 23531 272780
rect 23279 272529 23531 272530
rect 27300 272770 33980 272890
rect 34220 272770 34460 273010
rect 34700 272770 34940 273010
rect 35180 272770 37180 273010
rect 37420 272770 37660 273010
rect 37900 272770 38140 273010
rect 38380 272770 40500 273010
rect 40740 272770 40980 273010
rect 41220 272770 41460 273010
rect 41700 272770 41780 273010
rect 27300 272680 41780 272770
rect 27300 272590 28370 272680
rect 28460 272670 41780 272680
rect 28460 272590 28750 272670
rect 27300 272580 28750 272590
rect 28840 272580 30190 272670
rect 30280 272580 41780 272670
rect 20229 272519 20491 272520
rect 7109 272310 10231 272311
rect 7109 269190 7110 272310
rect 10230 269190 10231 272310
rect 12359 272280 12631 272281
rect 12359 272010 12360 272280
rect 12630 272010 12631 272280
rect 12359 272009 12631 272010
rect 13999 272280 14271 272281
rect 13999 272010 14000 272280
rect 14270 272010 14271 272280
rect 27300 272450 41780 272580
rect 27300 272390 33980 272450
rect 27300 272270 27480 272390
rect 27600 272270 33980 272390
rect 27300 272210 33980 272270
rect 34220 272210 34460 272450
rect 34700 272210 34940 272450
rect 35180 272210 37180 272450
rect 37420 272210 37660 272450
rect 37900 272210 38140 272450
rect 38380 272210 40500 272450
rect 40740 272210 40980 272450
rect 41220 272210 41460 272450
rect 41700 272210 41780 272450
rect 27300 272130 41780 272210
rect 13999 272009 14271 272010
rect 15609 272040 15871 272041
rect 12869 271990 13121 271991
rect 12869 271740 12870 271990
rect 13120 271740 13121 271990
rect 15609 271780 15610 272040
rect 15870 271780 15871 272040
rect 15609 271779 15871 271780
rect 12869 271739 13121 271740
rect 21329 271750 21581 271751
rect 14519 271600 14781 271601
rect 14519 271340 14520 271600
rect 14780 271340 14781 271600
rect 14519 271339 14781 271340
rect 16069 271600 16331 271601
rect 16069 271340 16070 271600
rect 16330 271340 16331 271600
rect 21329 271500 21330 271750
rect 21580 271500 21581 271750
rect 24560 271750 26320 271790
rect 24320 271710 26320 271750
rect 24320 271630 25860 271710
rect 25940 271630 26080 271710
rect 26160 271630 26220 271710
rect 26300 271630 26320 271710
rect 24320 271570 26320 271630
rect 21329 271499 21581 271500
rect 16069 271339 16331 271340
rect 22849 271490 23101 271491
rect 22849 271240 22850 271490
rect 23100 271240 23101 271490
rect 22849 271239 23101 271240
rect 12859 270090 13111 270091
rect 12859 269840 12860 270090
rect 13110 269840 13111 270090
rect 12859 269839 13111 269840
rect 34459 269440 34701 269441
rect 34459 269200 34460 269440
rect 34700 269200 34701 269440
rect 34459 269199 34701 269200
rect 37659 269440 37901 269441
rect 37659 269200 37660 269440
rect 37900 269200 37901 269440
rect 37659 269199 37901 269200
rect 40979 269440 41221 269441
rect 40979 269200 40980 269440
rect 41220 269200 41221 269440
rect 40979 269199 41221 269200
rect 7109 269189 10231 269190
rect 6740 268622 6980 269078
rect 6740 265278 6891 268622
rect 6955 265278 6980 268622
rect 8450 269010 8810 269189
rect 8450 268990 14160 269010
rect 8450 268900 14040 268990
rect 14140 268900 14160 268990
rect 8450 268800 14160 268900
rect 8450 268710 14040 268800
rect 14140 268710 14160 268800
rect 8450 268690 14160 268710
rect 8450 268511 8810 268690
rect 33000 268600 92000 268800
rect 7109 268510 10231 268511
rect 7109 265390 7110 268510
rect 10230 265390 10231 268510
rect 33000 268300 34000 268600
rect 34300 268300 34800 268600
rect 35100 268300 37300 268600
rect 37600 268300 38000 268600
rect 38300 268300 40600 268600
rect 40900 268300 41300 268600
rect 41600 268300 44700 268600
rect 45000 268300 92000 268600
rect 33000 268100 92000 268300
rect 33000 267800 34000 268100
rect 34300 267800 34800 268100
rect 35100 267800 37300 268100
rect 37600 267800 38000 268100
rect 38300 267800 40600 268100
rect 40900 267800 41300 268100
rect 41600 267800 44700 268100
rect 45000 267800 92000 268100
rect 33000 267600 92000 267800
rect 33000 267330 34000 267600
rect 14510 267300 34000 267330
rect 34300 267300 34800 267600
rect 35100 267300 37300 267600
rect 37600 267300 38000 267600
rect 38300 267300 40600 267600
rect 40900 267300 41300 267600
rect 41600 267300 44700 267600
rect 45000 267300 92000 267600
rect 14510 267120 14540 267300
rect 14640 267280 21980 267300
rect 14640 267120 15000 267280
rect 15160 267120 15220 267280
rect 15380 267120 15440 267280
rect 15600 267120 15660 267280
rect 15820 267120 21980 267280
rect 14510 267060 21980 267120
rect 22220 267060 22320 267300
rect 22560 267100 92000 267300
rect 22560 267060 34000 267100
rect 14510 266940 34000 267060
rect 14510 266880 21980 266940
rect 14510 266700 14540 266880
rect 14640 266860 21980 266880
rect 14640 266700 15000 266860
rect 15160 266700 15220 266860
rect 15380 266700 15440 266860
rect 15600 266700 15660 266860
rect 15820 266700 21980 266860
rect 22220 266700 22320 266940
rect 22560 266800 34000 266940
rect 34300 266800 34800 267100
rect 35100 266800 37300 267100
rect 37600 266800 38000 267100
rect 38300 266800 40600 267100
rect 40900 266800 41300 267100
rect 41600 266800 44700 267100
rect 45000 266800 92000 267100
rect 22560 266700 92000 266800
rect 14510 266670 92000 266700
rect 33000 266600 92000 266670
rect 7109 265389 10231 265390
rect 20600 266200 27800 266400
rect 20600 266000 20700 266200
rect 20900 266000 22700 266200
rect 22900 266000 23100 266200
rect 23300 266000 23500 266200
rect 23700 266000 23900 266200
rect 24100 266000 24300 266200
rect 24500 266000 24700 266200
rect 24900 266000 25100 266200
rect 25300 266000 25500 266200
rect 25700 266000 25900 266200
rect 26100 266000 26300 266200
rect 26500 266000 26700 266200
rect 26900 266000 27100 266200
rect 27300 266000 27500 266200
rect 27700 266000 27800 266200
rect 20600 265800 27800 266000
rect 20600 265600 20700 265800
rect 20900 265600 22700 265800
rect 22900 265600 23100 265800
rect 23300 265600 23500 265800
rect 23700 265600 23900 265800
rect 24100 265600 24300 265800
rect 24500 265600 24700 265800
rect 24900 265600 25100 265800
rect 25300 265600 25500 265800
rect 25700 265600 25900 265800
rect 26100 265600 26300 265800
rect 26500 265600 26700 265800
rect 26900 265600 27100 265800
rect 27300 265600 27500 265800
rect 27700 265600 27800 265800
rect 20600 265400 27800 265600
rect 6740 265020 6980 265278
rect 20600 265200 20700 265400
rect 20900 265200 22700 265400
rect 22900 265200 23100 265400
rect 23300 265200 23500 265400
rect 23700 265200 23900 265400
rect 24100 265200 24300 265400
rect 24500 265200 24700 265400
rect 24900 265200 25100 265400
rect 25300 265200 25500 265400
rect 25700 265200 25900 265400
rect 26100 265200 26300 265400
rect 26500 265200 26700 265400
rect 26900 265200 27100 265400
rect 27300 265200 27500 265400
rect 27700 265200 27800 265400
rect 6740 265000 13280 265020
rect 6740 264930 13080 265000
rect 13150 264930 13280 265000
rect 6740 264890 13280 264930
rect 6740 264820 13190 264890
rect 13260 264820 13280 264890
rect 6740 264800 13280 264820
rect 20600 265000 27800 265200
rect 20600 264800 20700 265000
rect 20900 264800 22700 265000
rect 22900 264800 23100 265000
rect 23300 264800 23500 265000
rect 23700 264800 23900 265000
rect 24100 264800 24300 265000
rect 24500 264800 24700 265000
rect 24900 264800 25100 265000
rect 25300 264800 25500 265000
rect 25700 264800 25900 265000
rect 26100 264800 26300 265000
rect 26500 264800 26700 265000
rect 26900 264800 27100 265000
rect 27300 264800 27500 265000
rect 27700 264800 27800 265000
rect 20600 264600 27800 264800
rect 33000 266300 34000 266600
rect 34300 266300 34800 266600
rect 35100 266300 37300 266600
rect 37600 266300 38000 266600
rect 38300 266300 40600 266600
rect 40900 266300 41300 266600
rect 41600 266300 44700 266600
rect 45000 266300 92000 266600
rect 33000 266100 92000 266300
rect 33000 265800 34000 266100
rect 34300 265800 34800 266100
rect 35100 265800 37300 266100
rect 37600 265800 38000 266100
rect 38300 265800 40600 266100
rect 40900 265800 41300 266100
rect 41600 265800 44700 266100
rect 45000 265800 92000 266100
rect 33000 265600 92000 265800
rect 33000 265300 34000 265600
rect 34300 265300 34800 265600
rect 35100 265300 37300 265600
rect 37600 265300 38000 265600
rect 38300 265300 40600 265600
rect 40900 265300 41300 265600
rect 41600 265300 44700 265600
rect 45000 265300 92000 265600
rect 33000 265100 92000 265300
rect 33000 264800 34000 265100
rect 34300 264800 34800 265100
rect 35100 264800 37300 265100
rect 37600 264800 38000 265100
rect 38300 264800 40600 265100
rect 40900 264800 41300 265100
rect 41600 264800 44700 265100
rect 45000 264800 92000 265100
rect 33000 264600 92000 264800
rect 33000 264300 34000 264600
rect 34300 264300 34800 264600
rect 35100 264300 37300 264600
rect 37600 264300 38000 264600
rect 38300 264300 40600 264600
rect 40900 264300 41300 264600
rect 41600 264300 44700 264600
rect 45000 264300 92000 264600
rect 33000 264100 92000 264300
rect 33000 263800 34000 264100
rect 34300 263800 34800 264100
rect 35100 263800 37300 264100
rect 37600 263800 38000 264100
rect 38300 263800 40600 264100
rect 40900 263800 41300 264100
rect 41600 263800 44700 264100
rect 45000 263800 92000 264100
rect 33000 263600 92000 263800
rect 33000 263300 34000 263600
rect 34300 263300 34800 263600
rect 35100 263300 37300 263600
rect 37600 263300 38000 263600
rect 38300 263300 40600 263600
rect 40900 263300 41300 263600
rect 41600 263300 44700 263600
rect 45000 263300 92000 263600
rect 33000 263100 92000 263300
rect 33000 262800 34000 263100
rect 34300 262800 34800 263100
rect 35100 262800 37300 263100
rect 37600 262800 38000 263100
rect 38300 262800 40600 263100
rect 40900 262800 41300 263100
rect 41600 262800 44700 263100
rect 45000 262800 92000 263100
rect 33000 262600 92000 262800
rect 33000 262300 34000 262600
rect 34300 262300 34800 262600
rect 35100 262300 37300 262600
rect 37600 262300 38000 262600
rect 38300 262300 40600 262600
rect 40900 262300 41300 262600
rect 41600 262300 44700 262600
rect 45000 262300 92000 262600
rect 33000 262100 92000 262300
rect 33000 261800 34000 262100
rect 34300 261800 34800 262100
rect 35100 261800 37300 262100
rect 37600 261800 38000 262100
rect 38300 261800 40600 262100
rect 40900 261800 41300 262100
rect 41600 261800 44700 262100
rect 45000 261800 92000 262100
rect 33000 261600 92000 261800
rect 33000 261300 34000 261600
rect 34300 261300 34800 261600
rect 35100 261300 37300 261600
rect 37600 261300 38000 261600
rect 38300 261300 40600 261600
rect 40900 261300 41300 261600
rect 41600 261300 44700 261600
rect 45000 261300 92000 261600
rect 33000 261100 92000 261300
rect 33000 260800 34000 261100
rect 34300 260800 34800 261100
rect 35100 260800 37300 261100
rect 37600 260800 38000 261100
rect 38300 260800 40600 261100
rect 40900 260800 41300 261100
rect 41600 260800 44700 261100
rect 45000 260800 92000 261100
rect 33000 260600 92000 260800
rect 9600 252400 74200 252600
rect 5700 252320 6060 252340
rect 5700 252200 5820 252320
rect 5940 252200 6060 252320
rect 5700 252120 6060 252200
rect 5700 252000 5820 252120
rect 5940 252000 6060 252120
rect 5700 251920 6060 252000
rect 5700 251800 5820 251920
rect 5940 251800 6060 251920
rect 5700 251720 6060 251800
rect 5700 251600 5820 251720
rect 5940 251600 6060 251720
rect 5700 251520 6060 251600
rect 5700 251400 5820 251520
rect 5940 251400 6060 251520
rect 5700 249200 6060 251400
rect 9600 252200 9800 252400
rect 10000 252200 10200 252400
rect 10400 252200 10600 252400
rect 10800 252200 11000 252400
rect 11200 252200 11400 252400
rect 11600 252200 59500 252400
rect 9600 252100 59500 252200
rect 59800 252100 60100 252400
rect 60400 252100 60700 252400
rect 61000 252100 61400 252400
rect 61700 252100 62000 252400
rect 62300 252100 62600 252400
rect 62900 252100 63200 252400
rect 63500 252100 63800 252400
rect 64100 252100 64400 252400
rect 64700 252100 65100 252400
rect 65400 252100 65700 252400
rect 66000 252100 66300 252400
rect 66600 252100 66900 252400
rect 67200 252100 67500 252400
rect 67800 252100 68100 252400
rect 68400 252100 68700 252400
rect 69000 252100 69300 252400
rect 69600 252100 69900 252400
rect 70200 252100 70600 252400
rect 70900 252100 71300 252400
rect 71600 252100 72000 252400
rect 72300 252100 72800 252400
rect 73100 252100 73500 252400
rect 73800 252100 74200 252400
rect 9600 252000 74200 252100
rect 9600 251800 9800 252000
rect 10000 251800 10200 252000
rect 10400 251800 10600 252000
rect 10800 251800 11000 252000
rect 11200 251800 11400 252000
rect 11600 251800 74200 252000
rect 9600 251700 74200 251800
rect 9600 251600 59500 251700
rect 9600 251400 9800 251600
rect 10000 251400 10200 251600
rect 10400 251400 10600 251600
rect 10800 251400 11000 251600
rect 11200 251400 11400 251600
rect 11600 251400 59500 251600
rect 59800 251400 60100 251700
rect 60400 251400 60700 251700
rect 61000 251400 61400 251700
rect 61700 251400 62000 251700
rect 62300 251400 62600 251700
rect 62900 251400 63200 251700
rect 63500 251400 63800 251700
rect 64100 251400 64400 251700
rect 64700 251400 65100 251700
rect 65400 251400 65700 251700
rect 66000 251400 66300 251700
rect 66600 251400 66900 251700
rect 67200 251400 67500 251700
rect 67800 251400 68100 251700
rect 68400 251400 68700 251700
rect 69000 251400 69300 251700
rect 69600 251400 69900 251700
rect 70200 251400 70600 251700
rect 70900 251400 71300 251700
rect 71600 251400 72000 251700
rect 72300 251400 72800 251700
rect 73100 251400 73500 251700
rect 73800 251400 74200 251700
rect 9600 251200 74200 251400
rect 5700 249000 20000 249200
rect 5700 248800 5800 249000
rect 6000 248800 6200 249000
rect 6400 248800 6600 249000
rect 6800 248800 7000 249000
rect 7200 248800 7400 249000
rect 7600 248800 7800 249000
rect 8000 248800 19300 249000
rect 19500 248800 19700 249000
rect 19900 248800 20000 249000
rect 5700 248600 20000 248800
rect 5700 248400 5800 248600
rect 6000 248400 6200 248600
rect 6400 248400 6600 248600
rect 6800 248400 7000 248600
rect 7200 248400 7400 248600
rect 7600 248400 7800 248600
rect 8000 248400 19300 248600
rect 19500 248400 19700 248600
rect 19900 248400 20000 248600
rect 5700 248200 20000 248400
rect 5700 248000 5800 248200
rect 6000 248000 6200 248200
rect 6400 248000 6600 248200
rect 6800 248000 7000 248200
rect 7200 248000 7400 248200
rect 7600 248000 7800 248200
rect 8000 248000 19300 248200
rect 19500 248000 19700 248200
rect 19900 248000 20000 248200
rect 5700 247800 20000 248000
rect 5700 247600 5800 247800
rect 6000 247600 6200 247800
rect 6400 247600 6600 247800
rect 6800 247600 7000 247800
rect 7200 247600 7400 247800
rect 7600 247600 7800 247800
rect 8000 247600 19300 247800
rect 19500 247600 19700 247800
rect 19900 247600 20000 247800
rect 5700 247400 20000 247600
rect 5700 247200 5800 247400
rect 6000 247200 6200 247400
rect 6400 247200 6600 247400
rect 6800 247200 7000 247400
rect 7200 247200 7400 247400
rect 7600 247200 7800 247400
rect 8000 247200 19300 247400
rect 19500 247200 19700 247400
rect 19900 247200 20000 247400
rect 5700 247000 20000 247200
rect 5700 246800 5800 247000
rect 6000 246800 6200 247000
rect 6400 246800 6600 247000
rect 6800 246800 7000 247000
rect 7200 246800 7400 247000
rect 7600 246800 7800 247000
rect 8000 246800 19300 247000
rect 19500 246800 19700 247000
rect 19900 246800 20000 247000
rect 5700 246600 20000 246800
rect 5700 246400 5800 246600
rect 6000 246400 6200 246600
rect 6400 246400 6600 246600
rect 6800 246400 7000 246600
rect 7200 246400 7400 246600
rect 7600 246400 7800 246600
rect 8000 246400 19300 246600
rect 19500 246400 19700 246600
rect 19900 246400 20000 246600
rect 5700 246200 20000 246400
rect 5700 246000 5800 246200
rect 6000 246000 6200 246200
rect 6400 246000 6600 246200
rect 6800 246000 7000 246200
rect 7200 246000 7400 246200
rect 7600 246000 7800 246200
rect 8000 246000 19300 246200
rect 19500 246000 19700 246200
rect 19900 246000 20000 246200
rect 5700 245800 20000 246000
rect 5700 245600 5800 245800
rect 6000 245600 6200 245800
rect 6400 245600 6600 245800
rect 6800 245600 7000 245800
rect 7200 245600 7400 245800
rect 7600 245600 7800 245800
rect 8000 245600 19300 245800
rect 19500 245600 19700 245800
rect 19900 245600 20000 245800
rect 5700 245400 20000 245600
rect 5700 245200 5800 245400
rect 6000 245200 6200 245400
rect 6400 245200 6600 245400
rect 6800 245200 7000 245400
rect 7200 245200 7400 245400
rect 7600 245200 7800 245400
rect 8000 245200 19300 245400
rect 19500 245200 19700 245400
rect 19900 245200 20000 245400
rect 5700 245000 20000 245200
rect 5700 244800 5800 245000
rect 6000 244800 6200 245000
rect 6400 244800 6600 245000
rect 6800 244800 7000 245000
rect 7200 244800 7400 245000
rect 7600 244800 7800 245000
rect 8000 244800 19300 245000
rect 19500 244800 19700 245000
rect 19900 244800 20000 245000
rect 5700 244600 20000 244800
rect 5700 244400 5800 244600
rect 6000 244400 6200 244600
rect 6400 244400 6600 244600
rect 6800 244400 7000 244600
rect 7200 244400 7400 244600
rect 7600 244400 7800 244600
rect 8000 244400 19300 244600
rect 19500 244400 19700 244600
rect 19900 244400 20000 244600
rect 5700 244200 20000 244400
rect 9600 241800 11600 244200
rect 9600 241600 9800 241800
rect 10000 241600 10200 241800
rect 10400 241600 10800 241800
rect 11000 241600 11200 241800
rect 11400 241600 11600 241800
rect 9600 241200 11600 241600
rect 9600 241000 9800 241200
rect 10000 241000 10200 241200
rect 10400 241000 10800 241200
rect 11000 241000 11200 241200
rect 11400 241000 11600 241200
rect 9600 240800 11600 241000
rect 16020 242000 35300 242120
rect 16020 241800 16100 242000
rect 16300 241800 33900 242000
rect 16020 241700 33900 241800
rect 34200 241700 34400 242000
rect 34700 241700 34900 242000
rect 35200 241700 35300 242000
rect 16020 241500 16100 241700
rect 16300 241500 35300 241700
rect 16020 241400 35300 241500
rect 16020 241200 16100 241400
rect 16300 241200 35300 241400
rect 16020 241100 33900 241200
rect 16020 240900 16100 241100
rect 16300 240900 33900 241100
rect 34200 240900 34400 241200
rect 34700 240900 34900 241200
rect 35200 240900 35300 241200
rect 16020 240800 35300 240900
rect 59999 218800 60401 218801
rect 59999 218400 60000 218800
rect 60400 218400 60401 218800
rect 59999 218399 60401 218400
rect 60799 218800 61201 218801
rect 60799 218400 60800 218800
rect 61200 218400 61201 218800
rect 60799 218399 61201 218400
rect 61599 218800 62001 218801
rect 61599 218400 61600 218800
rect 62000 218400 62001 218800
rect 61599 218399 62001 218400
rect 62399 218800 62801 218801
rect 62399 218400 62400 218800
rect 62800 218400 62801 218800
rect 62399 218399 62801 218400
rect 63199 218800 63601 218801
rect 63199 218400 63200 218800
rect 63600 218400 63601 218800
rect 63199 218399 63601 218400
rect 63999 218800 64401 218801
rect 63999 218400 64000 218800
rect 64400 218400 64401 218800
rect 63999 218399 64401 218400
rect 68999 218800 69401 218801
rect 68999 218400 69000 218800
rect 69400 218400 69401 218800
rect 68999 218399 69401 218400
rect 69799 218800 70201 218801
rect 69799 218400 69800 218800
rect 70200 218400 70201 218800
rect 69799 218399 70201 218400
rect 70599 218800 71001 218801
rect 70599 218400 70600 218800
rect 71000 218400 71001 218800
rect 70599 218399 71001 218400
rect 71399 218800 71801 218801
rect 71399 218400 71400 218800
rect 71800 218400 71801 218800
rect 71399 218399 71801 218400
rect 72199 218800 72601 218801
rect 72199 218400 72200 218800
rect 72600 218400 72601 218800
rect 72199 218399 72601 218400
rect 72999 218800 73401 218801
rect 72999 218400 73000 218800
rect 73400 218400 73401 218800
rect 72999 218399 73401 218400
rect 59999 218000 60401 218001
rect 59999 217600 60000 218000
rect 60400 217600 60401 218000
rect 59999 217599 60401 217600
rect 60799 218000 61201 218001
rect 60799 217600 60800 218000
rect 61200 217600 61201 218000
rect 60799 217599 61201 217600
rect 61599 218000 62001 218001
rect 61599 217600 61600 218000
rect 62000 217600 62001 218000
rect 61599 217599 62001 217600
rect 62399 218000 62801 218001
rect 62399 217600 62400 218000
rect 62800 217600 62801 218000
rect 62399 217599 62801 217600
rect 63199 218000 63601 218001
rect 63199 217600 63200 218000
rect 63600 217600 63601 218000
rect 63199 217599 63601 217600
rect 63999 218000 64401 218001
rect 63999 217600 64000 218000
rect 64400 217600 64401 218000
rect 63999 217599 64401 217600
rect 68999 218000 69401 218001
rect 68999 217600 69000 218000
rect 69400 217600 69401 218000
rect 68999 217599 69401 217600
rect 69799 218000 70201 218001
rect 69799 217600 69800 218000
rect 70200 217600 70201 218000
rect 69799 217599 70201 217600
rect 70599 218000 71001 218001
rect 70599 217600 70600 218000
rect 71000 217600 71001 218000
rect 70599 217599 71001 217600
rect 71399 218000 71801 218001
rect 71399 217600 71400 218000
rect 71800 217600 71801 218000
rect 71399 217599 71801 217600
rect 72199 218000 72601 218001
rect 72199 217600 72200 218000
rect 72600 217600 72601 218000
rect 72199 217599 72601 217600
rect 72999 218000 73401 218001
rect 72999 217600 73000 218000
rect 73400 217600 73401 218000
rect 72999 217599 73401 217600
rect 59999 217200 60401 217201
rect 59999 216800 60000 217200
rect 60400 216800 60401 217200
rect 59999 216799 60401 216800
rect 60799 217200 61201 217201
rect 60799 216800 60800 217200
rect 61200 216800 61201 217200
rect 60799 216799 61201 216800
rect 61599 217200 62001 217201
rect 61599 216800 61600 217200
rect 62000 216800 62001 217200
rect 61599 216799 62001 216800
rect 62399 217200 62801 217201
rect 62399 216800 62400 217200
rect 62800 216800 62801 217200
rect 62399 216799 62801 216800
rect 63199 217200 63601 217201
rect 63199 216800 63200 217200
rect 63600 216800 63601 217200
rect 63199 216799 63601 216800
rect 63999 217200 64401 217201
rect 63999 216800 64000 217200
rect 64400 216800 64401 217200
rect 63999 216799 64401 216800
rect 68999 217200 69401 217201
rect 68999 216800 69000 217200
rect 69400 216800 69401 217200
rect 68999 216799 69401 216800
rect 69799 217200 70201 217201
rect 69799 216800 69800 217200
rect 70200 216800 70201 217200
rect 69799 216799 70201 216800
rect 70599 217200 71001 217201
rect 70599 216800 70600 217200
rect 71000 216800 71001 217200
rect 70599 216799 71001 216800
rect 71399 217200 71801 217201
rect 71399 216800 71400 217200
rect 71800 216800 71801 217200
rect 71399 216799 71801 216800
rect 72199 217200 72601 217201
rect 72199 216800 72200 217200
rect 72600 216800 72601 217200
rect 72199 216799 72601 216800
rect 72999 217200 73401 217201
rect 72999 216800 73000 217200
rect 73400 216800 73401 217200
rect 72999 216799 73401 216800
rect 59999 216400 60401 216401
rect 59999 216000 60000 216400
rect 60400 216000 60401 216400
rect 59999 215999 60401 216000
rect 60799 216400 61201 216401
rect 60799 216000 60800 216400
rect 61200 216000 61201 216400
rect 60799 215999 61201 216000
rect 61599 216400 62001 216401
rect 61599 216000 61600 216400
rect 62000 216000 62001 216400
rect 61599 215999 62001 216000
rect 62399 216400 62801 216401
rect 62399 216000 62400 216400
rect 62800 216000 62801 216400
rect 62399 215999 62801 216000
rect 63199 216400 63601 216401
rect 63199 216000 63200 216400
rect 63600 216000 63601 216400
rect 63199 215999 63601 216000
rect 63999 216400 64401 216401
rect 63999 216000 64000 216400
rect 64400 216000 64401 216400
rect 63999 215999 64401 216000
rect 68999 216400 69401 216401
rect 68999 216000 69000 216400
rect 69400 216000 69401 216400
rect 68999 215999 69401 216000
rect 69799 216400 70201 216401
rect 69799 216000 69800 216400
rect 70200 216000 70201 216400
rect 69799 215999 70201 216000
rect 70599 216400 71001 216401
rect 70599 216000 70600 216400
rect 71000 216000 71001 216400
rect 70599 215999 71001 216000
rect 71399 216400 71801 216401
rect 71399 216000 71400 216400
rect 71800 216000 71801 216400
rect 71399 215999 71801 216000
rect 72199 216400 72601 216401
rect 72199 216000 72200 216400
rect 72600 216000 72601 216400
rect 72199 215999 72601 216000
rect 72999 216400 73401 216401
rect 72999 216000 73000 216400
rect 73400 216000 73401 216400
rect 72999 215999 73401 216000
rect 59999 215600 60401 215601
rect 59999 215200 60000 215600
rect 60400 215200 60401 215600
rect 59999 215199 60401 215200
rect 60799 215600 61201 215601
rect 60799 215200 60800 215600
rect 61200 215200 61201 215600
rect 60799 215199 61201 215200
rect 61599 215600 62001 215601
rect 61599 215200 61600 215600
rect 62000 215200 62001 215600
rect 61599 215199 62001 215200
rect 62399 215600 62801 215601
rect 62399 215200 62400 215600
rect 62800 215200 62801 215600
rect 62399 215199 62801 215200
rect 63199 215600 63601 215601
rect 63199 215200 63200 215600
rect 63600 215200 63601 215600
rect 63199 215199 63601 215200
rect 63999 215600 64401 215601
rect 63999 215200 64000 215600
rect 64400 215200 64401 215600
rect 63999 215199 64401 215200
rect 68999 215600 69401 215601
rect 68999 215200 69000 215600
rect 69400 215200 69401 215600
rect 68999 215199 69401 215200
rect 69799 215600 70201 215601
rect 69799 215200 69800 215600
rect 70200 215200 70201 215600
rect 69799 215199 70201 215200
rect 70599 215600 71001 215601
rect 70599 215200 70600 215600
rect 71000 215200 71001 215600
rect 70599 215199 71001 215200
rect 71399 215600 71801 215601
rect 71399 215200 71400 215600
rect 71800 215200 71801 215600
rect 71399 215199 71801 215200
rect 72199 215600 72601 215601
rect 72199 215200 72200 215600
rect 72600 215200 72601 215600
rect 72199 215199 72601 215200
rect 72999 215600 73401 215601
rect 72999 215200 73000 215600
rect 73400 215200 73401 215600
rect 72999 215199 73401 215200
rect 59999 214800 60401 214801
rect 59999 214400 60000 214800
rect 60400 214400 60401 214800
rect 59999 214399 60401 214400
rect 60799 214800 61201 214801
rect 60799 214400 60800 214800
rect 61200 214400 61201 214800
rect 60799 214399 61201 214400
rect 61599 214800 62001 214801
rect 61599 214400 61600 214800
rect 62000 214400 62001 214800
rect 61599 214399 62001 214400
rect 62399 214800 62801 214801
rect 62399 214400 62400 214800
rect 62800 214400 62801 214800
rect 62399 214399 62801 214400
rect 63199 214800 63601 214801
rect 63199 214400 63200 214800
rect 63600 214400 63601 214800
rect 63199 214399 63601 214400
rect 63999 214800 64401 214801
rect 63999 214400 64000 214800
rect 64400 214400 64401 214800
rect 63999 214399 64401 214400
rect 68999 214800 69401 214801
rect 68999 214400 69000 214800
rect 69400 214400 69401 214800
rect 68999 214399 69401 214400
rect 69799 214800 70201 214801
rect 69799 214400 69800 214800
rect 70200 214400 70201 214800
rect 69799 214399 70201 214400
rect 70599 214800 71001 214801
rect 70599 214400 70600 214800
rect 71000 214400 71001 214800
rect 70599 214399 71001 214400
rect 71399 214800 71801 214801
rect 71399 214400 71400 214800
rect 71800 214400 71801 214800
rect 71399 214399 71801 214400
rect 72199 214800 72601 214801
rect 72199 214400 72200 214800
rect 72600 214400 72601 214800
rect 72199 214399 72601 214400
rect 72999 214800 73401 214801
rect 72999 214400 73000 214800
rect 73400 214400 73401 214800
rect 72999 214399 73401 214400
rect 68999 210200 69401 210201
rect 59999 210000 60401 210001
rect 59999 209600 60000 210000
rect 60400 209600 60401 210000
rect 59999 209599 60401 209600
rect 60799 210000 61201 210001
rect 60799 209600 60800 210000
rect 61200 209600 61201 210000
rect 60799 209599 61201 209600
rect 61599 210000 62001 210001
rect 61599 209600 61600 210000
rect 62000 209600 62001 210000
rect 61599 209599 62001 209600
rect 62399 210000 62801 210001
rect 62399 209600 62400 210000
rect 62800 209600 62801 210000
rect 62399 209599 62801 209600
rect 63199 210000 63601 210001
rect 63199 209600 63200 210000
rect 63600 209600 63601 210000
rect 63199 209599 63601 209600
rect 63999 210000 64401 210001
rect 63999 209600 64000 210000
rect 64400 209600 64401 210000
rect 68999 209800 69000 210200
rect 69400 209800 69401 210200
rect 68999 209799 69401 209800
rect 69799 210200 70201 210201
rect 69799 209800 69800 210200
rect 70200 209800 70201 210200
rect 69799 209799 70201 209800
rect 70599 210200 71001 210201
rect 70599 209800 70600 210200
rect 71000 209800 71001 210200
rect 70599 209799 71001 209800
rect 71399 210200 71801 210201
rect 71399 209800 71400 210200
rect 71800 209800 71801 210200
rect 71399 209799 71801 209800
rect 72199 210200 72601 210201
rect 72199 209800 72200 210200
rect 72600 209800 72601 210200
rect 72199 209799 72601 209800
rect 72999 210200 73401 210201
rect 72999 209800 73000 210200
rect 73400 209800 73401 210200
rect 72999 209799 73401 209800
rect 63999 209599 64401 209600
rect 68999 209400 69401 209401
rect 59999 209200 60401 209201
rect 59999 208800 60000 209200
rect 60400 208800 60401 209200
rect 59999 208799 60401 208800
rect 60799 209200 61201 209201
rect 60799 208800 60800 209200
rect 61200 208800 61201 209200
rect 60799 208799 61201 208800
rect 61599 209200 62001 209201
rect 61599 208800 61600 209200
rect 62000 208800 62001 209200
rect 61599 208799 62001 208800
rect 62399 209200 62801 209201
rect 62399 208800 62400 209200
rect 62800 208800 62801 209200
rect 62399 208799 62801 208800
rect 63199 209200 63601 209201
rect 63199 208800 63200 209200
rect 63600 208800 63601 209200
rect 63199 208799 63601 208800
rect 63999 209200 64401 209201
rect 63999 208800 64000 209200
rect 64400 208800 64401 209200
rect 68999 209000 69000 209400
rect 69400 209000 69401 209400
rect 68999 208999 69401 209000
rect 69799 209400 70201 209401
rect 69799 209000 69800 209400
rect 70200 209000 70201 209400
rect 69799 208999 70201 209000
rect 70599 209400 71001 209401
rect 70599 209000 70600 209400
rect 71000 209000 71001 209400
rect 70599 208999 71001 209000
rect 71399 209400 71801 209401
rect 71399 209000 71400 209400
rect 71800 209000 71801 209400
rect 71399 208999 71801 209000
rect 72199 209400 72601 209401
rect 72199 209000 72200 209400
rect 72600 209000 72601 209400
rect 72199 208999 72601 209000
rect 72999 209400 73401 209401
rect 72999 209000 73000 209400
rect 73400 209000 73401 209400
rect 72999 208999 73401 209000
rect 63999 208799 64401 208800
rect 68999 208600 69401 208601
rect 59999 208400 60401 208401
rect 59999 208000 60000 208400
rect 60400 208000 60401 208400
rect 59999 207999 60401 208000
rect 60799 208400 61201 208401
rect 60799 208000 60800 208400
rect 61200 208000 61201 208400
rect 60799 207999 61201 208000
rect 61599 208400 62001 208401
rect 61599 208000 61600 208400
rect 62000 208000 62001 208400
rect 61599 207999 62001 208000
rect 62399 208400 62801 208401
rect 62399 208000 62400 208400
rect 62800 208000 62801 208400
rect 62399 207999 62801 208000
rect 63199 208400 63601 208401
rect 63199 208000 63200 208400
rect 63600 208000 63601 208400
rect 63199 207999 63601 208000
rect 63999 208400 64401 208401
rect 63999 208000 64000 208400
rect 64400 208000 64401 208400
rect 68999 208200 69000 208600
rect 69400 208200 69401 208600
rect 68999 208199 69401 208200
rect 69799 208600 70201 208601
rect 69799 208200 69800 208600
rect 70200 208200 70201 208600
rect 69799 208199 70201 208200
rect 70599 208600 71001 208601
rect 70599 208200 70600 208600
rect 71000 208200 71001 208600
rect 70599 208199 71001 208200
rect 71399 208600 71801 208601
rect 71399 208200 71400 208600
rect 71800 208200 71801 208600
rect 71399 208199 71801 208200
rect 72199 208600 72601 208601
rect 72199 208200 72200 208600
rect 72600 208200 72601 208600
rect 72199 208199 72601 208200
rect 72999 208600 73401 208601
rect 72999 208200 73000 208600
rect 73400 208200 73401 208600
rect 72999 208199 73401 208200
rect 63999 207999 64401 208000
rect 68999 207800 69401 207801
rect 59999 207600 60401 207601
rect 59999 207200 60000 207600
rect 60400 207200 60401 207600
rect 59999 207199 60401 207200
rect 60799 207600 61201 207601
rect 60799 207200 60800 207600
rect 61200 207200 61201 207600
rect 60799 207199 61201 207200
rect 61599 207600 62001 207601
rect 61599 207200 61600 207600
rect 62000 207200 62001 207600
rect 61599 207199 62001 207200
rect 62399 207600 62801 207601
rect 62399 207200 62400 207600
rect 62800 207200 62801 207600
rect 62399 207199 62801 207200
rect 63199 207600 63601 207601
rect 63199 207200 63200 207600
rect 63600 207200 63601 207600
rect 63199 207199 63601 207200
rect 63999 207600 64401 207601
rect 63999 207200 64000 207600
rect 64400 207200 64401 207600
rect 68999 207400 69000 207800
rect 69400 207400 69401 207800
rect 68999 207399 69401 207400
rect 69799 207800 70201 207801
rect 69799 207400 69800 207800
rect 70200 207400 70201 207800
rect 69799 207399 70201 207400
rect 70599 207800 71001 207801
rect 70599 207400 70600 207800
rect 71000 207400 71001 207800
rect 70599 207399 71001 207400
rect 71399 207800 71801 207801
rect 71399 207400 71400 207800
rect 71800 207400 71801 207800
rect 71399 207399 71801 207400
rect 72199 207800 72601 207801
rect 72199 207400 72200 207800
rect 72600 207400 72601 207800
rect 72199 207399 72601 207400
rect 72999 207800 73401 207801
rect 72999 207400 73000 207800
rect 73400 207400 73401 207800
rect 72999 207399 73401 207400
rect 63999 207199 64401 207200
rect 68999 207000 69401 207001
rect 59999 206800 60401 206801
rect 59999 206400 60000 206800
rect 60400 206400 60401 206800
rect 59999 206399 60401 206400
rect 60799 206800 61201 206801
rect 60799 206400 60800 206800
rect 61200 206400 61201 206800
rect 60799 206399 61201 206400
rect 61599 206800 62001 206801
rect 61599 206400 61600 206800
rect 62000 206400 62001 206800
rect 61599 206399 62001 206400
rect 62399 206800 62801 206801
rect 62399 206400 62400 206800
rect 62800 206400 62801 206800
rect 62399 206399 62801 206400
rect 63199 206800 63601 206801
rect 63199 206400 63200 206800
rect 63600 206400 63601 206800
rect 63199 206399 63601 206400
rect 63999 206800 64401 206801
rect 63999 206400 64000 206800
rect 64400 206400 64401 206800
rect 68999 206600 69000 207000
rect 69400 206600 69401 207000
rect 68999 206599 69401 206600
rect 69799 207000 70201 207001
rect 69799 206600 69800 207000
rect 70200 206600 70201 207000
rect 69799 206599 70201 206600
rect 70599 207000 71001 207001
rect 70599 206600 70600 207000
rect 71000 206600 71001 207000
rect 70599 206599 71001 206600
rect 71399 207000 71801 207001
rect 71399 206600 71400 207000
rect 71800 206600 71801 207000
rect 71399 206599 71801 206600
rect 72199 207000 72601 207001
rect 72199 206600 72200 207000
rect 72600 206600 72601 207000
rect 72199 206599 72601 206600
rect 72999 207000 73401 207001
rect 72999 206600 73000 207000
rect 73400 206600 73401 207000
rect 72999 206599 73401 206600
rect 63999 206399 64401 206400
rect 68999 206200 69401 206201
rect 59999 206000 60401 206001
rect 59999 205600 60000 206000
rect 60400 205600 60401 206000
rect 59999 205599 60401 205600
rect 60799 206000 61201 206001
rect 60799 205600 60800 206000
rect 61200 205600 61201 206000
rect 60799 205599 61201 205600
rect 61599 206000 62001 206001
rect 61599 205600 61600 206000
rect 62000 205600 62001 206000
rect 61599 205599 62001 205600
rect 62399 206000 62801 206001
rect 62399 205600 62400 206000
rect 62800 205600 62801 206000
rect 62399 205599 62801 205600
rect 63199 206000 63601 206001
rect 63199 205600 63200 206000
rect 63600 205600 63601 206000
rect 63199 205599 63601 205600
rect 63999 206000 64401 206001
rect 63999 205600 64000 206000
rect 64400 205600 64401 206000
rect 68999 205800 69000 206200
rect 69400 205800 69401 206200
rect 68999 205799 69401 205800
rect 69799 206200 70201 206201
rect 69799 205800 69800 206200
rect 70200 205800 70201 206200
rect 69799 205799 70201 205800
rect 70599 206200 71001 206201
rect 70599 205800 70600 206200
rect 71000 205800 71001 206200
rect 70599 205799 71001 205800
rect 71399 206200 71801 206201
rect 71399 205800 71400 206200
rect 71800 205800 71801 206200
rect 71399 205799 71801 205800
rect 72199 206200 72601 206201
rect 72199 205800 72200 206200
rect 72600 205800 72601 206200
rect 72199 205799 72601 205800
rect 72999 206200 73401 206201
rect 72999 205800 73000 206200
rect 73400 205800 73401 206200
rect 72999 205799 73401 205800
rect 63999 205599 64401 205600
rect 83800 177600 92000 260600
rect 285399 219400 285801 219401
rect 285399 219000 285400 219400
rect 285800 219000 285801 219400
rect 285399 218999 285801 219000
rect 286199 219400 286601 219401
rect 286199 219000 286200 219400
rect 286600 219000 286601 219400
rect 286199 218999 286601 219000
rect 286999 219400 287401 219401
rect 286999 219000 287000 219400
rect 287400 219000 287401 219400
rect 286999 218999 287401 219000
rect 287799 219400 288201 219401
rect 287799 219000 287800 219400
rect 288200 219000 288201 219400
rect 287799 218999 288201 219000
rect 288599 219400 289001 219401
rect 288599 219000 288600 219400
rect 289000 219000 289001 219400
rect 288599 218999 289001 219000
rect 289399 219400 289801 219401
rect 289399 219000 289400 219400
rect 289800 219000 289801 219400
rect 289399 218999 289801 219000
rect 285399 218600 285801 218601
rect 285399 218200 285400 218600
rect 285800 218200 285801 218600
rect 285399 218199 285801 218200
rect 286199 218600 286601 218601
rect 286199 218200 286200 218600
rect 286600 218200 286601 218600
rect 286199 218199 286601 218200
rect 286999 218600 287401 218601
rect 286999 218200 287000 218600
rect 287400 218200 287401 218600
rect 286999 218199 287401 218200
rect 287799 218600 288201 218601
rect 287799 218200 287800 218600
rect 288200 218200 288201 218600
rect 287799 218199 288201 218200
rect 288599 218600 289001 218601
rect 288599 218200 288600 218600
rect 289000 218200 289001 218600
rect 288599 218199 289001 218200
rect 289399 218600 289801 218601
rect 289399 218200 289400 218600
rect 289800 218200 289801 218600
rect 289399 218199 289801 218200
rect 285399 217800 285801 217801
rect 285399 217400 285400 217800
rect 285800 217400 285801 217800
rect 285399 217399 285801 217400
rect 286199 217800 286601 217801
rect 286199 217400 286200 217800
rect 286600 217400 286601 217800
rect 286199 217399 286601 217400
rect 286999 217800 287401 217801
rect 286999 217400 287000 217800
rect 287400 217400 287401 217800
rect 286999 217399 287401 217400
rect 287799 217800 288201 217801
rect 287799 217400 287800 217800
rect 288200 217400 288201 217800
rect 287799 217399 288201 217400
rect 288599 217800 289001 217801
rect 288599 217400 288600 217800
rect 289000 217400 289001 217800
rect 288599 217399 289001 217400
rect 289399 217800 289801 217801
rect 289399 217400 289400 217800
rect 289800 217400 289801 217800
rect 289399 217399 289801 217400
rect 285399 217000 285801 217001
rect 285399 216600 285400 217000
rect 285800 216600 285801 217000
rect 285399 216599 285801 216600
rect 286199 217000 286601 217001
rect 286199 216600 286200 217000
rect 286600 216600 286601 217000
rect 286199 216599 286601 216600
rect 286999 217000 287401 217001
rect 286999 216600 287000 217000
rect 287400 216600 287401 217000
rect 286999 216599 287401 216600
rect 287799 217000 288201 217001
rect 287799 216600 287800 217000
rect 288200 216600 288201 217000
rect 287799 216599 288201 216600
rect 288599 217000 289001 217001
rect 288599 216600 288600 217000
rect 289000 216600 289001 217000
rect 288599 216599 289001 216600
rect 289399 217000 289801 217001
rect 289399 216600 289400 217000
rect 289800 216600 289801 217000
rect 289399 216599 289801 216600
rect 285399 216200 285801 216201
rect 285399 215800 285400 216200
rect 285800 215800 285801 216200
rect 285399 215799 285801 215800
rect 286199 216200 286601 216201
rect 286199 215800 286200 216200
rect 286600 215800 286601 216200
rect 286199 215799 286601 215800
rect 286999 216200 287401 216201
rect 286999 215800 287000 216200
rect 287400 215800 287401 216200
rect 286999 215799 287401 215800
rect 287799 216200 288201 216201
rect 287799 215800 287800 216200
rect 288200 215800 288201 216200
rect 287799 215799 288201 215800
rect 288599 216200 289001 216201
rect 288599 215800 288600 216200
rect 289000 215800 289001 216200
rect 288599 215799 289001 215800
rect 289399 216200 289801 216201
rect 289399 215800 289400 216200
rect 289800 215800 289801 216200
rect 289399 215799 289801 215800
rect 285399 215400 285801 215401
rect 285399 215000 285400 215400
rect 285800 215000 285801 215400
rect 285399 214999 285801 215000
rect 286199 215400 286601 215401
rect 286199 215000 286200 215400
rect 286600 215000 286601 215400
rect 286199 214999 286601 215000
rect 286999 215400 287401 215401
rect 286999 215000 287000 215400
rect 287400 215000 287401 215400
rect 286999 214999 287401 215000
rect 287799 215400 288201 215401
rect 287799 215000 287800 215400
rect 288200 215000 288201 215400
rect 287799 214999 288201 215000
rect 288599 215400 289001 215401
rect 288599 215000 288600 215400
rect 289000 215000 289001 215400
rect 288599 214999 289001 215000
rect 289399 215400 289801 215401
rect 289399 215000 289400 215400
rect 289800 215000 289801 215400
rect 289399 214999 289801 215000
rect 285199 214600 285601 214601
rect 285199 214200 285200 214600
rect 285600 214200 285601 214600
rect 285199 214199 285601 214200
rect 285999 214600 286401 214601
rect 285999 214200 286000 214600
rect 286400 214200 286401 214600
rect 285999 214199 286401 214200
rect 286799 214600 287201 214601
rect 286799 214200 286800 214600
rect 287200 214200 287201 214600
rect 286799 214199 287201 214200
rect 287599 214600 288001 214601
rect 287599 214200 287600 214600
rect 288000 214200 288001 214600
rect 287599 214199 288001 214200
rect 288399 214600 288801 214601
rect 288399 214200 288400 214600
rect 288800 214200 288801 214600
rect 288399 214199 288801 214200
rect 289199 214600 289601 214601
rect 289199 214200 289200 214600
rect 289600 214200 289601 214600
rect 289199 214199 289601 214200
rect 285199 213800 285601 213801
rect 285199 213400 285200 213800
rect 285600 213400 285601 213800
rect 285199 213399 285601 213400
rect 285999 213800 286401 213801
rect 285999 213400 286000 213800
rect 286400 213400 286401 213800
rect 285999 213399 286401 213400
rect 286799 213800 287201 213801
rect 286799 213400 286800 213800
rect 287200 213400 287201 213800
rect 286799 213399 287201 213400
rect 287599 213800 288001 213801
rect 287599 213400 287600 213800
rect 288000 213400 288001 213800
rect 287599 213399 288001 213400
rect 288399 213800 288801 213801
rect 288399 213400 288400 213800
rect 288800 213400 288801 213800
rect 288399 213399 288801 213400
rect 289199 213800 289601 213801
rect 289199 213400 289200 213800
rect 289600 213400 289601 213800
rect 289199 213399 289601 213400
rect 285199 213000 285601 213001
rect 285199 212600 285200 213000
rect 285600 212600 285601 213000
rect 285199 212599 285601 212600
rect 285999 213000 286401 213001
rect 285999 212600 286000 213000
rect 286400 212600 286401 213000
rect 285999 212599 286401 212600
rect 286799 213000 287201 213001
rect 286799 212600 286800 213000
rect 287200 212600 287201 213000
rect 286799 212599 287201 212600
rect 287599 213000 288001 213001
rect 287599 212600 287600 213000
rect 288000 212600 288001 213000
rect 287599 212599 288001 212600
rect 288399 213000 288801 213001
rect 288399 212600 288400 213000
rect 288800 212600 288801 213000
rect 288399 212599 288801 212600
rect 289199 213000 289601 213001
rect 289199 212600 289200 213000
rect 289600 212600 289601 213000
rect 289199 212599 289601 212600
rect 285199 212200 285601 212201
rect 285199 211800 285200 212200
rect 285600 211800 285601 212200
rect 285199 211799 285601 211800
rect 285999 212200 286401 212201
rect 285999 211800 286000 212200
rect 286400 211800 286401 212200
rect 285999 211799 286401 211800
rect 286799 212200 287201 212201
rect 286799 211800 286800 212200
rect 287200 211800 287201 212200
rect 286799 211799 287201 211800
rect 287599 212200 288001 212201
rect 287599 211800 287600 212200
rect 288000 211800 288001 212200
rect 287599 211799 288001 211800
rect 288399 212200 288801 212201
rect 288399 211800 288400 212200
rect 288800 211800 288801 212200
rect 288399 211799 288801 211800
rect 289199 212200 289601 212201
rect 289199 211800 289200 212200
rect 289600 211800 289601 212200
rect 289199 211799 289601 211800
rect 285199 211400 285601 211401
rect 285199 211000 285200 211400
rect 285600 211000 285601 211400
rect 285199 210999 285601 211000
rect 285999 211400 286401 211401
rect 285999 211000 286000 211400
rect 286400 211000 286401 211400
rect 285999 210999 286401 211000
rect 286799 211400 287201 211401
rect 286799 211000 286800 211400
rect 287200 211000 287201 211400
rect 286799 210999 287201 211000
rect 287599 211400 288001 211401
rect 287599 211000 287600 211400
rect 288000 211000 288001 211400
rect 287599 210999 288001 211000
rect 288399 211400 288801 211401
rect 288399 211000 288400 211400
rect 288800 211000 288801 211400
rect 288399 210999 288801 211000
rect 289199 211400 289601 211401
rect 289199 211000 289200 211400
rect 289600 211000 289601 211400
rect 289199 210999 289601 211000
rect 285199 210600 285601 210601
rect 285199 210200 285200 210600
rect 285600 210200 285601 210600
rect 285199 210199 285601 210200
rect 285999 210600 286401 210601
rect 285999 210200 286000 210600
rect 286400 210200 286401 210600
rect 285999 210199 286401 210200
rect 286799 210600 287201 210601
rect 286799 210200 286800 210600
rect 287200 210200 287201 210600
rect 286799 210199 287201 210200
rect 287599 210600 288001 210601
rect 287599 210200 287600 210600
rect 288000 210200 288001 210600
rect 287599 210199 288001 210200
rect 288399 210600 288801 210601
rect 288399 210200 288400 210600
rect 288800 210200 288801 210600
rect 288399 210199 288801 210200
rect 289199 210600 289601 210601
rect 289199 210200 289200 210600
rect 289600 210200 289601 210600
rect 289199 210199 289601 210200
rect 285199 209800 285601 209801
rect 285199 209400 285200 209800
rect 285600 209400 285601 209800
rect 285199 209399 285601 209400
rect 285999 209800 286401 209801
rect 285999 209400 286000 209800
rect 286400 209400 286401 209800
rect 285999 209399 286401 209400
rect 286799 209800 287201 209801
rect 286799 209400 286800 209800
rect 287200 209400 287201 209800
rect 286799 209399 287201 209400
rect 287599 209800 288001 209801
rect 287599 209400 287600 209800
rect 288000 209400 288001 209800
rect 287599 209399 288001 209400
rect 288399 209800 288801 209801
rect 288399 209400 288400 209800
rect 288800 209400 288801 209800
rect 288399 209399 288801 209400
rect 289199 209800 289601 209801
rect 289199 209400 289200 209800
rect 289600 209400 289601 209800
rect 289199 209399 289601 209400
rect 285199 209000 285601 209001
rect 285199 208600 285200 209000
rect 285600 208600 285601 209000
rect 285199 208599 285601 208600
rect 285999 209000 286401 209001
rect 285999 208600 286000 209000
rect 286400 208600 286401 209000
rect 285999 208599 286401 208600
rect 286799 209000 287201 209001
rect 286799 208600 286800 209000
rect 287200 208600 287201 209000
rect 286799 208599 287201 208600
rect 287599 209000 288001 209001
rect 287599 208600 287600 209000
rect 288000 208600 288001 209000
rect 287599 208599 288001 208600
rect 288399 209000 288801 209001
rect 288399 208600 288400 209000
rect 288800 208600 288801 209000
rect 288399 208599 288801 208600
rect 289199 209000 289601 209001
rect 289199 208600 289200 209000
rect 289600 208600 289601 209000
rect 289199 208599 289601 208600
rect 285199 208200 285601 208201
rect 285199 207800 285200 208200
rect 285600 207800 285601 208200
rect 285199 207799 285601 207800
rect 285999 208200 286401 208201
rect 285999 207800 286000 208200
rect 286400 207800 286401 208200
rect 285999 207799 286401 207800
rect 286799 208200 287201 208201
rect 286799 207800 286800 208200
rect 287200 207800 287201 208200
rect 286799 207799 287201 207800
rect 287599 208200 288001 208201
rect 287599 207800 287600 208200
rect 288000 207800 288001 208200
rect 287599 207799 288001 207800
rect 288399 208200 288801 208201
rect 288399 207800 288400 208200
rect 288800 207800 288801 208200
rect 288399 207799 288801 207800
rect 289199 208200 289601 208201
rect 289199 207800 289200 208200
rect 289600 207800 289601 208200
rect 289199 207799 289601 207800
rect 285199 207400 285601 207401
rect 285199 207000 285200 207400
rect 285600 207000 285601 207400
rect 285199 206999 285601 207000
rect 285999 207400 286401 207401
rect 285999 207000 286000 207400
rect 286400 207000 286401 207400
rect 285999 206999 286401 207000
rect 286799 207400 287201 207401
rect 286799 207000 286800 207400
rect 287200 207000 287201 207400
rect 286799 206999 287201 207000
rect 287599 207400 288001 207401
rect 287599 207000 287600 207400
rect 288000 207000 288001 207400
rect 287599 206999 288001 207000
rect 288399 207400 288801 207401
rect 288399 207000 288400 207400
rect 288800 207000 288801 207400
rect 288399 206999 288801 207000
rect 289199 207400 289601 207401
rect 289199 207000 289200 207400
rect 289600 207000 289601 207400
rect 289199 206999 289601 207000
rect 285199 206600 285601 206601
rect 285199 206200 285200 206600
rect 285600 206200 285601 206600
rect 285199 206199 285601 206200
rect 285999 206600 286401 206601
rect 285999 206200 286000 206600
rect 286400 206200 286401 206600
rect 285999 206199 286401 206200
rect 286799 206600 287201 206601
rect 286799 206200 286800 206600
rect 287200 206200 287201 206600
rect 286799 206199 287201 206200
rect 287599 206600 288001 206601
rect 287599 206200 287600 206600
rect 288000 206200 288001 206600
rect 287599 206199 288001 206200
rect 288399 206600 288801 206601
rect 288399 206200 288400 206600
rect 288800 206200 288801 206600
rect 288399 206199 288801 206200
rect 289199 206600 289601 206601
rect 289199 206200 289200 206600
rect 289600 206200 289601 206600
rect 289199 206199 289601 206200
rect 285199 205800 285601 205801
rect 285199 205400 285200 205800
rect 285600 205400 285601 205800
rect 285199 205399 285601 205400
rect 285999 205800 286401 205801
rect 285999 205400 286000 205800
rect 286400 205400 286401 205800
rect 285999 205399 286401 205400
rect 286799 205800 287201 205801
rect 286799 205400 286800 205800
rect 287200 205400 287201 205800
rect 286799 205399 287201 205400
rect 287599 205800 288001 205801
rect 287599 205400 287600 205800
rect 288000 205400 288001 205800
rect 287599 205399 288001 205400
rect 288399 205800 288801 205801
rect 288399 205400 288400 205800
rect 288800 205400 288801 205800
rect 288399 205399 288801 205400
rect 289199 205800 289601 205801
rect 289199 205400 289200 205800
rect 289600 205400 289601 205800
rect 289199 205399 289601 205400
rect 83800 177200 86000 177600
rect 86400 177200 86800 177600
rect 87200 177200 87600 177600
rect 88000 177200 88400 177600
rect 88800 177200 89200 177600
rect 89600 177200 90000 177600
rect 90400 177200 92000 177600
rect 83800 176800 92000 177200
rect 83800 176400 86000 176800
rect 86400 176400 86800 176800
rect 87200 176400 87600 176800
rect 88000 176400 88400 176800
rect 88800 176400 89200 176800
rect 89600 176400 90000 176800
rect 90400 176400 92000 176800
rect 83800 176000 92000 176400
rect 83800 175600 86000 176000
rect 86400 175600 86800 176000
rect 87200 175600 87600 176000
rect 88000 175600 88400 176000
rect 88800 175600 89200 176000
rect 89600 175600 90000 176000
rect 90400 175600 92000 176000
rect 83800 175200 92000 175600
rect 83800 174800 86000 175200
rect 86400 174800 86800 175200
rect 87200 174800 87600 175200
rect 88000 174800 88400 175200
rect 88800 174800 89200 175200
rect 89600 174800 90000 175200
rect 90400 174800 92000 175200
rect 83800 174400 92000 174800
rect 83800 174000 86000 174400
rect 86400 174000 86800 174400
rect 87200 174000 87600 174400
rect 88000 174000 88400 174400
rect 88800 174000 89200 174400
rect 89600 174000 90000 174400
rect 90400 174000 92000 174400
rect 83800 173600 92000 174000
rect 83800 173200 86000 173600
rect 86400 173200 86800 173600
rect 87200 173200 87600 173600
rect 88000 173200 88400 173600
rect 88800 173200 89200 173600
rect 89600 173200 90000 173600
rect 90400 173200 92000 173600
rect 83800 172800 92000 173200
rect 83800 172400 86000 172800
rect 86400 172400 86800 172800
rect 87200 172400 87600 172800
rect 88000 172400 88400 172800
rect 88800 172400 89200 172800
rect 89600 172400 90000 172800
rect 90400 172400 92000 172800
rect 83800 172000 92000 172400
rect 83800 171600 86000 172000
rect 86400 171600 86800 172000
rect 87200 171600 87600 172000
rect 88000 171600 88400 172000
rect 88800 171600 89200 172000
rect 89600 171600 90000 172000
rect 90400 171600 92000 172000
rect 83800 171200 92000 171600
rect 83800 170800 86000 171200
rect 86400 170800 86800 171200
rect 87200 170800 87600 171200
rect 88000 170800 88400 171200
rect 88800 170800 89200 171200
rect 89600 170800 90000 171200
rect 90400 170800 92000 171200
rect 83800 170400 92000 170800
rect 83800 170000 86000 170400
rect 86400 170000 86800 170400
rect 87200 170000 87600 170400
rect 88000 170000 88400 170400
rect 88800 170000 89200 170400
rect 89600 170000 90000 170400
rect 90400 170000 92000 170400
rect 83800 169600 92000 170000
rect 83800 169200 86000 169600
rect 86400 169200 86800 169600
rect 87200 169200 87600 169600
rect 88000 169200 88400 169600
rect 88800 169200 89200 169600
rect 89600 169200 90000 169600
rect 90400 169200 92000 169600
rect 83800 168800 92000 169200
rect 83800 168400 86000 168800
rect 86400 168400 86800 168800
rect 87200 168400 87600 168800
rect 88000 168400 88400 168800
rect 88800 168400 89200 168800
rect 89600 168400 90000 168800
rect 90400 168400 92000 168800
rect 83800 168000 92000 168400
rect 83800 167600 86000 168000
rect 86400 167600 86800 168000
rect 87200 167600 87600 168000
rect 88000 167600 88400 168000
rect 88800 167600 89200 168000
rect 89600 167600 90000 168000
rect 90400 167600 92000 168000
rect 83800 167200 92000 167600
rect 83800 166800 86000 167200
rect 86400 166800 86800 167200
rect 87200 166800 87600 167200
rect 88000 166800 88400 167200
rect 88800 166800 89200 167200
rect 89600 166800 90000 167200
rect 90400 166800 92000 167200
rect 83800 166400 92000 166800
rect 83800 166000 86000 166400
rect 86400 166000 86800 166400
rect 87200 166000 87600 166400
rect 88000 166000 88400 166400
rect 88800 166000 89200 166400
rect 89600 166000 90000 166400
rect 90400 166000 92000 166400
rect 83800 165600 92000 166000
rect 83800 165200 86000 165600
rect 86400 165200 86800 165600
rect 87200 165200 87600 165600
rect 88000 165200 88400 165600
rect 88800 165200 89200 165600
rect 89600 165200 90000 165600
rect 90400 165200 92000 165600
rect 83800 164800 92000 165200
rect 83800 164400 86000 164800
rect 86400 164400 86800 164800
rect 87200 164400 87600 164800
rect 88000 164400 88400 164800
rect 88800 164400 89200 164800
rect 89600 164400 90000 164800
rect 90400 164400 92000 164800
rect 83800 164000 92000 164400
rect 83800 163600 86000 164000
rect 86400 163600 86800 164000
rect 87200 163600 87600 164000
rect 88000 163600 88400 164000
rect 88800 163600 89200 164000
rect 89600 163600 90000 164000
rect 90400 163600 92000 164000
rect 83800 162900 92000 163600
rect 297000 177600 306000 343300
rect 569100 302000 570220 302200
rect 569100 301800 569300 302000
rect 569500 301800 569800 302000
rect 570000 301800 570220 302000
rect 569100 301600 570220 301800
rect 511500 301400 517000 301600
rect 511500 301200 511700 301400
rect 511900 301200 512100 301400
rect 512300 301200 512500 301400
rect 512700 301200 512900 301400
rect 513100 301200 513300 301400
rect 513500 301200 513700 301400
rect 513900 301200 514100 301400
rect 514300 301200 514500 301400
rect 514700 301200 514900 301400
rect 515100 301200 515300 301400
rect 515500 301200 515700 301400
rect 515900 301200 516100 301400
rect 516300 301200 516500 301400
rect 516700 301200 517000 301400
rect 511500 301000 517000 301200
rect 511500 300800 511700 301000
rect 511900 300800 512100 301000
rect 512300 300800 512500 301000
rect 512700 300800 512900 301000
rect 513100 300800 513300 301000
rect 513500 300800 513700 301000
rect 513900 300800 514100 301000
rect 514300 300800 514500 301000
rect 514700 300800 514900 301000
rect 515100 300800 515300 301000
rect 515500 300800 515700 301000
rect 515900 300800 516100 301000
rect 516300 300800 516500 301000
rect 516700 300800 517000 301000
rect 511500 300600 517000 300800
rect 511500 300400 511700 300600
rect 511900 300400 512100 300600
rect 512300 300400 512500 300600
rect 512700 300400 512900 300600
rect 513100 300400 513300 300600
rect 513500 300400 513700 300600
rect 513900 300400 514100 300600
rect 514300 300400 514500 300600
rect 514700 300400 514900 300600
rect 515100 300400 515300 300600
rect 515500 300400 515700 300600
rect 515900 300400 516100 300600
rect 516300 300400 516500 300600
rect 516700 300400 517000 300600
rect 511500 288800 517000 300400
rect 569100 301400 569300 301600
rect 569500 301400 569800 301600
rect 570000 301400 570220 301600
rect 569100 301200 570220 301400
rect 569100 301000 569300 301200
rect 569500 301000 569800 301200
rect 570000 301000 570220 301200
rect 569100 300800 570220 301000
rect 569100 300600 569300 300800
rect 569500 300600 569800 300800
rect 570000 300600 570220 300800
rect 569100 300400 570220 300600
rect 569100 300200 569300 300400
rect 569500 300200 569800 300400
rect 570000 300200 570220 300400
rect 530599 298992 550539 299052
rect 530599 298862 530639 298992
rect 530739 298862 530899 298992
rect 530999 298921 550129 298992
rect 530999 298862 533197 298921
rect 530599 298857 533197 298862
rect 536541 298857 536997 298921
rect 540341 298857 540797 298921
rect 544141 298857 544597 298921
rect 547941 298862 550129 298921
rect 550239 298862 550389 298992
rect 550499 298862 550539 298992
rect 547941 298857 550539 298862
rect 530599 298812 550539 298857
rect 533308 298702 536430 298703
rect 533308 295582 533309 298702
rect 536429 297552 536430 298702
rect 537108 298702 540230 298703
rect 537108 297552 537109 298702
rect 536429 297192 537109 297552
rect 536429 295582 536430 297192
rect 533308 295581 536430 295582
rect 536649 295372 536819 297192
rect 537108 295582 537109 297192
rect 540229 297552 540230 298702
rect 540908 298702 544030 298703
rect 540908 297552 540909 298702
rect 540229 297192 540909 297552
rect 540229 295582 540230 297192
rect 537108 295581 540230 295582
rect 540908 295582 540909 297192
rect 544029 297552 544030 298702
rect 544708 298702 547830 298703
rect 544708 297552 544709 298702
rect 544029 297192 544709 297552
rect 544029 295582 544030 297192
rect 540908 295581 544030 295582
rect 534849 295182 536819 295372
rect 544289 295392 544449 297192
rect 544708 295582 544709 297192
rect 547829 295582 547830 298702
rect 544708 295581 547830 295582
rect 544289 295262 545069 295392
rect 534849 294500 535139 295182
rect 537069 294682 537339 294812
rect 537069 294602 537089 294682
rect 537169 294602 537239 294682
rect 537319 294602 537339 294682
rect 528200 294400 535200 294500
rect 528200 294200 528300 294400
rect 528500 294200 528700 294400
rect 528900 294200 529100 294400
rect 529300 294200 529500 294400
rect 529700 294200 529900 294400
rect 530100 294200 535200 294400
rect 528200 294100 535200 294200
rect 528200 293900 528300 294100
rect 528500 293900 528700 294100
rect 528900 293900 529100 294100
rect 529300 293900 529500 294100
rect 529700 293900 529900 294100
rect 530100 293900 535200 294100
rect 528200 293700 535200 293900
rect 528200 293500 528300 293700
rect 528500 293500 528700 293700
rect 528900 293500 529100 293700
rect 529300 293500 529500 293700
rect 529700 293500 529900 293700
rect 530100 293500 535200 293700
rect 528200 293300 535200 293500
rect 528200 293100 528300 293300
rect 528500 293100 528700 293300
rect 528900 293100 529100 293300
rect 529300 293100 529500 293300
rect 529700 293100 529900 293300
rect 530100 293100 535200 293300
rect 528200 292900 535200 293100
rect 528200 292700 528300 292900
rect 528500 292700 528700 292900
rect 528900 292700 529100 292900
rect 529300 292700 529500 292900
rect 529700 292700 529900 292900
rect 530100 292700 535200 292900
rect 528200 292600 535200 292700
rect 537069 294142 537339 294602
rect 537069 294062 537089 294142
rect 537169 294062 537239 294142
rect 537319 294062 537339 294142
rect 537069 293602 537339 294062
rect 537069 293522 537089 293602
rect 537169 293522 537239 293602
rect 537319 293522 537339 293602
rect 534849 291652 535139 292600
rect 534849 291542 534869 291652
rect 534959 291542 535029 291652
rect 535119 291542 535139 291652
rect 534849 291322 535139 291542
rect 511500 288600 511700 288800
rect 511900 288600 512100 288800
rect 512300 288600 512500 288800
rect 512700 288600 512900 288800
rect 513100 288600 513300 288800
rect 513500 288600 513700 288800
rect 513900 288600 514100 288800
rect 514300 288600 514500 288800
rect 514700 288600 514900 288800
rect 515100 288600 515300 288800
rect 515500 288600 515700 288800
rect 515900 288600 516100 288800
rect 516300 288600 516500 288800
rect 516700 288600 517000 288800
rect 511500 288400 517000 288600
rect 511500 288200 511700 288400
rect 511900 288200 512100 288400
rect 512300 288200 512500 288400
rect 512700 288200 512900 288400
rect 513100 288200 513300 288400
rect 513500 288200 513700 288400
rect 513900 288200 514100 288400
rect 514300 288200 514500 288400
rect 514700 288200 514900 288400
rect 515100 288200 515300 288400
rect 515500 288200 515700 288400
rect 515900 288200 516100 288400
rect 516300 288200 516500 288400
rect 516700 288200 517000 288400
rect 537069 288372 537339 293522
rect 539559 294682 539829 294862
rect 539559 294602 539579 294682
rect 539659 294602 539729 294682
rect 539809 294602 539829 294682
rect 539559 294142 539829 294602
rect 539559 294062 539579 294142
rect 539659 294062 539729 294142
rect 539809 294062 539829 294142
rect 539559 293602 539829 294062
rect 539559 293522 539579 293602
rect 539659 293522 539729 293602
rect 539809 293522 539829 293602
rect 538359 293002 538589 293022
rect 538359 292922 538379 293002
rect 538459 292922 538489 293002
rect 538569 292922 538589 293002
rect 538359 292392 538589 292922
rect 538359 292312 538379 292392
rect 538459 292312 538489 292392
rect 538569 292312 538589 292392
rect 538359 291832 538589 292312
rect 538359 291752 538379 291832
rect 538459 291752 538489 291832
rect 538569 291752 538589 291832
rect 538359 289132 538589 291752
rect 538359 289052 538379 289132
rect 538459 289052 538489 289132
rect 538569 289052 538589 289132
rect 538359 289032 538589 289052
rect 537069 288292 537089 288372
rect 537169 288292 537239 288372
rect 537319 288292 537339 288372
rect 539559 288392 539829 293522
rect 542039 294682 542309 294872
rect 542039 294602 542059 294682
rect 542139 294602 542209 294682
rect 542289 294602 542309 294682
rect 542039 294142 542309 294602
rect 542039 294062 542059 294142
rect 542139 294062 542209 294142
rect 542289 294062 542309 294142
rect 542039 293602 542309 294062
rect 542039 293522 542069 293602
rect 542149 293522 542209 293602
rect 542289 293522 542309 293602
rect 540769 293002 540999 293022
rect 540769 292922 540789 293002
rect 540869 292922 540899 293002
rect 540979 292922 540999 293002
rect 540769 292412 540999 292922
rect 540769 292332 540789 292412
rect 540869 292332 540899 292412
rect 540979 292332 540999 292412
rect 540769 291832 540999 292332
rect 540769 291752 540789 291832
rect 540869 291752 540899 291832
rect 540979 291752 540999 291832
rect 540769 289132 540999 291752
rect 540769 289052 540789 289132
rect 540869 289052 540899 289132
rect 540979 289052 540999 289132
rect 540769 289032 540999 289052
rect 539559 288312 539579 288392
rect 539659 288312 539729 288392
rect 539809 288312 539829 288392
rect 539559 288292 539829 288312
rect 542039 288392 542309 293522
rect 543229 292992 543459 293032
rect 543229 292912 543249 292992
rect 543329 292912 543359 292992
rect 543439 292912 543459 292992
rect 543229 292412 543459 292912
rect 543229 292332 543249 292412
rect 543329 292332 543359 292412
rect 543439 292332 543459 292412
rect 543229 291832 543459 292332
rect 543229 291752 543249 291832
rect 543329 291752 543359 291832
rect 543439 291752 543459 291832
rect 543229 289142 543459 291752
rect 544779 291602 545069 295262
rect 544779 291522 544799 291602
rect 544879 291522 544969 291602
rect 545049 291522 545069 291602
rect 544779 291112 545069 291522
rect 545700 291300 549100 291400
rect 545700 291200 547200 291300
rect 543229 289062 543249 289142
rect 543329 289062 543359 289142
rect 543439 289062 543459 289142
rect 543229 289042 543459 289062
rect 545700 291000 545900 291200
rect 546100 291000 546200 291200
rect 546400 291000 546500 291200
rect 546700 291000 546800 291200
rect 547000 291100 547200 291200
rect 547400 291100 549100 291300
rect 547000 291000 549100 291100
rect 545700 290800 547200 291000
rect 547400 290800 549100 291000
rect 545700 290700 549100 290800
rect 545700 290500 547200 290700
rect 547400 290500 549100 290700
rect 545700 290400 549100 290500
rect 545700 290200 547200 290400
rect 547400 290200 549100 290400
rect 545700 290100 549100 290200
rect 545700 289900 545800 290100
rect 546000 289900 546100 290100
rect 546300 289900 546400 290100
rect 546600 289900 546800 290100
rect 547000 289900 549100 290100
rect 542039 288312 542059 288392
rect 542139 288312 542199 288392
rect 542279 288312 542309 288392
rect 542039 288292 542309 288312
rect 545700 288900 549100 289900
rect 545700 288600 545900 288900
rect 546200 288600 546400 288900
rect 546700 288600 546900 288900
rect 547200 288600 547400 288900
rect 547700 288600 547900 288900
rect 548200 288600 548400 288900
rect 548700 288600 549100 288900
rect 545700 288400 549100 288600
rect 537069 288262 537339 288292
rect 511500 288000 517000 288200
rect 511500 287800 511700 288000
rect 511900 287800 512100 288000
rect 512300 287800 512500 288000
rect 512700 287800 512900 288000
rect 513100 287800 513300 288000
rect 513500 287800 513700 288000
rect 513900 287800 514100 288000
rect 514300 287800 514500 288000
rect 514700 287800 514900 288000
rect 515100 287800 515300 288000
rect 515500 287800 515700 288000
rect 515900 287800 516100 288000
rect 516300 287800 516500 288000
rect 516700 287800 517000 288000
rect 511500 287600 517000 287800
rect 511500 287400 511700 287600
rect 511900 287400 512100 287600
rect 512300 287400 512500 287600
rect 512700 287400 512900 287600
rect 513100 287400 513300 287600
rect 513500 287400 513700 287600
rect 513900 287400 514100 287600
rect 514300 287400 514500 287600
rect 514700 287400 514900 287600
rect 515100 287400 515300 287600
rect 515500 287400 515700 287600
rect 515900 287400 516100 287600
rect 516300 287400 516500 287600
rect 516700 287400 517000 287600
rect 511500 287200 517000 287400
rect 511500 287000 511700 287200
rect 511900 287000 512100 287200
rect 512300 287000 512500 287200
rect 512700 287000 512900 287200
rect 513100 287000 513300 287200
rect 513500 287000 513700 287200
rect 513900 287000 514100 287200
rect 514300 287000 514500 287200
rect 514700 287000 514900 287200
rect 515100 287000 515300 287200
rect 515500 287000 515700 287200
rect 515900 287000 516100 287200
rect 516300 287000 516500 287200
rect 516700 287000 517000 287200
rect 511500 286800 517000 287000
rect 511500 286600 511700 286800
rect 511900 286600 512100 286800
rect 512300 286600 512500 286800
rect 512700 286600 512900 286800
rect 513100 286600 513300 286800
rect 513500 286600 513700 286800
rect 513900 286600 514100 286800
rect 514300 286600 514500 286800
rect 514700 286600 514900 286800
rect 515100 286600 515300 286800
rect 515500 286600 515700 286800
rect 515900 286600 516100 286800
rect 516300 286600 516500 286800
rect 516700 286600 517000 286800
rect 511500 283200 517000 286600
rect 545700 288100 545900 288400
rect 546200 288100 546400 288400
rect 546700 288100 546900 288400
rect 547200 288100 547400 288400
rect 547700 288100 547900 288400
rect 548200 288100 548400 288400
rect 548700 288100 549100 288400
rect 545700 287900 549100 288100
rect 545700 287600 545900 287900
rect 546200 287600 546400 287900
rect 546700 287600 546900 287900
rect 547200 287600 547400 287900
rect 547700 287600 547900 287900
rect 548200 287600 548400 287900
rect 548700 287600 549100 287900
rect 542388 286442 542510 286443
rect 542388 286342 542389 286442
rect 542509 286342 542510 286442
rect 542388 286341 542510 286342
rect 511500 283000 511900 283200
rect 512100 283000 512300 283200
rect 512500 283000 512700 283200
rect 512900 283000 513100 283200
rect 513300 283000 513500 283200
rect 513700 283000 513900 283200
rect 514100 283000 514300 283200
rect 514500 283000 514700 283200
rect 514900 283000 515100 283200
rect 515300 283000 515500 283200
rect 515700 283000 515900 283200
rect 516100 283000 516300 283200
rect 516500 283000 516700 283200
rect 516900 283000 517000 283200
rect 511500 282800 517000 283000
rect 511500 282600 511900 282800
rect 512100 282600 512300 282800
rect 512500 282600 512700 282800
rect 512900 282600 513100 282800
rect 513300 282600 513500 282800
rect 513700 282600 513900 282800
rect 514100 282600 514300 282800
rect 514500 282600 514700 282800
rect 514900 282600 515100 282800
rect 515300 282600 515500 282800
rect 515700 282600 515900 282800
rect 516100 282600 516300 282800
rect 516500 282600 516700 282800
rect 516900 282600 517000 282800
rect 511500 282400 517000 282600
rect 511500 282200 511900 282400
rect 512100 282200 512300 282400
rect 512500 282200 512700 282400
rect 512900 282200 513100 282400
rect 513300 282200 513500 282400
rect 513700 282200 513900 282400
rect 514100 282200 514300 282400
rect 514500 282200 514700 282400
rect 514900 282200 515100 282400
rect 515300 282200 515500 282400
rect 515700 282200 515900 282400
rect 516100 282200 516300 282400
rect 516500 282200 516700 282400
rect 516900 282200 517000 282400
rect 511500 282000 517000 282200
rect 511500 281800 511900 282000
rect 512100 281800 512300 282000
rect 512500 281800 512700 282000
rect 512900 281800 513100 282000
rect 513300 281800 513500 282000
rect 513700 281800 513900 282000
rect 514100 281800 514300 282000
rect 514500 281800 514700 282000
rect 514900 281800 515100 282000
rect 515300 281800 515500 282000
rect 515700 281800 515900 282000
rect 516100 281800 516300 282000
rect 516500 281800 516700 282000
rect 516900 281800 517000 282000
rect 511500 281600 517000 281800
rect 511500 281400 511900 281600
rect 512100 281400 512300 281600
rect 512500 281400 512700 281600
rect 512900 281400 513100 281600
rect 513300 281400 513500 281600
rect 513700 281400 513900 281600
rect 514100 281400 514300 281600
rect 514500 281400 514700 281600
rect 514900 281400 515100 281600
rect 515300 281400 515500 281600
rect 515700 281400 515900 281600
rect 516100 281400 516300 281600
rect 516500 281400 516700 281600
rect 516900 281400 517000 281600
rect 511500 281200 517000 281400
rect 511500 281000 511900 281200
rect 512100 281000 512300 281200
rect 512500 281000 512700 281200
rect 512900 281000 513100 281200
rect 513300 281000 513500 281200
rect 513700 281000 513900 281200
rect 514100 281000 514300 281200
rect 514500 281000 514700 281200
rect 514900 281000 515100 281200
rect 515300 281000 515500 281200
rect 515700 281000 515900 281200
rect 516100 281000 516300 281200
rect 516500 281000 516700 281200
rect 516900 281000 517000 281200
rect 511500 280800 517000 281000
rect 511500 280600 511900 280800
rect 512100 280600 512300 280800
rect 512500 280600 512700 280800
rect 512900 280600 513100 280800
rect 513300 280600 513500 280800
rect 513700 280600 513900 280800
rect 514100 280600 514300 280800
rect 514500 280600 514700 280800
rect 514900 280600 515100 280800
rect 515300 280600 515500 280800
rect 515700 280600 515900 280800
rect 516100 280600 516300 280800
rect 516500 280600 516700 280800
rect 516900 280600 517000 280800
rect 511500 195600 517000 280600
rect 545700 285400 549100 287600
rect 569100 288900 570220 300200
rect 569100 288600 569200 288900
rect 569500 288600 569800 288900
rect 570100 288600 570220 288900
rect 569100 288400 570220 288600
rect 569100 288100 569200 288400
rect 569500 288100 569800 288400
rect 570100 288100 570220 288400
rect 572799 288700 573101 288701
rect 572799 288400 572800 288700
rect 573100 288400 573101 288700
rect 572799 288399 573101 288400
rect 573299 288700 573601 288701
rect 573299 288400 573300 288700
rect 573600 288400 573601 288700
rect 573299 288399 573601 288400
rect 573799 288700 574101 288701
rect 573799 288400 573800 288700
rect 574100 288400 574101 288700
rect 573799 288399 574101 288400
rect 574299 288700 574601 288701
rect 574299 288400 574300 288700
rect 574600 288400 574601 288700
rect 574299 288399 574601 288400
rect 569100 287900 570220 288100
rect 569100 287600 569200 287900
rect 569500 287600 569800 287900
rect 570100 287600 570220 287900
rect 572799 288200 573101 288201
rect 572799 287900 572800 288200
rect 573100 287900 573101 288200
rect 572799 287899 573101 287900
rect 573299 288200 573601 288201
rect 573299 287900 573300 288200
rect 573600 287900 573601 288200
rect 573299 287899 573601 287900
rect 573799 288200 574101 288201
rect 573799 287900 573800 288200
rect 574100 287900 574101 288200
rect 573799 287899 574101 287900
rect 574299 288200 574601 288201
rect 574299 287900 574300 288200
rect 574600 287900 574601 288200
rect 574299 287899 574601 287900
rect 569100 287400 570220 287600
rect 545700 285200 545800 285400
rect 546000 285200 546200 285400
rect 546400 285200 546600 285400
rect 546800 285200 547000 285400
rect 547200 285200 547400 285400
rect 547600 285200 547800 285400
rect 548000 285200 548200 285400
rect 548400 285200 548600 285400
rect 548800 285200 549100 285400
rect 545700 285000 549100 285200
rect 545700 284800 545800 285000
rect 546000 284800 546200 285000
rect 546400 284800 546600 285000
rect 546800 284800 547000 285000
rect 547200 284800 547400 285000
rect 547600 284800 547800 285000
rect 548000 284800 548200 285000
rect 548400 284800 548600 285000
rect 548800 284800 549100 285000
rect 545700 248600 549100 284800
rect 545700 248400 546000 248600
rect 546200 248400 546400 248600
rect 546600 248400 546800 248600
rect 547000 248400 547200 248600
rect 547400 248400 547600 248600
rect 547800 248400 548000 248600
rect 548200 248400 548400 248600
rect 548600 248400 548800 248600
rect 549000 248400 549100 248600
rect 545700 248200 549100 248400
rect 545700 248000 546000 248200
rect 546200 248000 546400 248200
rect 546600 248000 546800 248200
rect 547000 248000 547200 248200
rect 547400 248000 547600 248200
rect 547800 248000 548000 248200
rect 548200 248000 548400 248200
rect 548600 248000 548800 248200
rect 549000 248000 549100 248200
rect 545700 247800 549100 248000
rect 545700 247600 546000 247800
rect 546200 247600 546400 247800
rect 546600 247600 546800 247800
rect 547000 247600 547200 247800
rect 547400 247600 547600 247800
rect 547800 247600 548000 247800
rect 548200 247600 548400 247800
rect 548600 247600 548800 247800
rect 549000 247600 549100 247800
rect 545700 247400 549100 247600
rect 545700 247200 546000 247400
rect 546200 247200 546400 247400
rect 546600 247200 546800 247400
rect 547000 247200 547200 247400
rect 547400 247200 547600 247400
rect 547800 247200 548000 247400
rect 548200 247200 548400 247400
rect 548600 247200 548800 247400
rect 549000 247200 549100 247400
rect 545700 247000 549100 247200
rect 545700 246800 546000 247000
rect 546200 246800 546400 247000
rect 546600 246800 546800 247000
rect 547000 246800 547200 247000
rect 547400 246800 547600 247000
rect 547800 246800 548000 247000
rect 548200 246800 548400 247000
rect 548600 246800 548800 247000
rect 549000 246800 549100 247000
rect 545700 246600 549100 246800
rect 545700 246400 546000 246600
rect 546200 246400 546400 246600
rect 546600 246400 546800 246600
rect 547000 246400 547200 246600
rect 547400 246400 547600 246600
rect 547800 246400 548000 246600
rect 548200 246400 548400 246600
rect 548600 246400 548800 246600
rect 549000 246400 549100 246600
rect 545700 246200 549100 246400
rect 545700 246000 546000 246200
rect 546200 246000 546400 246200
rect 546600 246000 546800 246200
rect 547000 246000 547200 246200
rect 547400 246000 547600 246200
rect 547800 246000 548000 246200
rect 548200 246000 548400 246200
rect 548600 246000 548800 246200
rect 549000 246000 549100 246200
rect 545700 245800 549100 246000
rect 545700 245600 546000 245800
rect 546200 245600 546400 245800
rect 546600 245600 546800 245800
rect 547000 245600 547200 245800
rect 547400 245600 547600 245800
rect 547800 245600 548000 245800
rect 548200 245600 548400 245800
rect 548600 245600 548800 245800
rect 549000 245600 549100 245800
rect 545700 245400 549100 245600
rect 545700 245200 546000 245400
rect 546200 245200 546400 245400
rect 546600 245200 546800 245400
rect 547000 245200 547200 245400
rect 547400 245200 547600 245400
rect 547800 245200 548000 245400
rect 548200 245200 548400 245400
rect 548600 245200 548800 245400
rect 549000 245200 549100 245400
rect 545700 245000 549100 245200
rect 545700 244800 546000 245000
rect 546200 244800 546400 245000
rect 546600 244800 546800 245000
rect 547000 244800 547200 245000
rect 547400 244800 547600 245000
rect 547800 244800 548000 245000
rect 548200 244800 548400 245000
rect 548600 244800 548800 245000
rect 549000 244800 549100 245000
rect 545700 244600 549100 244800
rect 545700 244400 546000 244600
rect 546200 244400 546400 244600
rect 546600 244400 546800 244600
rect 547000 244400 547200 244600
rect 547400 244400 547600 244600
rect 547800 244400 548000 244600
rect 548200 244400 548400 244600
rect 548600 244400 548800 244600
rect 549000 244400 549100 244600
rect 545700 244200 549100 244400
rect 545700 244000 546000 244200
rect 546200 244000 546400 244200
rect 546600 244000 546800 244200
rect 547000 244000 547200 244200
rect 547400 244000 547600 244200
rect 547800 244000 548000 244200
rect 548200 244000 548400 244200
rect 548600 244000 548800 244200
rect 549000 244000 549100 244200
rect 545700 243800 549100 244000
rect 545700 243600 546000 243800
rect 546200 243600 546400 243800
rect 546600 243600 546800 243800
rect 547000 243600 547200 243800
rect 547400 243600 547600 243800
rect 547800 243600 548000 243800
rect 548200 243600 548400 243800
rect 548600 243600 548800 243800
rect 549000 243600 549100 243800
rect 545700 243400 549100 243600
rect 545700 243200 546000 243400
rect 546200 243200 546400 243400
rect 546600 243200 546800 243400
rect 547000 243200 547200 243400
rect 547400 243200 547600 243400
rect 547800 243200 548000 243400
rect 548200 243200 548400 243400
rect 548600 243200 548800 243400
rect 549000 243200 549100 243400
rect 545700 243000 549100 243200
rect 545700 242800 546000 243000
rect 546200 242800 546400 243000
rect 546600 242800 546800 243000
rect 547000 242800 547200 243000
rect 547400 242800 547600 243000
rect 547800 242800 548000 243000
rect 548200 242800 548400 243000
rect 548600 242800 548800 243000
rect 549000 242800 549100 243000
rect 545700 242600 549100 242800
rect 545700 242400 546000 242600
rect 546200 242400 546400 242600
rect 546600 242400 546800 242600
rect 547000 242400 547200 242600
rect 547400 242400 547600 242600
rect 547800 242400 548000 242600
rect 548200 242400 548400 242600
rect 548600 242400 548800 242600
rect 549000 242400 549100 242600
rect 545700 242200 549100 242400
rect 545700 242000 546000 242200
rect 546200 242000 546400 242200
rect 546600 242000 546800 242200
rect 547000 242000 547200 242200
rect 547400 242000 547600 242200
rect 547800 242000 548000 242200
rect 548200 242000 548400 242200
rect 548600 242000 548800 242200
rect 549000 242000 549100 242200
rect 545700 241800 549100 242000
rect 545700 241600 546000 241800
rect 546200 241600 546400 241800
rect 546600 241600 546800 241800
rect 547000 241600 547200 241800
rect 547400 241600 547600 241800
rect 547800 241600 548000 241800
rect 548200 241600 548400 241800
rect 548600 241600 548800 241800
rect 549000 241600 549100 241800
rect 545700 241400 549100 241600
rect 545700 241200 546000 241400
rect 546200 241200 546400 241400
rect 546600 241200 546800 241400
rect 547000 241200 547200 241400
rect 547400 241200 547600 241400
rect 547800 241200 548000 241400
rect 548200 241200 548400 241400
rect 548600 241200 548800 241400
rect 549000 241200 549100 241400
rect 545700 241000 549100 241200
rect 545700 240800 546000 241000
rect 546200 240800 546400 241000
rect 546600 240800 546800 241000
rect 547000 240800 547200 241000
rect 547400 240800 547600 241000
rect 547800 240800 548000 241000
rect 548200 240800 548400 241000
rect 548600 240800 548800 241000
rect 549000 240800 549100 241000
rect 545700 240600 549100 240800
rect 545700 240400 546000 240600
rect 546200 240400 546400 240600
rect 546600 240400 546800 240600
rect 547000 240400 547200 240600
rect 547400 240400 547600 240600
rect 547800 240400 548000 240600
rect 548200 240400 548400 240600
rect 548600 240400 548800 240600
rect 549000 240400 549100 240600
rect 545700 240200 549100 240400
rect 545700 240000 546000 240200
rect 546200 240000 546400 240200
rect 546600 240000 546800 240200
rect 547000 240000 547200 240200
rect 547400 240000 547600 240200
rect 547800 240000 548000 240200
rect 548200 240000 548400 240200
rect 548600 240000 548800 240200
rect 549000 240000 549100 240200
rect 545700 239800 549100 240000
rect 545700 239600 546000 239800
rect 546200 239600 546400 239800
rect 546600 239600 546800 239800
rect 547000 239600 547200 239800
rect 547400 239600 547600 239800
rect 547800 239600 548000 239800
rect 548200 239600 548400 239800
rect 548600 239600 548800 239800
rect 549000 239600 549100 239800
rect 545700 239400 549100 239600
rect 545700 239200 546000 239400
rect 546200 239200 546400 239400
rect 546600 239200 546800 239400
rect 547000 239200 547200 239400
rect 547400 239200 547600 239400
rect 547800 239200 548000 239400
rect 548200 239200 548400 239400
rect 548600 239200 548800 239400
rect 549000 239200 549100 239400
rect 545700 239000 549100 239200
rect 545700 238800 546000 239000
rect 546200 238800 546400 239000
rect 546600 238800 546800 239000
rect 547000 238800 547200 239000
rect 547400 238800 547600 239000
rect 547800 238800 548000 239000
rect 548200 238800 548400 239000
rect 548600 238800 548800 239000
rect 549000 238800 549100 239000
rect 545700 238600 549100 238800
rect 545700 238400 546000 238600
rect 546200 238400 546400 238600
rect 546600 238400 546800 238600
rect 547000 238400 547200 238600
rect 547400 238400 547600 238600
rect 547800 238400 548000 238600
rect 548200 238400 548400 238600
rect 548600 238400 548800 238600
rect 549000 238400 549100 238600
rect 545700 238200 549100 238400
rect 545700 238000 546000 238200
rect 546200 238000 546400 238200
rect 546600 238000 546800 238200
rect 547000 238000 547200 238200
rect 547400 238000 547600 238200
rect 547800 238000 548000 238200
rect 548200 238000 548400 238200
rect 548600 238000 548800 238200
rect 549000 238000 549100 238200
rect 545700 237800 549100 238000
rect 545700 237600 546000 237800
rect 546200 237600 546400 237800
rect 546600 237600 546800 237800
rect 547000 237600 547200 237800
rect 547400 237600 547600 237800
rect 547800 237600 548000 237800
rect 548200 237600 548400 237800
rect 548600 237600 548800 237800
rect 549000 237600 549100 237800
rect 545700 237400 549100 237600
rect 545700 237200 546000 237400
rect 546200 237200 546400 237400
rect 546600 237200 546800 237400
rect 547000 237200 547200 237400
rect 547400 237200 547600 237400
rect 547800 237200 548000 237400
rect 548200 237200 548400 237400
rect 548600 237200 548800 237400
rect 549000 237200 549100 237400
rect 545700 237000 549100 237200
rect 545700 236800 546000 237000
rect 546200 236800 546400 237000
rect 546600 236800 546800 237000
rect 547000 236800 547200 237000
rect 547400 236800 547600 237000
rect 547800 236800 548000 237000
rect 548200 236800 548400 237000
rect 548600 236800 548800 237000
rect 549000 236800 549100 237000
rect 545700 236600 549100 236800
rect 545700 236400 546000 236600
rect 546200 236400 546400 236600
rect 546600 236400 546800 236600
rect 547000 236400 547200 236600
rect 547400 236400 547600 236600
rect 547800 236400 548000 236600
rect 548200 236400 548400 236600
rect 548600 236400 548800 236600
rect 549000 236400 549100 236600
rect 545700 236200 549100 236400
rect 545700 236000 546000 236200
rect 546200 236000 546400 236200
rect 546600 236000 546800 236200
rect 547000 236000 547200 236200
rect 547400 236000 547600 236200
rect 547800 236000 548000 236200
rect 548200 236000 548400 236200
rect 548600 236000 548800 236200
rect 549000 236000 549100 236200
rect 545700 235800 549100 236000
rect 545700 235600 546000 235800
rect 546200 235600 546400 235800
rect 546600 235600 546800 235800
rect 547000 235600 547200 235800
rect 547400 235600 547600 235800
rect 547800 235600 548000 235800
rect 548200 235600 548400 235800
rect 548600 235600 548800 235800
rect 549000 235600 549100 235800
rect 545700 235400 549100 235600
rect 545700 235200 546000 235400
rect 546200 235200 546400 235400
rect 546600 235200 546800 235400
rect 547000 235200 547200 235400
rect 547400 235200 547600 235400
rect 547800 235200 548000 235400
rect 548200 235200 548400 235400
rect 548600 235200 548800 235400
rect 549000 235200 549100 235400
rect 545700 235000 549100 235200
rect 545700 234800 546000 235000
rect 546200 234800 546400 235000
rect 546600 234800 546800 235000
rect 547000 234800 547200 235000
rect 547400 234800 547600 235000
rect 547800 234800 548000 235000
rect 548200 234800 548400 235000
rect 548600 234800 548800 235000
rect 549000 234800 549100 235000
rect 545700 234700 549100 234800
rect 545700 234500 546000 234700
rect 546200 234500 546400 234700
rect 546600 234500 546800 234700
rect 547000 234500 547200 234700
rect 547400 234500 547600 234700
rect 547800 234500 548000 234700
rect 548200 234500 548400 234700
rect 548600 234500 548800 234700
rect 549000 234500 549100 234700
rect 545700 234400 549100 234500
rect 545700 234200 546000 234400
rect 546200 234200 546400 234400
rect 546600 234200 546800 234400
rect 547000 234200 547200 234400
rect 547400 234200 547600 234400
rect 547800 234200 548000 234400
rect 548200 234200 548400 234400
rect 548600 234200 548800 234400
rect 549000 234200 549100 234400
rect 545700 234000 549100 234200
rect 545700 233800 546000 234000
rect 546200 233800 546400 234000
rect 546600 233800 546800 234000
rect 547000 233800 547200 234000
rect 547400 233800 547600 234000
rect 547800 233800 548000 234000
rect 548200 233800 548400 234000
rect 548600 233800 548800 234000
rect 549000 233800 549100 234000
rect 545700 233700 549100 233800
rect 511500 195200 512000 195600
rect 512400 195200 512800 195600
rect 513200 195200 513600 195600
rect 514000 195200 514400 195600
rect 514800 195200 515200 195600
rect 515600 195200 516000 195600
rect 516400 195200 517000 195600
rect 511500 194800 517000 195200
rect 511500 194400 512000 194800
rect 512400 194400 512800 194800
rect 513200 194400 513600 194800
rect 514000 194400 514400 194800
rect 514800 194400 515200 194800
rect 515600 194400 516000 194800
rect 516400 194400 517000 194800
rect 511500 194000 517000 194400
rect 511500 193600 512000 194000
rect 512400 193600 512800 194000
rect 513200 193600 513600 194000
rect 514000 193600 514400 194000
rect 514800 193600 515200 194000
rect 515600 193600 516000 194000
rect 516400 193600 517000 194000
rect 511500 193200 517000 193600
rect 511500 192800 512000 193200
rect 512400 192800 512800 193200
rect 513200 192800 513600 193200
rect 514000 192800 514400 193200
rect 514800 192800 515200 193200
rect 515600 192800 516000 193200
rect 516400 192800 517000 193200
rect 511500 192400 517000 192800
rect 511500 192000 512000 192400
rect 512400 192000 512800 192400
rect 513200 192000 513600 192400
rect 514000 192000 514400 192400
rect 514800 192000 515200 192400
rect 515600 192000 516000 192400
rect 516400 192000 517000 192400
rect 511500 191600 517000 192000
rect 511500 191200 512000 191600
rect 512400 191200 512800 191600
rect 513200 191200 513600 191600
rect 514000 191200 514400 191600
rect 514800 191200 515200 191600
rect 515600 191200 516000 191600
rect 516400 191200 517000 191600
rect 511500 190800 517000 191200
rect 511500 190400 512000 190800
rect 512400 190400 512800 190800
rect 513200 190400 513600 190800
rect 514000 190400 514400 190800
rect 514800 190400 515200 190800
rect 515600 190400 516000 190800
rect 516400 190400 517000 190800
rect 511500 190000 517000 190400
rect 511500 189600 512000 190000
rect 512400 189600 512800 190000
rect 513200 189600 513600 190000
rect 514000 189600 514400 190000
rect 514800 189600 515200 190000
rect 515600 189600 516000 190000
rect 516400 189600 517000 190000
rect 511500 189200 517000 189600
rect 511500 188800 512000 189200
rect 512400 188800 512800 189200
rect 513200 188800 513600 189200
rect 514000 188800 514400 189200
rect 514800 188800 515200 189200
rect 515600 188800 516000 189200
rect 516400 188800 517000 189200
rect 511500 188400 517000 188800
rect 511500 188000 512000 188400
rect 512400 188000 512800 188400
rect 513200 188000 513600 188400
rect 514000 188000 514400 188400
rect 514800 188000 515200 188400
rect 515600 188000 516000 188400
rect 516400 188000 517000 188400
rect 511500 187600 517000 188000
rect 511500 187200 512000 187600
rect 512400 187200 512800 187600
rect 513200 187200 513600 187600
rect 514000 187200 514400 187600
rect 514800 187200 515200 187600
rect 515600 187200 516000 187600
rect 516400 187200 517000 187600
rect 511500 186800 517000 187200
rect 511500 186400 512000 186800
rect 512400 186400 512800 186800
rect 513200 186400 513600 186800
rect 514000 186400 514400 186800
rect 514800 186400 515200 186800
rect 515600 186400 516000 186800
rect 516400 186400 517000 186800
rect 511500 186000 517000 186400
rect 511500 185600 512000 186000
rect 512400 185600 512800 186000
rect 513200 185600 513600 186000
rect 514000 185600 514400 186000
rect 514800 185600 515200 186000
rect 515600 185600 516000 186000
rect 516400 185600 517000 186000
rect 511500 185200 517000 185600
rect 511500 184800 512000 185200
rect 512400 184800 512800 185200
rect 513200 184800 513600 185200
rect 514000 184800 514400 185200
rect 514800 184800 515200 185200
rect 515600 184800 516000 185200
rect 516400 184800 517000 185200
rect 511500 184400 517000 184800
rect 511500 184000 512000 184400
rect 512400 184000 512800 184400
rect 513200 184000 513600 184400
rect 514000 184000 514400 184400
rect 514800 184000 515200 184400
rect 515600 184000 516000 184400
rect 516400 184000 517000 184400
rect 511500 183600 517000 184000
rect 511500 183200 512000 183600
rect 512400 183200 512800 183600
rect 513200 183200 513600 183600
rect 514000 183200 514400 183600
rect 514800 183200 515200 183600
rect 515600 183200 516000 183600
rect 516400 183200 517000 183600
rect 511500 182800 517000 183200
rect 511500 182400 512000 182800
rect 512400 182400 512800 182800
rect 513200 182400 513600 182800
rect 514000 182400 514400 182800
rect 514800 182400 515200 182800
rect 515600 182400 516000 182800
rect 516400 182400 517000 182800
rect 511500 182000 517000 182400
rect 511500 181600 512000 182000
rect 512400 181600 512800 182000
rect 513200 181600 513600 182000
rect 514000 181600 514400 182000
rect 514800 181600 515200 182000
rect 515600 181600 516000 182000
rect 516400 181600 517000 182000
rect 511500 181150 517000 181600
rect 297000 177200 299400 177600
rect 299800 177200 300200 177600
rect 300600 177200 301000 177600
rect 301400 177200 301800 177600
rect 302200 177200 302600 177600
rect 303000 177200 303400 177600
rect 303800 177200 306000 177600
rect 297000 176800 306000 177200
rect 297000 176400 299400 176800
rect 299800 176400 300200 176800
rect 300600 176400 301000 176800
rect 301400 176400 301800 176800
rect 302200 176400 302600 176800
rect 303000 176400 303400 176800
rect 303800 176400 306000 176800
rect 297000 176000 306000 176400
rect 297000 175600 299400 176000
rect 299800 175600 300200 176000
rect 300600 175600 301000 176000
rect 301400 175600 301800 176000
rect 302200 175600 302600 176000
rect 303000 175600 303400 176000
rect 303800 175600 306000 176000
rect 297000 175200 306000 175600
rect 297000 174800 299400 175200
rect 299800 174800 300200 175200
rect 300600 174800 301000 175200
rect 301400 174800 301800 175200
rect 302200 174800 302600 175200
rect 303000 174800 303400 175200
rect 303800 174800 306000 175200
rect 297000 174400 306000 174800
rect 297000 174000 299400 174400
rect 299800 174000 300200 174400
rect 300600 174000 301000 174400
rect 301400 174000 301800 174400
rect 302200 174000 302600 174400
rect 303000 174000 303400 174400
rect 303800 174000 306000 174400
rect 297000 173600 306000 174000
rect 297000 173200 299400 173600
rect 299800 173200 300200 173600
rect 300600 173200 301000 173600
rect 301400 173200 301800 173600
rect 302200 173200 302600 173600
rect 303000 173200 303400 173600
rect 303800 173200 306000 173600
rect 297000 172800 306000 173200
rect 297000 172400 299400 172800
rect 299800 172400 300200 172800
rect 300600 172400 301000 172800
rect 301400 172400 301800 172800
rect 302200 172400 302600 172800
rect 303000 172400 303400 172800
rect 303800 172400 306000 172800
rect 297000 172000 306000 172400
rect 297000 171600 299400 172000
rect 299800 171600 300200 172000
rect 300600 171600 301000 172000
rect 301400 171600 301800 172000
rect 302200 171600 302600 172000
rect 303000 171600 303400 172000
rect 303800 171600 306000 172000
rect 297000 171200 306000 171600
rect 297000 170800 299400 171200
rect 299800 170800 300200 171200
rect 300600 170800 301000 171200
rect 301400 170800 301800 171200
rect 302200 170800 302600 171200
rect 303000 170800 303400 171200
rect 303800 170800 306000 171200
rect 297000 170400 306000 170800
rect 297000 170000 299400 170400
rect 299800 170000 300200 170400
rect 300600 170000 301000 170400
rect 301400 170000 301800 170400
rect 302200 170000 302600 170400
rect 303000 170000 303400 170400
rect 303800 170000 306000 170400
rect 297000 169600 306000 170000
rect 297000 169200 299400 169600
rect 299800 169200 300200 169600
rect 300600 169200 301000 169600
rect 301400 169200 301800 169600
rect 302200 169200 302600 169600
rect 303000 169200 303400 169600
rect 303800 169200 306000 169600
rect 297000 168800 306000 169200
rect 297000 168400 299400 168800
rect 299800 168400 300200 168800
rect 300600 168400 301000 168800
rect 301400 168400 301800 168800
rect 302200 168400 302600 168800
rect 303000 168400 303400 168800
rect 303800 168400 306000 168800
rect 297000 168000 306000 168400
rect 297000 167600 299400 168000
rect 299800 167600 300200 168000
rect 300600 167600 301000 168000
rect 301400 167600 301800 168000
rect 302200 167600 302600 168000
rect 303000 167600 303400 168000
rect 303800 167600 306000 168000
rect 297000 167200 306000 167600
rect 297000 166800 299400 167200
rect 299800 166800 300200 167200
rect 300600 166800 301000 167200
rect 301400 166800 301800 167200
rect 302200 166800 302600 167200
rect 303000 166800 303400 167200
rect 303800 166800 306000 167200
rect 297000 166400 306000 166800
rect 297000 166000 299400 166400
rect 299800 166000 300200 166400
rect 300600 166000 301000 166400
rect 301400 166000 301800 166400
rect 302200 166000 302600 166400
rect 303000 166000 303400 166400
rect 303800 166000 306000 166400
rect 297000 165600 306000 166000
rect 297000 165200 299400 165600
rect 299800 165200 300200 165600
rect 300600 165200 301000 165600
rect 301400 165200 301800 165600
rect 302200 165200 302600 165600
rect 303000 165200 303400 165600
rect 303800 165200 306000 165600
rect 297000 164800 306000 165200
rect 297000 164400 299400 164800
rect 299800 164400 300200 164800
rect 300600 164400 301000 164800
rect 301400 164400 301800 164800
rect 302200 164400 302600 164800
rect 303000 164400 303400 164800
rect 303800 164400 306000 164800
rect 297000 164000 306000 164400
rect 297000 163600 299400 164000
rect 299800 163600 300200 164000
rect 300600 163600 301000 164000
rect 301400 163600 301800 164000
rect 302200 163600 302600 164000
rect 303000 163600 303400 164000
rect 303800 163600 306000 164000
rect 297000 162900 306000 163600
<< rmetal4 >>
rect 515500 697940 521000 698500
<< via4 >>
rect 12900 673800 13200 674100
rect 13700 673800 14000 674100
rect 12900 673300 13200 673600
rect 13700 673300 14000 673600
rect 12900 672800 13200 673100
rect 13700 672800 14000 673100
rect 2500 648300 2800 648600
rect 3000 648300 3300 648600
rect 3500 648300 3800 648600
rect 23400 648200 23700 648500
rect 24100 648200 24400 648500
rect 2500 647800 2800 648100
rect 3000 647800 3300 648100
rect 3500 647800 3800 648100
rect 2500 647300 2800 647600
rect 3000 647300 3300 647600
rect 3500 647300 3800 647600
rect 23400 647600 23700 647900
rect 24100 647600 24400 647900
rect 2500 646800 2800 647100
rect 3000 646800 3300 647100
rect 3500 646800 3800 647100
rect 23400 647000 23700 647300
rect 24100 647000 24400 647300
rect 2500 646300 2800 646600
rect 3000 646300 3300 646600
rect 3500 646300 3800 646600
rect 23400 646300 23700 646600
rect 24100 646300 24400 646600
rect 2500 645800 2800 646100
rect 3000 645800 3300 646100
rect 3500 645800 3800 646100
rect 23400 645700 23700 646000
rect 24100 645700 24400 646000
rect 2500 645300 2800 645600
rect 3000 645300 3300 645600
rect 3500 645300 3800 645600
rect 2500 644800 2800 645100
rect 3000 644800 3300 645100
rect 3500 644800 3800 645100
rect 23400 645100 23700 645400
rect 24100 645100 24400 645400
rect 2500 644300 2800 644600
rect 3000 644300 3300 644600
rect 3500 644300 3800 644600
rect 23400 644500 23700 644800
rect 24100 644500 24400 644800
rect 2500 643800 2800 644100
rect 3000 643800 3300 644100
rect 3500 643800 3800 644100
rect 23400 643900 23700 644200
rect 24100 643900 24400 644200
rect 2500 643300 2800 643600
rect 3000 643300 3300 643600
rect 3500 643300 3800 643600
rect 23400 643300 23700 643600
rect 24100 643300 24400 643600
rect 2500 642800 2800 643100
rect 3000 642800 3300 643100
rect 3500 642800 3800 643100
rect 2500 642300 2800 642600
rect 3000 642300 3300 642600
rect 3500 642300 3800 642600
rect 23400 642600 23700 642900
rect 24100 642600 24400 642900
rect 2500 641800 2800 642100
rect 3000 641800 3300 642100
rect 3500 641800 3800 642100
rect 23400 642000 23700 642300
rect 24100 642000 24400 642300
rect 2500 641300 2800 641600
rect 3000 641300 3300 641600
rect 3500 641300 3800 641600
rect 23400 641400 23700 641700
rect 24100 641400 24400 641700
rect 2500 640800 2800 641100
rect 3000 640800 3300 641100
rect 3500 640800 3800 641100
rect 23400 640800 23700 641100
rect 24100 640800 24400 641100
rect 2500 640300 2800 640600
rect 3000 640300 3300 640600
rect 3500 640300 3800 640600
rect 23400 640200 23700 640500
rect 24100 640200 24400 640500
rect 2500 639800 2800 640100
rect 3000 639800 3300 640100
rect 3500 639800 3800 640100
rect 2500 639300 2800 639600
rect 3000 639300 3300 639600
rect 3500 639300 3800 639600
rect 23400 639600 23700 639900
rect 24100 639600 24400 639900
rect 2500 638800 2800 639100
rect 3000 638800 3300 639100
rect 3500 638800 3800 639100
rect 23400 639000 23700 639300
rect 24100 639000 24400 639300
rect 2500 638300 2800 638600
rect 3000 638300 3300 638600
rect 3500 638300 3800 638600
rect 23400 638400 23700 638700
rect 24100 638400 24400 638700
rect 2500 637800 2800 638100
rect 3000 637800 3300 638100
rect 3500 637800 3800 638100
rect 23400 637800 23700 638100
rect 24100 637800 24400 638100
rect 2500 637300 2800 637600
rect 3000 637300 3300 637600
rect 3500 637300 3800 637600
rect 2500 636800 2800 637100
rect 3000 636800 3300 637100
rect 3500 636800 3800 637100
rect 23400 637100 23700 637400
rect 24100 637100 24400 637400
rect 2500 636300 2800 636600
rect 3000 636300 3300 636600
rect 3500 636300 3800 636600
rect 23400 636400 23700 636700
rect 24100 636400 24400 636700
rect 2500 635800 2800 636100
rect 3000 635800 3300 636100
rect 3500 635800 3800 636100
rect 23400 635700 23700 636000
rect 24100 635700 24400 636000
rect 2500 635300 2800 635600
rect 3000 635300 3300 635600
rect 3500 635300 3800 635600
rect 2500 634800 2800 635100
rect 3000 634800 3300 635100
rect 3500 634800 3800 635100
rect 23400 634900 23700 635200
rect 24100 634900 24400 635200
rect 2500 634300 2800 634600
rect 3000 634300 3300 634600
rect 3500 634300 3800 634600
rect 23400 634200 23700 634500
rect 24100 634200 24400 634500
rect 32800 673700 33100 674000
rect 33300 673700 33600 674000
rect 33800 673700 34100 674000
rect 34300 673700 34600 674000
rect 34800 673700 35100 674000
rect 35300 673700 35600 674000
rect 35800 673700 36100 674000
rect 36300 673700 36600 674000
rect 36800 673700 37100 674000
rect 37300 673700 37600 674000
rect 37800 673700 38100 674000
rect 38300 673700 38600 674000
rect 38800 673700 39100 674000
rect 39300 673700 39600 674000
rect 39800 673700 40100 674000
rect 40300 673700 40600 674000
rect 32800 672900 33100 673200
rect 33300 672900 33600 673200
rect 33800 672900 34100 673200
rect 34300 672900 34600 673200
rect 34800 672900 35100 673200
rect 35300 672900 35600 673200
rect 35800 672900 36100 673200
rect 36300 672900 36600 673200
rect 36800 672900 37100 673200
rect 37300 672900 37600 673200
rect 37800 672900 38100 673200
rect 38300 672900 38600 673200
rect 38800 672900 39100 673200
rect 39300 672900 39600 673200
rect 39800 672900 40100 673200
rect 40300 672900 40600 673200
rect 50100 673700 50400 674000
rect 50100 673300 50400 673600
rect 50100 672900 50400 673200
rect 32800 670400 33100 670700
rect 33300 670400 33600 670700
rect 33800 670400 34100 670700
rect 34300 670400 34600 670700
rect 34800 670400 35100 670700
rect 35300 670400 35600 670700
rect 35800 670400 36100 670700
rect 36300 670400 36600 670700
rect 36800 670400 37100 670700
rect 37300 670400 37600 670700
rect 37800 670400 38100 670700
rect 38300 670400 38600 670700
rect 38800 670400 39100 670700
rect 39300 670400 39600 670700
rect 39800 670400 40100 670700
rect 40300 670400 40600 670700
rect 32800 669700 33100 670000
rect 33300 669700 33600 670000
rect 33800 669700 34100 670000
rect 34300 669700 34600 670000
rect 34800 669700 35100 670000
rect 35300 669700 35600 670000
rect 35800 669700 36100 670000
rect 36300 669700 36600 670000
rect 36800 669700 37100 670000
rect 37300 669700 37600 670000
rect 37800 669700 38100 670000
rect 38300 669700 38600 670000
rect 38800 669700 39100 670000
rect 39300 669700 39600 670000
rect 39800 669700 40100 670000
rect 40300 669700 40600 670000
rect 32800 667100 33100 667400
rect 33300 667100 33600 667400
rect 33800 667100 34100 667400
rect 34300 667100 34600 667400
rect 34800 667100 35100 667400
rect 35300 667100 35600 667400
rect 35800 667100 36100 667400
rect 36300 667100 36600 667400
rect 36800 667100 37100 667400
rect 37300 667100 37600 667400
rect 37800 667100 38100 667400
rect 38300 667100 38600 667400
rect 38800 667100 39100 667400
rect 39300 667100 39600 667400
rect 39800 667100 40100 667400
rect 40300 667100 40600 667400
rect 32800 666400 33100 666700
rect 33300 666400 33600 666700
rect 33800 666400 34100 666700
rect 34300 666400 34600 666700
rect 34800 666400 35100 666700
rect 35300 666400 35600 666700
rect 35800 666400 36100 666700
rect 36300 666400 36600 666700
rect 36800 666400 37100 666700
rect 37300 666400 37600 666700
rect 37800 666400 38100 666700
rect 38300 666400 38600 666700
rect 38800 666400 39100 666700
rect 39300 666400 39600 666700
rect 39800 666400 40100 666700
rect 40300 666400 40600 666700
rect 549900 684600 550200 684900
rect 550400 684600 550700 684900
rect 550900 684600 551200 684900
rect 551400 684600 551700 684900
rect 551900 684600 552200 684900
rect 552400 684600 552700 684900
rect 549900 684100 550200 684400
rect 550400 684100 550700 684400
rect 550900 684100 551200 684400
rect 551400 684100 551700 684400
rect 551900 684100 552200 684400
rect 552400 684100 552700 684400
rect 549900 683600 550200 683900
rect 550400 683600 550700 683900
rect 550900 683600 551200 683900
rect 551400 683600 551700 683900
rect 551900 683600 552200 683900
rect 552400 683600 552700 683900
rect 573200 684600 573500 684900
rect 573800 684600 574100 684900
rect 573200 684100 573500 684400
rect 573800 684100 574100 684400
rect 576800 684400 577100 684700
rect 577300 684400 577600 684700
rect 577800 684400 578100 684700
rect 578300 684400 578600 684700
rect 573200 683600 573500 683900
rect 573800 683600 574100 683900
rect 576800 683900 577100 684200
rect 577300 683900 577600 684200
rect 577800 683900 578100 684200
rect 578300 683900 578600 684200
rect 58000 648300 58300 648600
rect 58500 648300 58800 648600
rect 59000 648300 59300 648600
rect 59500 648300 59800 648600
rect 60000 648300 60300 648600
rect 60500 648300 60800 648600
rect 61000 648300 61300 648600
rect 61500 648300 61800 648600
rect 58000 647800 58300 648100
rect 58500 647800 58800 648100
rect 59000 647800 59300 648100
rect 59500 647800 59800 648100
rect 60000 647800 60300 648100
rect 60500 647800 60800 648100
rect 61000 647800 61300 648100
rect 61500 647800 61800 648100
rect 58000 647300 58300 647600
rect 58500 647300 58800 647600
rect 59000 647300 59300 647600
rect 59500 647300 59800 647600
rect 60000 647300 60300 647600
rect 60500 647300 60800 647600
rect 61000 647300 61300 647600
rect 61500 647300 61800 647600
rect 58000 646800 58300 647100
rect 58500 646800 58800 647100
rect 59000 646800 59300 647100
rect 59500 646800 59800 647100
rect 60000 646800 60300 647100
rect 60500 646800 60800 647100
rect 61000 646800 61300 647100
rect 61500 646800 61800 647100
rect 58000 646300 58300 646600
rect 58500 646300 58800 646600
rect 59000 646300 59300 646600
rect 59500 646300 59800 646600
rect 60000 646300 60300 646600
rect 60500 646300 60800 646600
rect 61000 646300 61300 646600
rect 61500 646300 61800 646600
rect 58000 645800 58300 646100
rect 58500 645800 58800 646100
rect 59000 645800 59300 646100
rect 59500 645800 59800 646100
rect 60000 645800 60300 646100
rect 60500 645800 60800 646100
rect 61000 645800 61300 646100
rect 61500 645800 61800 646100
rect 58000 645300 58300 645600
rect 58500 645300 58800 645600
rect 59000 645300 59300 645600
rect 59500 645300 59800 645600
rect 60000 645300 60300 645600
rect 60500 645300 60800 645600
rect 61000 645300 61300 645600
rect 61500 645300 61800 645600
rect 58000 644800 58300 645100
rect 58500 644800 58800 645100
rect 59000 644800 59300 645100
rect 59500 644800 59800 645100
rect 60000 644800 60300 645100
rect 60500 644800 60800 645100
rect 61000 644800 61300 645100
rect 61500 644800 61800 645100
rect 58000 644300 58300 644600
rect 58500 644300 58800 644600
rect 59000 644300 59300 644600
rect 59500 644300 59800 644600
rect 60000 644300 60300 644600
rect 60500 644300 60800 644600
rect 61000 644300 61300 644600
rect 61500 644300 61800 644600
rect 58000 643800 58300 644100
rect 58500 643800 58800 644100
rect 59000 643800 59300 644100
rect 59500 643800 59800 644100
rect 60000 643800 60300 644100
rect 60500 643800 60800 644100
rect 61000 643800 61300 644100
rect 61500 643800 61800 644100
rect 58000 643300 58300 643600
rect 58500 643300 58800 643600
rect 59000 643300 59300 643600
rect 59500 643300 59800 643600
rect 60000 643300 60300 643600
rect 60500 643300 60800 643600
rect 61000 643300 61300 643600
rect 61500 643300 61800 643600
rect 58000 642800 58300 643100
rect 58500 642800 58800 643100
rect 59000 642800 59300 643100
rect 59500 642800 59800 643100
rect 60000 642800 60300 643100
rect 60500 642800 60800 643100
rect 61000 642800 61300 643100
rect 61500 642800 61800 643100
rect 58000 642300 58300 642600
rect 58500 642300 58800 642600
rect 59000 642300 59300 642600
rect 59500 642300 59800 642600
rect 60000 642300 60300 642600
rect 60500 642300 60800 642600
rect 61000 642300 61300 642600
rect 61500 642300 61800 642600
rect 58000 641800 58300 642100
rect 58500 641800 58800 642100
rect 59000 641800 59300 642100
rect 59500 641800 59800 642100
rect 60000 641800 60300 642100
rect 60500 641800 60800 642100
rect 61000 641800 61300 642100
rect 61500 641800 61800 642100
rect 58000 641300 58300 641600
rect 58500 641300 58800 641600
rect 59000 641300 59300 641600
rect 59500 641300 59800 641600
rect 60000 641300 60300 641600
rect 60500 641300 60800 641600
rect 61000 641300 61300 641600
rect 61500 641300 61800 641600
rect 58000 640800 58300 641100
rect 58500 640800 58800 641100
rect 59000 640800 59300 641100
rect 59500 640800 59800 641100
rect 60000 640800 60300 641100
rect 60500 640800 60800 641100
rect 61000 640800 61300 641100
rect 61500 640800 61800 641100
rect 58000 640300 58300 640600
rect 58500 640300 58800 640600
rect 59000 640300 59300 640600
rect 59500 640300 59800 640600
rect 60000 640300 60300 640600
rect 60500 640300 60800 640600
rect 61000 640300 61300 640600
rect 61500 640300 61800 640600
rect 58000 639800 58300 640100
rect 58500 639800 58800 640100
rect 59000 639800 59300 640100
rect 59500 639800 59800 640100
rect 60000 639800 60300 640100
rect 60500 639800 60800 640100
rect 61000 639800 61300 640100
rect 61500 639800 61800 640100
rect 58000 639300 58300 639600
rect 58500 639300 58800 639600
rect 59000 639300 59300 639600
rect 59500 639300 59800 639600
rect 60000 639300 60300 639600
rect 60500 639300 60800 639600
rect 61000 639300 61300 639600
rect 61500 639300 61800 639600
rect 58000 638800 58300 639100
rect 58500 638800 58800 639100
rect 59000 638800 59300 639100
rect 59500 638800 59800 639100
rect 60000 638800 60300 639100
rect 60500 638800 60800 639100
rect 61000 638800 61300 639100
rect 61500 638800 61800 639100
rect 58000 638300 58300 638600
rect 58500 638300 58800 638600
rect 59000 638300 59300 638600
rect 59500 638300 59800 638600
rect 60000 638300 60300 638600
rect 60500 638300 60800 638600
rect 61000 638300 61300 638600
rect 61500 638300 61800 638600
rect 58000 637800 58300 638100
rect 58500 637800 58800 638100
rect 59000 637800 59300 638100
rect 59500 637800 59800 638100
rect 60000 637800 60300 638100
rect 60500 637800 60800 638100
rect 61000 637800 61300 638100
rect 61500 637800 61800 638100
rect 58000 637300 58300 637600
rect 58500 637300 58800 637600
rect 59000 637300 59300 637600
rect 59500 637300 59800 637600
rect 60000 637300 60300 637600
rect 60500 637300 60800 637600
rect 61000 637300 61300 637600
rect 61500 637300 61800 637600
rect 58000 636800 58300 637100
rect 58500 636800 58800 637100
rect 59000 636800 59300 637100
rect 59500 636800 59800 637100
rect 60000 636800 60300 637100
rect 60500 636800 60800 637100
rect 61000 636800 61300 637100
rect 61500 636800 61800 637100
rect 58000 636300 58300 636600
rect 58500 636300 58800 636600
rect 59000 636300 59300 636600
rect 59500 636300 59800 636600
rect 60000 636300 60300 636600
rect 60500 636300 60800 636600
rect 61000 636300 61300 636600
rect 61500 636300 61800 636600
rect 58000 635800 58300 636100
rect 58500 635800 58800 636100
rect 59000 635800 59300 636100
rect 59500 635800 59800 636100
rect 60000 635800 60300 636100
rect 60500 635800 60800 636100
rect 61000 635800 61300 636100
rect 61500 635800 61800 636100
rect 58000 635300 58300 635600
rect 58500 635300 58800 635600
rect 59000 635300 59300 635600
rect 59500 635300 59800 635600
rect 60000 635300 60300 635600
rect 60500 635300 60800 635600
rect 61000 635300 61300 635600
rect 61500 635300 61800 635600
rect 58000 634800 58300 635100
rect 58500 634800 58800 635100
rect 59000 634800 59300 635100
rect 59500 634800 59800 635100
rect 60000 634800 60300 635100
rect 60500 634800 60800 635100
rect 61000 634800 61300 635100
rect 61500 634800 61800 635100
rect 58000 634300 58300 634600
rect 58500 634300 58800 634600
rect 59000 634300 59300 634600
rect 59500 634300 59800 634600
rect 60000 634300 60300 634600
rect 60500 634300 60800 634600
rect 61000 634300 61300 634600
rect 61500 634300 61800 634600
rect 289600 344100 289900 344400
rect 294800 343900 295100 344200
rect 289600 343600 289900 343900
rect 299000 343900 299400 344300
rect 299600 343900 300000 344300
rect 300200 343900 300600 344300
rect 300800 343900 301200 344300
rect 301400 343900 301800 344300
rect 302000 343900 302400 344300
rect 302600 343900 303000 344300
rect 303200 343900 303600 344300
rect 289600 343100 289900 343400
rect 299000 343300 299400 343700
rect 299600 343300 300000 343700
rect 300200 343300 300600 343700
rect 300800 343300 301200 343700
rect 301400 343300 301800 343700
rect 302000 343300 302400 343700
rect 302600 343300 303000 343700
rect 303200 343300 303600 343700
rect 287500 342000 287800 342300
rect 288000 342000 288300 342300
rect 288300 340500 288600 340800
rect 59400 289500 59700 289800
rect 59900 289500 60200 289800
rect 60400 289500 60700 289800
rect 60900 289500 61200 289800
rect 61400 289500 61700 289800
rect 61900 289500 62200 289800
rect 62400 289500 62700 289800
rect 62900 289500 63200 289800
rect 63400 289500 63700 289800
rect 63900 289500 64200 289800
rect 64400 289500 64700 289800
rect 64900 289500 65200 289800
rect 65400 289500 65700 289800
rect 65900 289500 66200 289800
rect 66400 289500 66700 289800
rect 66900 289500 67200 289800
rect 67400 289500 67700 289800
rect 67900 289500 68200 289800
rect 68400 289500 68700 289800
rect 68900 289500 69200 289800
rect 69400 289500 69700 289800
rect 69900 289500 70200 289800
rect 70400 289500 70700 289800
rect 70900 289500 71200 289800
rect 71400 289500 71700 289800
rect 71900 289500 72200 289800
rect 72400 289500 72700 289800
rect 72900 289500 73200 289800
rect 73400 289500 73700 289800
rect 59400 289000 59700 289300
rect 59900 289000 60200 289300
rect 60400 289000 60700 289300
rect 60900 289000 61200 289300
rect 61400 289000 61700 289300
rect 61900 289000 62200 289300
rect 62400 289000 62700 289300
rect 62900 289000 63200 289300
rect 63400 289000 63700 289300
rect 63900 289000 64200 289300
rect 64400 289000 64700 289300
rect 64900 289000 65200 289300
rect 65400 289000 65700 289300
rect 65900 289000 66200 289300
rect 66400 289000 66700 289300
rect 66900 289000 67200 289300
rect 67400 289000 67700 289300
rect 67900 289000 68200 289300
rect 68400 289000 68700 289300
rect 68900 289000 69200 289300
rect 69400 289000 69700 289300
rect 69900 289000 70200 289300
rect 70400 289000 70700 289300
rect 70900 289000 71200 289300
rect 71400 289000 71700 289300
rect 71900 289000 72200 289300
rect 72400 289000 72700 289300
rect 72900 289000 73200 289300
rect 73400 289000 73700 289300
rect 59400 288500 59700 288800
rect 59900 288500 60200 288800
rect 60400 288500 60700 288800
rect 60900 288500 61200 288800
rect 61400 288500 61700 288800
rect 61900 288500 62200 288800
rect 62400 288500 62700 288800
rect 62900 288500 63200 288800
rect 63400 288500 63700 288800
rect 63900 288500 64200 288800
rect 64400 288500 64700 288800
rect 64900 288500 65200 288800
rect 65400 288500 65700 288800
rect 65900 288500 66200 288800
rect 66400 288500 66700 288800
rect 66900 288500 67200 288800
rect 67400 288500 67700 288800
rect 67900 288500 68200 288800
rect 68400 288500 68700 288800
rect 68900 288500 69200 288800
rect 69400 288500 69700 288800
rect 69900 288500 70200 288800
rect 70400 288500 70700 288800
rect 70900 288500 71200 288800
rect 71400 288500 71700 288800
rect 71900 288500 72200 288800
rect 72400 288500 72700 288800
rect 72900 288500 73200 288800
rect 73400 288500 73700 288800
rect 59400 288000 59700 288300
rect 59900 288000 60200 288300
rect 60400 288000 60700 288300
rect 60900 288000 61200 288300
rect 61400 288000 61700 288300
rect 61900 288000 62200 288300
rect 62400 288000 62700 288300
rect 62900 288000 63200 288300
rect 63400 288000 63700 288300
rect 63900 288000 64200 288300
rect 64400 288000 64700 288300
rect 64900 288000 65200 288300
rect 65400 288000 65700 288300
rect 65900 288000 66200 288300
rect 66400 288000 66700 288300
rect 66900 288000 67200 288300
rect 67400 288000 67700 288300
rect 67900 288000 68200 288300
rect 68400 288000 68700 288300
rect 68900 288000 69200 288300
rect 69400 288000 69700 288300
rect 69900 288000 70200 288300
rect 70400 288000 70700 288300
rect 70900 288000 71200 288300
rect 71400 288000 71700 288300
rect 71900 288000 72200 288300
rect 72400 288000 72700 288300
rect 72900 288000 73200 288300
rect 73400 288000 73700 288300
rect 59400 287500 59700 287800
rect 59900 287500 60200 287800
rect 60400 287500 60700 287800
rect 60900 287500 61200 287800
rect 61400 287500 61700 287800
rect 61900 287500 62200 287800
rect 62400 287500 62700 287800
rect 62900 287500 63200 287800
rect 63400 287500 63700 287800
rect 63900 287500 64200 287800
rect 64400 287500 64700 287800
rect 64900 287500 65200 287800
rect 65400 287500 65700 287800
rect 65900 287500 66200 287800
rect 66400 287500 66700 287800
rect 66900 287500 67200 287800
rect 67400 287500 67700 287800
rect 67900 287500 68200 287800
rect 68400 287500 68700 287800
rect 68900 287500 69200 287800
rect 69400 287500 69700 287800
rect 69900 287500 70200 287800
rect 70400 287500 70700 287800
rect 70900 287500 71200 287800
rect 71400 287500 71700 287800
rect 71900 287500 72200 287800
rect 72400 287500 72700 287800
rect 72900 287500 73200 287800
rect 73400 287500 73700 287800
rect 59400 287000 59700 287300
rect 59900 287000 60200 287300
rect 60400 287000 60700 287300
rect 60900 287000 61200 287300
rect 61400 287000 61700 287300
rect 61900 287000 62200 287300
rect 62400 287000 62700 287300
rect 62900 287000 63200 287300
rect 63400 287000 63700 287300
rect 63900 287000 64200 287300
rect 64400 287000 64700 287300
rect 64900 287000 65200 287300
rect 65400 287000 65700 287300
rect 65900 287000 66200 287300
rect 66400 287000 66700 287300
rect 66900 287000 67200 287300
rect 67400 287000 67700 287300
rect 67900 287000 68200 287300
rect 68400 287000 68700 287300
rect 68900 287000 69200 287300
rect 69400 287000 69700 287300
rect 69900 287000 70200 287300
rect 70400 287000 70700 287300
rect 70900 287000 71200 287300
rect 71400 287000 71700 287300
rect 71900 287000 72200 287300
rect 72400 287000 72700 287300
rect 72900 287000 73200 287300
rect 73400 287000 73700 287300
rect 59400 286500 59700 286800
rect 59900 286500 60200 286800
rect 60400 286500 60700 286800
rect 60900 286500 61200 286800
rect 61400 286500 61700 286800
rect 61900 286500 62200 286800
rect 62400 286500 62700 286800
rect 62900 286500 63200 286800
rect 63400 286500 63700 286800
rect 63900 286500 64200 286800
rect 64400 286500 64700 286800
rect 64900 286500 65200 286800
rect 65400 286500 65700 286800
rect 65900 286500 66200 286800
rect 66400 286500 66700 286800
rect 66900 286500 67200 286800
rect 67400 286500 67700 286800
rect 67900 286500 68200 286800
rect 68400 286500 68700 286800
rect 68900 286500 69200 286800
rect 69400 286500 69700 286800
rect 69900 286500 70200 286800
rect 70400 286500 70700 286800
rect 70900 286500 71200 286800
rect 71400 286500 71700 286800
rect 71900 286500 72200 286800
rect 72400 286500 72700 286800
rect 72900 286500 73200 286800
rect 73400 286500 73700 286800
rect 59400 286000 59700 286300
rect 59900 286000 60200 286300
rect 60400 286000 60700 286300
rect 60900 286000 61200 286300
rect 61400 286000 61700 286300
rect 61900 286000 62200 286300
rect 62400 286000 62700 286300
rect 62900 286000 63200 286300
rect 63400 286000 63700 286300
rect 63900 286000 64200 286300
rect 64400 286000 64700 286300
rect 64900 286000 65200 286300
rect 65400 286000 65700 286300
rect 65900 286000 66200 286300
rect 66400 286000 66700 286300
rect 66900 286000 67200 286300
rect 67400 286000 67700 286300
rect 67900 286000 68200 286300
rect 68400 286000 68700 286300
rect 68900 286000 69200 286300
rect 69400 286000 69700 286300
rect 69900 286000 70200 286300
rect 70400 286000 70700 286300
rect 70900 286000 71200 286300
rect 71400 286000 71700 286300
rect 71900 286000 72200 286300
rect 72400 286000 72700 286300
rect 72900 286000 73200 286300
rect 73400 286000 73700 286300
rect 21980 278310 22220 278550
rect 22320 278310 22560 278550
rect 21980 277950 22220 278190
rect 22320 277950 22560 278190
rect 34000 278100 34300 278400
rect 34400 278100 34700 278400
rect 34800 278100 35100 278400
rect 34460 275900 34700 276140
rect 37660 275900 37900 276140
rect 40980 275900 41220 276140
rect 12870 275220 13120 275470
rect 14520 273870 14780 274130
rect 16070 273870 16330 274130
rect 22850 273820 23100 274070
rect 12360 273060 12630 273330
rect 12870 273320 13120 273570
rect 21330 273560 21580 273810
rect 14000 273060 14270 273330
rect 15610 273280 15870 273540
rect 24320 273470 24560 273550
rect 24320 273390 24400 273470
rect 24400 273390 24480 273470
rect 24480 273390 24560 273470
rect 24320 273310 24560 273390
rect 24320 272950 24560 273030
rect 14520 272610 14780 272870
rect 16070 272610 16330 272870
rect 24320 272870 24400 272950
rect 24400 272870 24480 272950
rect 24480 272870 24560 272950
rect 24320 272790 24560 272870
rect 18710 272520 18970 272780
rect 20230 272520 20490 272780
rect 21750 272530 22000 272780
rect 23280 272530 23530 272780
rect 33980 272770 34220 273010
rect 34460 272770 34700 273010
rect 34940 272770 35180 273010
rect 37180 272770 37420 273010
rect 37660 272770 37900 273010
rect 38140 272770 38380 273010
rect 40500 272770 40740 273010
rect 40980 272770 41220 273010
rect 41460 272770 41700 273010
rect 24320 272430 24560 272510
rect 24320 272350 24400 272430
rect 24400 272350 24480 272430
rect 24480 272350 24560 272430
rect 12360 272010 12630 272280
rect 14000 272010 14270 272280
rect 24320 272270 24560 272350
rect 33980 272210 34220 272450
rect 34460 272210 34700 272450
rect 34940 272210 35180 272450
rect 37180 272210 37420 272450
rect 37660 272210 37900 272450
rect 38140 272210 38380 272450
rect 40500 272210 40740 272450
rect 40980 272210 41220 272450
rect 41460 272210 41700 272450
rect 12870 271740 13120 271990
rect 15610 271780 15870 272040
rect 24320 271930 24560 271990
rect 24320 271810 24380 271930
rect 24380 271810 24500 271930
rect 24500 271810 24560 271930
rect 14520 271340 14780 271600
rect 16070 271340 16330 271600
rect 21330 271500 21580 271750
rect 24320 271750 24560 271810
rect 22850 271240 23100 271490
rect 12860 269840 13110 270090
rect 34460 269200 34700 269440
rect 37660 269200 37900 269440
rect 40980 269200 41220 269440
rect 34000 268300 34300 268600
rect 34800 268300 35100 268600
rect 37300 268300 37600 268600
rect 38000 268300 38300 268600
rect 40600 268300 40900 268600
rect 41300 268300 41600 268600
rect 34000 267800 34300 268100
rect 34800 267800 35100 268100
rect 37300 267800 37600 268100
rect 38000 267800 38300 268100
rect 40600 267800 40900 268100
rect 41300 267800 41600 268100
rect 34000 267300 34300 267600
rect 34800 267300 35100 267600
rect 37300 267300 37600 267600
rect 38000 267300 38300 267600
rect 40600 267300 40900 267600
rect 41300 267300 41600 267600
rect 21980 267060 22220 267300
rect 22320 267060 22560 267300
rect 21980 266700 22220 266940
rect 22320 266700 22560 266940
rect 34000 266800 34300 267100
rect 34800 266800 35100 267100
rect 37300 266800 37600 267100
rect 38000 266800 38300 267100
rect 40600 266800 40900 267100
rect 41300 266800 41600 267100
rect 34000 266300 34300 266600
rect 34800 266300 35100 266600
rect 37300 266300 37600 266600
rect 38000 266300 38300 266600
rect 40600 266300 40900 266600
rect 41300 266300 41600 266600
rect 34000 265800 34300 266100
rect 34800 265800 35100 266100
rect 37300 265800 37600 266100
rect 38000 265800 38300 266100
rect 40600 265800 40900 266100
rect 41300 265800 41600 266100
rect 34000 265300 34300 265600
rect 34800 265300 35100 265600
rect 37300 265300 37600 265600
rect 38000 265300 38300 265600
rect 40600 265300 40900 265600
rect 41300 265300 41600 265600
rect 34000 264800 34300 265100
rect 34800 264800 35100 265100
rect 37300 264800 37600 265100
rect 38000 264800 38300 265100
rect 40600 264800 40900 265100
rect 41300 264800 41600 265100
rect 34000 264300 34300 264600
rect 34800 264300 35100 264600
rect 37300 264300 37600 264600
rect 38000 264300 38300 264600
rect 40600 264300 40900 264600
rect 41300 264300 41600 264600
rect 34000 263800 34300 264100
rect 34800 263800 35100 264100
rect 37300 263800 37600 264100
rect 38000 263800 38300 264100
rect 40600 263800 40900 264100
rect 41300 263800 41600 264100
rect 34000 263300 34300 263600
rect 34800 263300 35100 263600
rect 37300 263300 37600 263600
rect 38000 263300 38300 263600
rect 40600 263300 40900 263600
rect 41300 263300 41600 263600
rect 34000 262800 34300 263100
rect 34800 262800 35100 263100
rect 37300 262800 37600 263100
rect 38000 262800 38300 263100
rect 40600 262800 40900 263100
rect 41300 262800 41600 263100
rect 34000 262300 34300 262600
rect 34800 262300 35100 262600
rect 37300 262300 37600 262600
rect 38000 262300 38300 262600
rect 40600 262300 40900 262600
rect 41300 262300 41600 262600
rect 34000 261800 34300 262100
rect 34800 261800 35100 262100
rect 37300 261800 37600 262100
rect 38000 261800 38300 262100
rect 40600 261800 40900 262100
rect 41300 261800 41600 262100
rect 34000 261300 34300 261600
rect 34800 261300 35100 261600
rect 37300 261300 37600 261600
rect 38000 261300 38300 261600
rect 40600 261300 40900 261600
rect 41300 261300 41600 261600
rect 34000 260800 34300 261100
rect 34800 260800 35100 261100
rect 37300 260800 37600 261100
rect 38000 260800 38300 261100
rect 40600 260800 40900 261100
rect 41300 260800 41600 261100
rect 59500 252100 59800 252400
rect 60100 252100 60400 252400
rect 60700 252100 61000 252400
rect 61400 252100 61700 252400
rect 62000 252100 62300 252400
rect 62600 252100 62900 252400
rect 63200 252100 63500 252400
rect 63800 252100 64100 252400
rect 64400 252100 64700 252400
rect 65100 252100 65400 252400
rect 65700 252100 66000 252400
rect 66300 252100 66600 252400
rect 66900 252100 67200 252400
rect 67500 252100 67800 252400
rect 68100 252100 68400 252400
rect 68700 252100 69000 252400
rect 69300 252100 69600 252400
rect 69900 252100 70200 252400
rect 70600 252100 70900 252400
rect 71300 252100 71600 252400
rect 72000 252100 72300 252400
rect 72800 252100 73100 252400
rect 73500 252100 73800 252400
rect 59500 251400 59800 251700
rect 60100 251400 60400 251700
rect 60700 251400 61000 251700
rect 61400 251400 61700 251700
rect 62000 251400 62300 251700
rect 62600 251400 62900 251700
rect 63200 251400 63500 251700
rect 63800 251400 64100 251700
rect 64400 251400 64700 251700
rect 65100 251400 65400 251700
rect 65700 251400 66000 251700
rect 66300 251400 66600 251700
rect 66900 251400 67200 251700
rect 67500 251400 67800 251700
rect 68100 251400 68400 251700
rect 68700 251400 69000 251700
rect 69300 251400 69600 251700
rect 69900 251400 70200 251700
rect 70600 251400 70900 251700
rect 71300 251400 71600 251700
rect 72000 251400 72300 251700
rect 72800 251400 73100 251700
rect 73500 251400 73800 251700
rect 33900 241700 34200 242000
rect 34400 241700 34700 242000
rect 34900 241700 35200 242000
rect 33900 240900 34200 241200
rect 34400 240900 34700 241200
rect 34900 240900 35200 241200
rect 60000 218400 60400 218800
rect 60800 218400 61200 218800
rect 61600 218400 62000 218800
rect 62400 218400 62800 218800
rect 63200 218400 63600 218800
rect 64000 218400 64400 218800
rect 69000 218400 69400 218800
rect 69800 218400 70200 218800
rect 70600 218400 71000 218800
rect 71400 218400 71800 218800
rect 72200 218400 72600 218800
rect 73000 218400 73400 218800
rect 60000 217600 60400 218000
rect 60800 217600 61200 218000
rect 61600 217600 62000 218000
rect 62400 217600 62800 218000
rect 63200 217600 63600 218000
rect 64000 217600 64400 218000
rect 69000 217600 69400 218000
rect 69800 217600 70200 218000
rect 70600 217600 71000 218000
rect 71400 217600 71800 218000
rect 72200 217600 72600 218000
rect 73000 217600 73400 218000
rect 60000 216800 60400 217200
rect 60800 216800 61200 217200
rect 61600 216800 62000 217200
rect 62400 216800 62800 217200
rect 63200 216800 63600 217200
rect 64000 216800 64400 217200
rect 69000 216800 69400 217200
rect 69800 216800 70200 217200
rect 70600 216800 71000 217200
rect 71400 216800 71800 217200
rect 72200 216800 72600 217200
rect 73000 216800 73400 217200
rect 60000 216000 60400 216400
rect 60800 216000 61200 216400
rect 61600 216000 62000 216400
rect 62400 216000 62800 216400
rect 63200 216000 63600 216400
rect 64000 216000 64400 216400
rect 69000 216000 69400 216400
rect 69800 216000 70200 216400
rect 70600 216000 71000 216400
rect 71400 216000 71800 216400
rect 72200 216000 72600 216400
rect 73000 216000 73400 216400
rect 60000 215200 60400 215600
rect 60800 215200 61200 215600
rect 61600 215200 62000 215600
rect 62400 215200 62800 215600
rect 63200 215200 63600 215600
rect 64000 215200 64400 215600
rect 69000 215200 69400 215600
rect 69800 215200 70200 215600
rect 70600 215200 71000 215600
rect 71400 215200 71800 215600
rect 72200 215200 72600 215600
rect 73000 215200 73400 215600
rect 60000 214400 60400 214800
rect 60800 214400 61200 214800
rect 61600 214400 62000 214800
rect 62400 214400 62800 214800
rect 63200 214400 63600 214800
rect 64000 214400 64400 214800
rect 69000 214400 69400 214800
rect 69800 214400 70200 214800
rect 70600 214400 71000 214800
rect 71400 214400 71800 214800
rect 72200 214400 72600 214800
rect 73000 214400 73400 214800
rect 60000 209600 60400 210000
rect 60800 209600 61200 210000
rect 61600 209600 62000 210000
rect 62400 209600 62800 210000
rect 63200 209600 63600 210000
rect 64000 209600 64400 210000
rect 69000 209800 69400 210200
rect 69800 209800 70200 210200
rect 70600 209800 71000 210200
rect 71400 209800 71800 210200
rect 72200 209800 72600 210200
rect 73000 209800 73400 210200
rect 60000 208800 60400 209200
rect 60800 208800 61200 209200
rect 61600 208800 62000 209200
rect 62400 208800 62800 209200
rect 63200 208800 63600 209200
rect 64000 208800 64400 209200
rect 69000 209000 69400 209400
rect 69800 209000 70200 209400
rect 70600 209000 71000 209400
rect 71400 209000 71800 209400
rect 72200 209000 72600 209400
rect 73000 209000 73400 209400
rect 60000 208000 60400 208400
rect 60800 208000 61200 208400
rect 61600 208000 62000 208400
rect 62400 208000 62800 208400
rect 63200 208000 63600 208400
rect 64000 208000 64400 208400
rect 69000 208200 69400 208600
rect 69800 208200 70200 208600
rect 70600 208200 71000 208600
rect 71400 208200 71800 208600
rect 72200 208200 72600 208600
rect 73000 208200 73400 208600
rect 60000 207200 60400 207600
rect 60800 207200 61200 207600
rect 61600 207200 62000 207600
rect 62400 207200 62800 207600
rect 63200 207200 63600 207600
rect 64000 207200 64400 207600
rect 69000 207400 69400 207800
rect 69800 207400 70200 207800
rect 70600 207400 71000 207800
rect 71400 207400 71800 207800
rect 72200 207400 72600 207800
rect 73000 207400 73400 207800
rect 60000 206400 60400 206800
rect 60800 206400 61200 206800
rect 61600 206400 62000 206800
rect 62400 206400 62800 206800
rect 63200 206400 63600 206800
rect 64000 206400 64400 206800
rect 69000 206600 69400 207000
rect 69800 206600 70200 207000
rect 70600 206600 71000 207000
rect 71400 206600 71800 207000
rect 72200 206600 72600 207000
rect 73000 206600 73400 207000
rect 60000 205600 60400 206000
rect 60800 205600 61200 206000
rect 61600 205600 62000 206000
rect 62400 205600 62800 206000
rect 63200 205600 63600 206000
rect 64000 205600 64400 206000
rect 69000 205800 69400 206200
rect 69800 205800 70200 206200
rect 70600 205800 71000 206200
rect 71400 205800 71800 206200
rect 72200 205800 72600 206200
rect 73000 205800 73400 206200
rect 285400 219000 285800 219400
rect 286200 219000 286600 219400
rect 287000 219000 287400 219400
rect 287800 219000 288200 219400
rect 288600 219000 289000 219400
rect 289400 219000 289800 219400
rect 285400 218200 285800 218600
rect 286200 218200 286600 218600
rect 287000 218200 287400 218600
rect 287800 218200 288200 218600
rect 288600 218200 289000 218600
rect 289400 218200 289800 218600
rect 285400 217400 285800 217800
rect 286200 217400 286600 217800
rect 287000 217400 287400 217800
rect 287800 217400 288200 217800
rect 288600 217400 289000 217800
rect 289400 217400 289800 217800
rect 285400 216600 285800 217000
rect 286200 216600 286600 217000
rect 287000 216600 287400 217000
rect 287800 216600 288200 217000
rect 288600 216600 289000 217000
rect 289400 216600 289800 217000
rect 285400 215800 285800 216200
rect 286200 215800 286600 216200
rect 287000 215800 287400 216200
rect 287800 215800 288200 216200
rect 288600 215800 289000 216200
rect 289400 215800 289800 216200
rect 285400 215000 285800 215400
rect 286200 215000 286600 215400
rect 287000 215000 287400 215400
rect 287800 215000 288200 215400
rect 288600 215000 289000 215400
rect 289400 215000 289800 215400
rect 285200 214200 285600 214600
rect 286000 214200 286400 214600
rect 286800 214200 287200 214600
rect 287600 214200 288000 214600
rect 288400 214200 288800 214600
rect 289200 214200 289600 214600
rect 285200 213400 285600 213800
rect 286000 213400 286400 213800
rect 286800 213400 287200 213800
rect 287600 213400 288000 213800
rect 288400 213400 288800 213800
rect 289200 213400 289600 213800
rect 285200 212600 285600 213000
rect 286000 212600 286400 213000
rect 286800 212600 287200 213000
rect 287600 212600 288000 213000
rect 288400 212600 288800 213000
rect 289200 212600 289600 213000
rect 285200 211800 285600 212200
rect 286000 211800 286400 212200
rect 286800 211800 287200 212200
rect 287600 211800 288000 212200
rect 288400 211800 288800 212200
rect 289200 211800 289600 212200
rect 285200 211000 285600 211400
rect 286000 211000 286400 211400
rect 286800 211000 287200 211400
rect 287600 211000 288000 211400
rect 288400 211000 288800 211400
rect 289200 211000 289600 211400
rect 285200 210200 285600 210600
rect 286000 210200 286400 210600
rect 286800 210200 287200 210600
rect 287600 210200 288000 210600
rect 288400 210200 288800 210600
rect 289200 210200 289600 210600
rect 285200 209400 285600 209800
rect 286000 209400 286400 209800
rect 286800 209400 287200 209800
rect 287600 209400 288000 209800
rect 288400 209400 288800 209800
rect 289200 209400 289600 209800
rect 285200 208600 285600 209000
rect 286000 208600 286400 209000
rect 286800 208600 287200 209000
rect 287600 208600 288000 209000
rect 288400 208600 288800 209000
rect 289200 208600 289600 209000
rect 285200 207800 285600 208200
rect 286000 207800 286400 208200
rect 286800 207800 287200 208200
rect 287600 207800 288000 208200
rect 288400 207800 288800 208200
rect 289200 207800 289600 208200
rect 285200 207000 285600 207400
rect 286000 207000 286400 207400
rect 286800 207000 287200 207400
rect 287600 207000 288000 207400
rect 288400 207000 288800 207400
rect 289200 207000 289600 207400
rect 285200 206200 285600 206600
rect 286000 206200 286400 206600
rect 286800 206200 287200 206600
rect 287600 206200 288000 206600
rect 288400 206200 288800 206600
rect 289200 206200 289600 206600
rect 285200 205400 285600 205800
rect 286000 205400 286400 205800
rect 286800 205400 287200 205800
rect 287600 205400 288000 205800
rect 288400 205400 288800 205800
rect 289200 205400 289600 205800
rect 545900 288600 546200 288900
rect 546400 288600 546700 288900
rect 546900 288600 547200 288900
rect 547400 288600 547700 288900
rect 547900 288600 548200 288900
rect 548400 288600 548700 288900
rect 545900 288100 546200 288400
rect 546400 288100 546700 288400
rect 546900 288100 547200 288400
rect 547400 288100 547700 288400
rect 547900 288100 548200 288400
rect 548400 288100 548700 288400
rect 545900 287600 546200 287900
rect 546400 287600 546700 287900
rect 546900 287600 547200 287900
rect 547400 287600 547700 287900
rect 547900 287600 548200 287900
rect 548400 287600 548700 287900
rect 569200 288600 569500 288900
rect 569800 288600 570100 288900
rect 569200 288100 569500 288400
rect 569800 288100 570100 288400
rect 572800 288400 573100 288700
rect 573300 288400 573600 288700
rect 573800 288400 574100 288700
rect 574300 288400 574600 288700
rect 569200 287600 569500 287900
rect 569800 287600 570100 287900
rect 572800 287900 573100 288200
rect 573300 287900 573600 288200
rect 573800 287900 574100 288200
rect 574300 287900 574600 288200
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 549700 684900 578640 685100
rect 549700 684600 549900 684900
rect 550200 684600 550400 684900
rect 550700 684600 550900 684900
rect 551200 684600 551400 684900
rect 551700 684600 551900 684900
rect 552200 684600 552400 684900
rect 552700 684600 573200 684900
rect 573500 684600 573800 684900
rect 574100 684700 578640 684900
rect 574100 684600 576800 684700
rect 549700 684400 576800 684600
rect 577100 684400 577300 684700
rect 577600 684400 577800 684700
rect 578100 684400 578300 684700
rect 578600 684400 578640 684700
rect 549700 684100 549900 684400
rect 550200 684100 550400 684400
rect 550700 684100 550900 684400
rect 551200 684100 551400 684400
rect 551700 684100 551900 684400
rect 552200 684100 552400 684400
rect 552700 684100 573200 684400
rect 573500 684100 573800 684400
rect 574100 684200 578640 684400
rect 574100 684100 576800 684200
rect 549700 683900 576800 684100
rect 577100 683900 577300 684200
rect 577600 683900 577800 684200
rect 578100 683900 578300 684200
rect 578600 683900 578640 684200
rect 549700 683600 549900 683900
rect 550200 683600 550400 683900
rect 550700 683600 550900 683900
rect 551200 683600 551400 683900
rect 551700 683600 551900 683900
rect 552200 683600 552400 683900
rect 552700 683600 573200 683900
rect 573500 683600 573800 683900
rect 574100 683600 578640 683900
rect 549700 683400 578640 683600
rect 12800 674100 51300 674200
rect 12800 673800 12900 674100
rect 13200 673800 13700 674100
rect 14000 674000 51300 674100
rect 14000 673800 32800 674000
rect 12800 673700 32800 673800
rect 33100 673700 33300 674000
rect 33600 673700 33800 674000
rect 34100 673700 34300 674000
rect 34600 673700 34800 674000
rect 35100 673700 35300 674000
rect 35600 673700 35800 674000
rect 36100 673700 36300 674000
rect 36600 673700 36800 674000
rect 37100 673700 37300 674000
rect 37600 673700 37800 674000
rect 38100 673700 38300 674000
rect 38600 673700 38800 674000
rect 39100 673700 39300 674000
rect 39600 673700 39800 674000
rect 40100 673700 40300 674000
rect 40600 673700 50100 674000
rect 50400 673700 51300 674000
rect 12800 673600 51300 673700
rect 12800 673300 12900 673600
rect 13200 673300 13700 673600
rect 14000 673300 50100 673600
rect 50400 673300 51300 673600
rect 12800 673200 51300 673300
rect 12800 673100 32800 673200
rect 12800 672800 12900 673100
rect 13200 672800 13700 673100
rect 14000 672900 32800 673100
rect 33100 672900 33300 673200
rect 33600 672900 33800 673200
rect 34100 672900 34300 673200
rect 34600 672900 34800 673200
rect 35100 672900 35300 673200
rect 35600 672900 35800 673200
rect 36100 672900 36300 673200
rect 36600 672900 36800 673200
rect 37100 672900 37300 673200
rect 37600 672900 37800 673200
rect 38100 672900 38300 673200
rect 38600 672900 38800 673200
rect 39100 672900 39300 673200
rect 39600 672900 39800 673200
rect 40100 672900 40300 673200
rect 40600 672900 50100 673200
rect 50400 672900 51300 673200
rect 14000 672800 51300 672900
rect 12800 672700 51300 672800
rect 32600 670700 48300 670900
rect 32600 670400 32800 670700
rect 33100 670400 33300 670700
rect 33600 670400 33800 670700
rect 34100 670400 34300 670700
rect 34600 670400 34800 670700
rect 35100 670400 35300 670700
rect 35600 670400 35800 670700
rect 36100 670400 36300 670700
rect 36600 670400 36800 670700
rect 37100 670400 37300 670700
rect 37600 670400 37800 670700
rect 38100 670400 38300 670700
rect 38600 670400 38800 670700
rect 39100 670400 39300 670700
rect 39600 670400 39800 670700
rect 40100 670400 40300 670700
rect 40600 670400 48300 670700
rect 32600 670000 48300 670400
rect 32600 669700 32800 670000
rect 33100 669700 33300 670000
rect 33600 669700 33800 670000
rect 34100 669700 34300 670000
rect 34600 669700 34800 670000
rect 35100 669700 35300 670000
rect 35600 669700 35800 670000
rect 36100 669700 36300 670000
rect 36600 669700 36800 670000
rect 37100 669700 37300 670000
rect 37600 669700 37800 670000
rect 38100 669700 38300 670000
rect 38600 669700 38800 670000
rect 39100 669700 39300 670000
rect 39600 669700 39800 670000
rect 40100 669700 40300 670000
rect 40600 669700 48300 670000
rect 32600 669500 48300 669700
rect 32600 667400 48300 667600
rect 32600 667100 32800 667400
rect 33100 667100 33300 667400
rect 33600 667100 33800 667400
rect 34100 667100 34300 667400
rect 34600 667100 34800 667400
rect 35100 667100 35300 667400
rect 35600 667100 35800 667400
rect 36100 667100 36300 667400
rect 36600 667100 36800 667400
rect 37100 667100 37300 667400
rect 37600 667100 37800 667400
rect 38100 667100 38300 667400
rect 38600 667100 38800 667400
rect 39100 667100 39300 667400
rect 39600 667100 39800 667400
rect 40100 667100 40300 667400
rect 40600 667100 48300 667400
rect 32600 666700 48300 667100
rect 32600 666400 32800 666700
rect 33100 666400 33300 666700
rect 33600 666400 33800 666700
rect 34100 666400 34300 666700
rect 34600 666400 34800 666700
rect 35100 666400 35300 666700
rect 35600 666400 35800 666700
rect 36100 666400 36300 666700
rect 36600 666400 36800 666700
rect 37100 666400 37300 666700
rect 37600 666400 37800 666700
rect 38100 666400 38300 666700
rect 38600 666400 38800 666700
rect 39100 666400 39300 666700
rect 39600 666400 39800 666700
rect 40100 666400 40300 666700
rect 40600 666400 48300 666700
rect 32600 666200 48300 666400
rect 2300 648600 62200 648800
rect 2300 648300 2500 648600
rect 2800 648300 3000 648600
rect 3300 648300 3500 648600
rect 3800 648500 58000 648600
rect 3800 648300 23400 648500
rect 2300 648200 23400 648300
rect 23700 648200 24100 648500
rect 24400 648300 58000 648500
rect 58300 648300 58500 648600
rect 58800 648300 59000 648600
rect 59300 648300 59500 648600
rect 59800 648300 60000 648600
rect 60300 648300 60500 648600
rect 60800 648300 61000 648600
rect 61300 648300 61500 648600
rect 61800 648300 62200 648600
rect 24400 648200 62200 648300
rect 2300 648100 62200 648200
rect 2300 647800 2500 648100
rect 2800 647800 3000 648100
rect 3300 647800 3500 648100
rect 3800 647900 58000 648100
rect 3800 647800 23400 647900
rect 2300 647600 23400 647800
rect 23700 647600 24100 647900
rect 24400 647800 58000 647900
rect 58300 647800 58500 648100
rect 58800 647800 59000 648100
rect 59300 647800 59500 648100
rect 59800 647800 60000 648100
rect 60300 647800 60500 648100
rect 60800 647800 61000 648100
rect 61300 647800 61500 648100
rect 61800 647800 62200 648100
rect 24400 647600 62200 647800
rect 2300 647300 2500 647600
rect 2800 647300 3000 647600
rect 3300 647300 3500 647600
rect 3800 647300 58000 647600
rect 58300 647300 58500 647600
rect 58800 647300 59000 647600
rect 59300 647300 59500 647600
rect 59800 647300 60000 647600
rect 60300 647300 60500 647600
rect 60800 647300 61000 647600
rect 61300 647300 61500 647600
rect 61800 647300 62200 647600
rect 2300 647100 23400 647300
rect 2300 646800 2500 647100
rect 2800 646800 3000 647100
rect 3300 646800 3500 647100
rect 3800 647000 23400 647100
rect 23700 647000 24100 647300
rect 24400 647100 62200 647300
rect 24400 647000 58000 647100
rect 3800 646800 58000 647000
rect 58300 646800 58500 647100
rect 58800 646800 59000 647100
rect 59300 646800 59500 647100
rect 59800 646800 60000 647100
rect 60300 646800 60500 647100
rect 60800 646800 61000 647100
rect 61300 646800 61500 647100
rect 61800 646800 62200 647100
rect 2300 646600 62200 646800
rect 2300 646300 2500 646600
rect 2800 646300 3000 646600
rect 3300 646300 3500 646600
rect 3800 646300 23400 646600
rect 23700 646300 24100 646600
rect 24400 646300 58000 646600
rect 58300 646300 58500 646600
rect 58800 646300 59000 646600
rect 59300 646300 59500 646600
rect 59800 646300 60000 646600
rect 60300 646300 60500 646600
rect 60800 646300 61000 646600
rect 61300 646300 61500 646600
rect 61800 646300 62200 646600
rect 2300 646100 62200 646300
rect 2300 645800 2500 646100
rect 2800 645800 3000 646100
rect 3300 645800 3500 646100
rect 3800 646000 58000 646100
rect 3800 645800 23400 646000
rect 2300 645700 23400 645800
rect 23700 645700 24100 646000
rect 24400 645800 58000 646000
rect 58300 645800 58500 646100
rect 58800 645800 59000 646100
rect 59300 645800 59500 646100
rect 59800 645800 60000 646100
rect 60300 645800 60500 646100
rect 60800 645800 61000 646100
rect 61300 645800 61500 646100
rect 61800 645800 62200 646100
rect 24400 645700 62200 645800
rect 2300 645600 62200 645700
rect 2300 645300 2500 645600
rect 2800 645300 3000 645600
rect 3300 645300 3500 645600
rect 3800 645400 58000 645600
rect 3800 645300 23400 645400
rect 2300 645100 23400 645300
rect 23700 645100 24100 645400
rect 24400 645300 58000 645400
rect 58300 645300 58500 645600
rect 58800 645300 59000 645600
rect 59300 645300 59500 645600
rect 59800 645300 60000 645600
rect 60300 645300 60500 645600
rect 60800 645300 61000 645600
rect 61300 645300 61500 645600
rect 61800 645300 62200 645600
rect 24400 645100 62200 645300
rect 2300 644800 2500 645100
rect 2800 644800 3000 645100
rect 3300 644800 3500 645100
rect 3800 644800 58000 645100
rect 58300 644800 58500 645100
rect 58800 644800 59000 645100
rect 59300 644800 59500 645100
rect 59800 644800 60000 645100
rect 60300 644800 60500 645100
rect 60800 644800 61000 645100
rect 61300 644800 61500 645100
rect 61800 644800 62200 645100
rect 2300 644600 23400 644800
rect 2300 644300 2500 644600
rect 2800 644300 3000 644600
rect 3300 644300 3500 644600
rect 3800 644500 23400 644600
rect 23700 644500 24100 644800
rect 24400 644600 62200 644800
rect 24400 644500 58000 644600
rect 3800 644300 58000 644500
rect 58300 644300 58500 644600
rect 58800 644300 59000 644600
rect 59300 644300 59500 644600
rect 59800 644300 60000 644600
rect 60300 644300 60500 644600
rect 60800 644300 61000 644600
rect 61300 644300 61500 644600
rect 61800 644300 62200 644600
rect 2300 644200 62200 644300
rect 2300 644100 23400 644200
rect 2300 643800 2500 644100
rect 2800 643800 3000 644100
rect 3300 643800 3500 644100
rect 3800 643900 23400 644100
rect 23700 643900 24100 644200
rect 24400 644100 62200 644200
rect 24400 643900 58000 644100
rect 3800 643800 58000 643900
rect 58300 643800 58500 644100
rect 58800 643800 59000 644100
rect 59300 643800 59500 644100
rect 59800 643800 60000 644100
rect 60300 643800 60500 644100
rect 60800 643800 61000 644100
rect 61300 643800 61500 644100
rect 61800 643800 62200 644100
rect 2300 643600 62200 643800
rect 2300 643300 2500 643600
rect 2800 643300 3000 643600
rect 3300 643300 3500 643600
rect 3800 643300 23400 643600
rect 23700 643300 24100 643600
rect 24400 643300 58000 643600
rect 58300 643300 58500 643600
rect 58800 643300 59000 643600
rect 59300 643300 59500 643600
rect 59800 643300 60000 643600
rect 60300 643300 60500 643600
rect 60800 643300 61000 643600
rect 61300 643300 61500 643600
rect 61800 643300 62200 643600
rect 2300 643100 62200 643300
rect 2300 642800 2500 643100
rect 2800 642800 3000 643100
rect 3300 642800 3500 643100
rect 3800 642900 58000 643100
rect 3800 642800 23400 642900
rect 2300 642600 23400 642800
rect 23700 642600 24100 642900
rect 24400 642800 58000 642900
rect 58300 642800 58500 643100
rect 58800 642800 59000 643100
rect 59300 642800 59500 643100
rect 59800 642800 60000 643100
rect 60300 642800 60500 643100
rect 60800 642800 61000 643100
rect 61300 642800 61500 643100
rect 61800 642800 62200 643100
rect 24400 642600 62200 642800
rect 2300 642300 2500 642600
rect 2800 642300 3000 642600
rect 3300 642300 3500 642600
rect 3800 642300 58000 642600
rect 58300 642300 58500 642600
rect 58800 642300 59000 642600
rect 59300 642300 59500 642600
rect 59800 642300 60000 642600
rect 60300 642300 60500 642600
rect 60800 642300 61000 642600
rect 61300 642300 61500 642600
rect 61800 642300 62200 642600
rect 2300 642100 23400 642300
rect 2300 641800 2500 642100
rect 2800 641800 3000 642100
rect 3300 641800 3500 642100
rect 3800 642000 23400 642100
rect 23700 642000 24100 642300
rect 24400 642100 62200 642300
rect 24400 642000 58000 642100
rect 3800 641800 58000 642000
rect 58300 641800 58500 642100
rect 58800 641800 59000 642100
rect 59300 641800 59500 642100
rect 59800 641800 60000 642100
rect 60300 641800 60500 642100
rect 60800 641800 61000 642100
rect 61300 641800 61500 642100
rect 61800 641800 62200 642100
rect 2300 641700 62200 641800
rect 2300 641600 23400 641700
rect 2300 641300 2500 641600
rect 2800 641300 3000 641600
rect 3300 641300 3500 641600
rect 3800 641400 23400 641600
rect 23700 641400 24100 641700
rect 24400 641600 62200 641700
rect 24400 641400 58000 641600
rect 3800 641300 58000 641400
rect 58300 641300 58500 641600
rect 58800 641300 59000 641600
rect 59300 641300 59500 641600
rect 59800 641300 60000 641600
rect 60300 641300 60500 641600
rect 60800 641300 61000 641600
rect 61300 641300 61500 641600
rect 61800 641300 62200 641600
rect 2300 641100 62200 641300
rect 2300 640800 2500 641100
rect 2800 640800 3000 641100
rect 3300 640800 3500 641100
rect 3800 640800 23400 641100
rect 23700 640800 24100 641100
rect 24400 640800 58000 641100
rect 58300 640800 58500 641100
rect 58800 640800 59000 641100
rect 59300 640800 59500 641100
rect 59800 640800 60000 641100
rect 60300 640800 60500 641100
rect 60800 640800 61000 641100
rect 61300 640800 61500 641100
rect 61800 640800 62200 641100
rect 2300 640600 62200 640800
rect 2300 640300 2500 640600
rect 2800 640300 3000 640600
rect 3300 640300 3500 640600
rect 3800 640500 58000 640600
rect 3800 640300 23400 640500
rect 2300 640200 23400 640300
rect 23700 640200 24100 640500
rect 24400 640300 58000 640500
rect 58300 640300 58500 640600
rect 58800 640300 59000 640600
rect 59300 640300 59500 640600
rect 59800 640300 60000 640600
rect 60300 640300 60500 640600
rect 60800 640300 61000 640600
rect 61300 640300 61500 640600
rect 61800 640300 62200 640600
rect 24400 640200 62200 640300
rect 2300 640100 62200 640200
rect 2300 639800 2500 640100
rect 2800 639800 3000 640100
rect 3300 639800 3500 640100
rect 3800 639900 58000 640100
rect 3800 639800 23400 639900
rect 2300 639600 23400 639800
rect 23700 639600 24100 639900
rect 24400 639800 58000 639900
rect 58300 639800 58500 640100
rect 58800 639800 59000 640100
rect 59300 639800 59500 640100
rect 59800 639800 60000 640100
rect 60300 639800 60500 640100
rect 60800 639800 61000 640100
rect 61300 639800 61500 640100
rect 61800 639800 62200 640100
rect 24400 639600 62200 639800
rect 2300 639300 2500 639600
rect 2800 639300 3000 639600
rect 3300 639300 3500 639600
rect 3800 639300 58000 639600
rect 58300 639300 58500 639600
rect 58800 639300 59000 639600
rect 59300 639300 59500 639600
rect 59800 639300 60000 639600
rect 60300 639300 60500 639600
rect 60800 639300 61000 639600
rect 61300 639300 61500 639600
rect 61800 639300 62200 639600
rect 2300 639100 23400 639300
rect 2300 638800 2500 639100
rect 2800 638800 3000 639100
rect 3300 638800 3500 639100
rect 3800 639000 23400 639100
rect 23700 639000 24100 639300
rect 24400 639100 62200 639300
rect 24400 639000 58000 639100
rect 3800 638800 58000 639000
rect 58300 638800 58500 639100
rect 58800 638800 59000 639100
rect 59300 638800 59500 639100
rect 59800 638800 60000 639100
rect 60300 638800 60500 639100
rect 60800 638800 61000 639100
rect 61300 638800 61500 639100
rect 61800 638800 62200 639100
rect 2300 638700 62200 638800
rect 2300 638600 23400 638700
rect 2300 638300 2500 638600
rect 2800 638300 3000 638600
rect 3300 638300 3500 638600
rect 3800 638400 23400 638600
rect 23700 638400 24100 638700
rect 24400 638600 62200 638700
rect 24400 638400 58000 638600
rect 3800 638300 58000 638400
rect 58300 638300 58500 638600
rect 58800 638300 59000 638600
rect 59300 638300 59500 638600
rect 59800 638300 60000 638600
rect 60300 638300 60500 638600
rect 60800 638300 61000 638600
rect 61300 638300 61500 638600
rect 61800 638300 62200 638600
rect 2300 638100 62200 638300
rect 2300 637800 2500 638100
rect 2800 637800 3000 638100
rect 3300 637800 3500 638100
rect 3800 637800 23400 638100
rect 23700 637800 24100 638100
rect 24400 637800 58000 638100
rect 58300 637800 58500 638100
rect 58800 637800 59000 638100
rect 59300 637800 59500 638100
rect 59800 637800 60000 638100
rect 60300 637800 60500 638100
rect 60800 637800 61000 638100
rect 61300 637800 61500 638100
rect 61800 637800 62200 638100
rect 2300 637600 62200 637800
rect 2300 637300 2500 637600
rect 2800 637300 3000 637600
rect 3300 637300 3500 637600
rect 3800 637400 58000 637600
rect 3800 637300 23400 637400
rect 2300 637100 23400 637300
rect 23700 637100 24100 637400
rect 24400 637300 58000 637400
rect 58300 637300 58500 637600
rect 58800 637300 59000 637600
rect 59300 637300 59500 637600
rect 59800 637300 60000 637600
rect 60300 637300 60500 637600
rect 60800 637300 61000 637600
rect 61300 637300 61500 637600
rect 61800 637300 62200 637600
rect 24400 637100 62200 637300
rect 2300 636800 2500 637100
rect 2800 636800 3000 637100
rect 3300 636800 3500 637100
rect 3800 636800 58000 637100
rect 58300 636800 58500 637100
rect 58800 636800 59000 637100
rect 59300 636800 59500 637100
rect 59800 636800 60000 637100
rect 60300 636800 60500 637100
rect 60800 636800 61000 637100
rect 61300 636800 61500 637100
rect 61800 636800 62200 637100
rect 2300 636700 62200 636800
rect 2300 636600 23400 636700
rect 2300 636300 2500 636600
rect 2800 636300 3000 636600
rect 3300 636300 3500 636600
rect 3800 636400 23400 636600
rect 23700 636400 24100 636700
rect 24400 636600 62200 636700
rect 24400 636400 58000 636600
rect 3800 636300 58000 636400
rect 58300 636300 58500 636600
rect 58800 636300 59000 636600
rect 59300 636300 59500 636600
rect 59800 636300 60000 636600
rect 60300 636300 60500 636600
rect 60800 636300 61000 636600
rect 61300 636300 61500 636600
rect 61800 636300 62200 636600
rect 2300 636100 62200 636300
rect 2300 635800 2500 636100
rect 2800 635800 3000 636100
rect 3300 635800 3500 636100
rect 3800 636000 58000 636100
rect 3800 635800 23400 636000
rect 2300 635700 23400 635800
rect 23700 635700 24100 636000
rect 24400 635800 58000 636000
rect 58300 635800 58500 636100
rect 58800 635800 59000 636100
rect 59300 635800 59500 636100
rect 59800 635800 60000 636100
rect 60300 635800 60500 636100
rect 60800 635800 61000 636100
rect 61300 635800 61500 636100
rect 61800 635800 62200 636100
rect 24400 635700 62200 635800
rect 2300 635600 62200 635700
rect 2300 635300 2500 635600
rect 2800 635300 3000 635600
rect 3300 635300 3500 635600
rect 3800 635300 58000 635600
rect 58300 635300 58500 635600
rect 58800 635300 59000 635600
rect 59300 635300 59500 635600
rect 59800 635300 60000 635600
rect 60300 635300 60500 635600
rect 60800 635300 61000 635600
rect 61300 635300 61500 635600
rect 61800 635300 62200 635600
rect 2300 635200 62200 635300
rect 2300 635100 23400 635200
rect 2300 634800 2500 635100
rect 2800 634800 3000 635100
rect 3300 634800 3500 635100
rect 3800 634900 23400 635100
rect 23700 634900 24100 635200
rect 24400 635100 62200 635200
rect 24400 634900 58000 635100
rect 3800 634800 58000 634900
rect 58300 634800 58500 635100
rect 58800 634800 59000 635100
rect 59300 634800 59500 635100
rect 59800 634800 60000 635100
rect 60300 634800 60500 635100
rect 60800 634800 61000 635100
rect 61300 634800 61500 635100
rect 61800 634800 62200 635100
rect 2300 634600 62200 634800
rect 2300 634300 2500 634600
rect 2800 634300 3000 634600
rect 3300 634300 3500 634600
rect 3800 634500 58000 634600
rect 3800 634300 23400 634500
rect 2300 634200 23400 634300
rect 23700 634200 24100 634500
rect 24400 634300 58000 634500
rect 58300 634300 58500 634600
rect 58800 634300 59000 634600
rect 59300 634300 59500 634600
rect 59800 634300 60000 634600
rect 60300 634300 60500 634600
rect 60800 634300 61000 634600
rect 61300 634300 61500 634600
rect 61800 634300 62200 634600
rect 24400 634200 62200 634300
rect 2300 633800 62200 634200
rect 289500 344400 306000 344600
rect 289500 344100 289600 344400
rect 289900 344300 306000 344400
rect 289900 344200 299000 344300
rect 289900 344100 294800 344200
rect 289500 343900 294800 344100
rect 295100 343900 299000 344200
rect 299400 343900 299600 344300
rect 300000 343900 300200 344300
rect 300600 343900 300800 344300
rect 301200 343900 301400 344300
rect 301800 343900 302000 344300
rect 302400 343900 302600 344300
rect 303000 343900 303200 344300
rect 303600 343900 306000 344300
rect 289500 343600 289600 343900
rect 289900 343700 306000 343900
rect 289900 343600 299000 343700
rect 289500 343400 299000 343600
rect 289500 343100 289600 343400
rect 289900 343300 299000 343400
rect 299400 343300 299600 343700
rect 300000 343300 300200 343700
rect 300600 343300 300800 343700
rect 301200 343300 301400 343700
rect 301800 343300 302000 343700
rect 302400 343300 302600 343700
rect 303000 343300 303200 343700
rect 303600 343300 306000 343700
rect 289900 343100 306000 343300
rect 289500 342900 306000 343100
rect 287200 342300 288600 342400
rect 287200 342000 287500 342300
rect 287800 342000 288000 342300
rect 288300 342000 288600 342300
rect 287200 340824 288600 342000
rect 287200 340800 288624 340824
rect 287200 340500 288300 340800
rect 288600 340500 288624 340800
rect 287200 340476 288624 340500
rect 287200 338500 288600 340476
rect 59200 289800 74200 290200
rect 59200 289500 59400 289800
rect 59700 289500 59900 289800
rect 60200 289500 60400 289800
rect 60700 289500 60900 289800
rect 61200 289500 61400 289800
rect 61700 289500 61900 289800
rect 62200 289500 62400 289800
rect 62700 289500 62900 289800
rect 63200 289500 63400 289800
rect 63700 289500 63900 289800
rect 64200 289500 64400 289800
rect 64700 289500 64900 289800
rect 65200 289500 65400 289800
rect 65700 289500 65900 289800
rect 66200 289500 66400 289800
rect 66700 289500 66900 289800
rect 67200 289500 67400 289800
rect 67700 289500 67900 289800
rect 68200 289500 68400 289800
rect 68700 289500 68900 289800
rect 69200 289500 69400 289800
rect 69700 289500 69900 289800
rect 70200 289500 70400 289800
rect 70700 289500 70900 289800
rect 71200 289500 71400 289800
rect 71700 289500 71900 289800
rect 72200 289500 72400 289800
rect 72700 289500 72900 289800
rect 73200 289500 73400 289800
rect 73700 289500 74200 289800
rect 59200 289300 74200 289500
rect 59200 289000 59400 289300
rect 59700 289000 59900 289300
rect 60200 289000 60400 289300
rect 60700 289000 60900 289300
rect 61200 289000 61400 289300
rect 61700 289000 61900 289300
rect 62200 289000 62400 289300
rect 62700 289000 62900 289300
rect 63200 289000 63400 289300
rect 63700 289000 63900 289300
rect 64200 289000 64400 289300
rect 64700 289000 64900 289300
rect 65200 289000 65400 289300
rect 65700 289000 65900 289300
rect 66200 289000 66400 289300
rect 66700 289000 66900 289300
rect 67200 289000 67400 289300
rect 67700 289000 67900 289300
rect 68200 289000 68400 289300
rect 68700 289000 68900 289300
rect 69200 289000 69400 289300
rect 69700 289000 69900 289300
rect 70200 289000 70400 289300
rect 70700 289000 70900 289300
rect 71200 289000 71400 289300
rect 71700 289000 71900 289300
rect 72200 289000 72400 289300
rect 72700 289000 72900 289300
rect 73200 289000 73400 289300
rect 73700 289000 74200 289300
rect 59200 288800 74200 289000
rect 59200 288500 59400 288800
rect 59700 288500 59900 288800
rect 60200 288500 60400 288800
rect 60700 288500 60900 288800
rect 61200 288500 61400 288800
rect 61700 288500 61900 288800
rect 62200 288500 62400 288800
rect 62700 288500 62900 288800
rect 63200 288500 63400 288800
rect 63700 288500 63900 288800
rect 64200 288500 64400 288800
rect 64700 288500 64900 288800
rect 65200 288500 65400 288800
rect 65700 288500 65900 288800
rect 66200 288500 66400 288800
rect 66700 288500 66900 288800
rect 67200 288500 67400 288800
rect 67700 288500 67900 288800
rect 68200 288500 68400 288800
rect 68700 288500 68900 288800
rect 69200 288500 69400 288800
rect 69700 288500 69900 288800
rect 70200 288500 70400 288800
rect 70700 288500 70900 288800
rect 71200 288500 71400 288800
rect 71700 288500 71900 288800
rect 72200 288500 72400 288800
rect 72700 288500 72900 288800
rect 73200 288500 73400 288800
rect 73700 288500 74200 288800
rect 59200 288300 74200 288500
rect 59200 288000 59400 288300
rect 59700 288000 59900 288300
rect 60200 288000 60400 288300
rect 60700 288000 60900 288300
rect 61200 288000 61400 288300
rect 61700 288000 61900 288300
rect 62200 288000 62400 288300
rect 62700 288000 62900 288300
rect 63200 288000 63400 288300
rect 63700 288000 63900 288300
rect 64200 288000 64400 288300
rect 64700 288000 64900 288300
rect 65200 288000 65400 288300
rect 65700 288000 65900 288300
rect 66200 288000 66400 288300
rect 66700 288000 66900 288300
rect 67200 288000 67400 288300
rect 67700 288000 67900 288300
rect 68200 288000 68400 288300
rect 68700 288000 68900 288300
rect 69200 288000 69400 288300
rect 69700 288000 69900 288300
rect 70200 288000 70400 288300
rect 70700 288000 70900 288300
rect 71200 288000 71400 288300
rect 71700 288000 71900 288300
rect 72200 288000 72400 288300
rect 72700 288000 72900 288300
rect 73200 288000 73400 288300
rect 73700 288000 74200 288300
rect 59200 287800 74200 288000
rect 59200 287500 59400 287800
rect 59700 287500 59900 287800
rect 60200 287500 60400 287800
rect 60700 287500 60900 287800
rect 61200 287500 61400 287800
rect 61700 287500 61900 287800
rect 62200 287500 62400 287800
rect 62700 287500 62900 287800
rect 63200 287500 63400 287800
rect 63700 287500 63900 287800
rect 64200 287500 64400 287800
rect 64700 287500 64900 287800
rect 65200 287500 65400 287800
rect 65700 287500 65900 287800
rect 66200 287500 66400 287800
rect 66700 287500 66900 287800
rect 67200 287500 67400 287800
rect 67700 287500 67900 287800
rect 68200 287500 68400 287800
rect 68700 287500 68900 287800
rect 69200 287500 69400 287800
rect 69700 287500 69900 287800
rect 70200 287500 70400 287800
rect 70700 287500 70900 287800
rect 71200 287500 71400 287800
rect 71700 287500 71900 287800
rect 72200 287500 72400 287800
rect 72700 287500 72900 287800
rect 73200 287500 73400 287800
rect 73700 287500 74200 287800
rect 59200 287300 74200 287500
rect 59200 287000 59400 287300
rect 59700 287000 59900 287300
rect 60200 287000 60400 287300
rect 60700 287000 60900 287300
rect 61200 287000 61400 287300
rect 61700 287000 61900 287300
rect 62200 287000 62400 287300
rect 62700 287000 62900 287300
rect 63200 287000 63400 287300
rect 63700 287000 63900 287300
rect 64200 287000 64400 287300
rect 64700 287000 64900 287300
rect 65200 287000 65400 287300
rect 65700 287000 65900 287300
rect 66200 287000 66400 287300
rect 66700 287000 66900 287300
rect 67200 287000 67400 287300
rect 67700 287000 67900 287300
rect 68200 287000 68400 287300
rect 68700 287000 68900 287300
rect 69200 287000 69400 287300
rect 69700 287000 69900 287300
rect 70200 287000 70400 287300
rect 70700 287000 70900 287300
rect 71200 287000 71400 287300
rect 71700 287000 71900 287300
rect 72200 287000 72400 287300
rect 72700 287000 72900 287300
rect 73200 287000 73400 287300
rect 73700 287000 74200 287300
rect 59200 286800 74200 287000
rect 59200 286500 59400 286800
rect 59700 286500 59900 286800
rect 60200 286500 60400 286800
rect 60700 286500 60900 286800
rect 61200 286500 61400 286800
rect 61700 286500 61900 286800
rect 62200 286500 62400 286800
rect 62700 286500 62900 286800
rect 63200 286500 63400 286800
rect 63700 286500 63900 286800
rect 64200 286500 64400 286800
rect 64700 286500 64900 286800
rect 65200 286500 65400 286800
rect 65700 286500 65900 286800
rect 66200 286500 66400 286800
rect 66700 286500 66900 286800
rect 67200 286500 67400 286800
rect 67700 286500 67900 286800
rect 68200 286500 68400 286800
rect 68700 286500 68900 286800
rect 69200 286500 69400 286800
rect 69700 286500 69900 286800
rect 70200 286500 70400 286800
rect 70700 286500 70900 286800
rect 71200 286500 71400 286800
rect 71700 286500 71900 286800
rect 72200 286500 72400 286800
rect 72700 286500 72900 286800
rect 73200 286500 73400 286800
rect 73700 286500 74200 286800
rect 59200 286300 74200 286500
rect 59200 286000 59400 286300
rect 59700 286000 59900 286300
rect 60200 286000 60400 286300
rect 60700 286000 60900 286300
rect 61200 286000 61400 286300
rect 61700 286000 61900 286300
rect 62200 286000 62400 286300
rect 62700 286000 62900 286300
rect 63200 286000 63400 286300
rect 63700 286000 63900 286300
rect 64200 286000 64400 286300
rect 64700 286000 64900 286300
rect 65200 286000 65400 286300
rect 65700 286000 65900 286300
rect 66200 286000 66400 286300
rect 66700 286000 66900 286300
rect 67200 286000 67400 286300
rect 67700 286000 67900 286300
rect 68200 286000 68400 286300
rect 68700 286000 68900 286300
rect 69200 286000 69400 286300
rect 69700 286000 69900 286300
rect 70200 286000 70400 286300
rect 70700 286000 70900 286300
rect 71200 286000 71400 286300
rect 71700 286000 71900 286300
rect 72200 286000 72400 286300
rect 72700 286000 72900 286300
rect 73200 286000 73400 286300
rect 73700 286000 74200 286300
rect 21950 278550 22590 278580
rect 21950 278310 21980 278550
rect 22220 278310 22320 278550
rect 22560 278310 22590 278550
rect 21950 278190 22590 278310
rect 21950 277950 21980 278190
rect 22220 277950 22320 278190
rect 22560 277950 22590 278190
rect 12830 275470 13160 275510
rect 12830 275220 12870 275470
rect 13120 275220 13160 275470
rect 21950 275460 22590 277950
rect 33800 278400 35300 279300
rect 33800 278100 34000 278400
rect 34300 278100 34400 278400
rect 34700 278100 34800 278400
rect 35100 278100 35300 278400
rect 33800 276140 35300 278100
rect 33800 275900 34460 276140
rect 34700 275900 35300 276140
rect 12830 273570 13160 275220
rect 12830 273360 12870 273570
rect 12310 273330 12870 273360
rect 12310 273060 12360 273330
rect 12630 273320 12870 273330
rect 13120 273360 13160 273570
rect 14490 274130 14810 274170
rect 14490 273870 14520 274130
rect 14780 273870 14810 274130
rect 14490 273360 14810 273870
rect 16040 274130 16360 274170
rect 16040 273870 16070 274130
rect 16330 273870 16360 274130
rect 16040 273570 16360 273870
rect 15580 273540 16360 273570
rect 15580 273360 15610 273540
rect 13120 273330 15610 273360
rect 13120 273320 14000 273330
rect 12630 273060 14000 273320
rect 14270 273280 15610 273330
rect 15870 273280 16360 273540
rect 14270 273060 16360 273280
rect 12310 272870 16360 273060
rect 21290 274070 23140 275460
rect 21290 273820 22850 274070
rect 23100 273820 23140 274070
rect 21290 273810 23140 273820
rect 21290 273560 21330 273810
rect 21580 273560 23140 273810
rect 21290 272880 23140 273560
rect 23980 273550 24620 273850
rect 23980 273310 24320 273550
rect 24560 273310 24620 273550
rect 23980 273030 24620 273310
rect 21290 272870 23600 272880
rect 12310 272610 14520 272870
rect 14780 272610 16070 272870
rect 16330 272610 16360 272870
rect 12310 272280 16360 272610
rect 18670 272780 23600 272870
rect 18670 272520 18710 272780
rect 18970 272520 20230 272780
rect 20490 272530 21750 272780
rect 22000 272530 23280 272780
rect 23530 272530 23600 272780
rect 20490 272520 23600 272530
rect 18670 272440 23600 272520
rect 23980 272790 24320 273030
rect 24560 272790 24620 273030
rect 23980 272510 24620 272790
rect 18670 272430 23140 272440
rect 12310 272010 12360 272280
rect 12630 272010 14000 272280
rect 14270 272040 16360 272280
rect 14270 272010 15610 272040
rect 12310 271990 15610 272010
rect 12310 271980 12870 271990
rect 12830 271740 12870 271980
rect 13120 271980 15610 271990
rect 13120 271740 13160 271980
rect 12830 270090 13160 271740
rect 14490 271600 14810 271980
rect 15580 271780 15610 271980
rect 15870 271780 16360 272040
rect 15580 271750 16360 271780
rect 14490 271340 14520 271600
rect 14780 271340 14810 271600
rect 14490 271190 14810 271340
rect 16040 271600 16360 271750
rect 16040 271340 16070 271600
rect 16330 271340 16360 271600
rect 16040 271300 16360 271340
rect 21290 271750 23140 272430
rect 21290 271500 21330 271750
rect 21580 271500 23140 271750
rect 21290 271490 23140 271500
rect 23980 272270 24320 272510
rect 24560 272270 24620 272510
rect 23980 271990 24620 272270
rect 23980 271750 24320 271990
rect 24560 271750 24620 271990
rect 23980 271490 24620 271750
rect 33800 273010 35300 275900
rect 33800 272770 33980 273010
rect 34220 272770 34460 273010
rect 34700 272770 34940 273010
rect 35180 272770 35300 273010
rect 33800 272450 35300 272770
rect 33800 272210 33980 272450
rect 34220 272210 34460 272450
rect 34700 272210 34940 272450
rect 35180 272210 35300 272450
rect 21290 271240 22850 271490
rect 23100 271240 23140 271490
rect 12830 269840 12860 270090
rect 13110 269840 13160 270090
rect 12830 269810 13160 269840
rect 21290 269820 23140 271240
rect 21950 267300 22590 269820
rect 21950 267060 21980 267300
rect 22220 267060 22320 267300
rect 22560 267060 22590 267300
rect 21950 266940 22590 267060
rect 21950 266700 21980 266940
rect 22220 266700 22320 266940
rect 22560 266700 22590 266940
rect 21950 266670 22590 266700
rect 33800 269440 35300 272210
rect 33800 269200 34460 269440
rect 34700 269200 35300 269440
rect 33800 268600 35300 269200
rect 33800 268300 34000 268600
rect 34300 268300 34800 268600
rect 35100 268300 35300 268600
rect 33800 268100 35300 268300
rect 33800 267800 34000 268100
rect 34300 267800 34800 268100
rect 35100 267800 35300 268100
rect 33800 267600 35300 267800
rect 33800 267300 34000 267600
rect 34300 267300 34800 267600
rect 35100 267300 35300 267600
rect 33800 267100 35300 267300
rect 33800 266800 34000 267100
rect 34300 266800 34800 267100
rect 35100 266800 35300 267100
rect 33800 266600 35300 266800
rect 33800 266300 34000 266600
rect 34300 266300 34800 266600
rect 35100 266300 35300 266600
rect 33800 266100 35300 266300
rect 33800 265800 34000 266100
rect 34300 265800 34800 266100
rect 35100 265800 35300 266100
rect 33800 265600 35300 265800
rect 33800 265300 34000 265600
rect 34300 265300 34800 265600
rect 35100 265300 35300 265600
rect 33800 265100 35300 265300
rect 33800 264800 34000 265100
rect 34300 264800 34800 265100
rect 35100 264800 35300 265100
rect 33800 264600 35300 264800
rect 33800 264300 34000 264600
rect 34300 264300 34800 264600
rect 35100 264300 35300 264600
rect 33800 264100 35300 264300
rect 33800 263800 34000 264100
rect 34300 263800 34800 264100
rect 35100 263800 35300 264100
rect 33800 263600 35300 263800
rect 33800 263300 34000 263600
rect 34300 263300 34800 263600
rect 35100 263300 35300 263600
rect 33800 263100 35300 263300
rect 33800 262800 34000 263100
rect 34300 262800 34800 263100
rect 35100 262800 35300 263100
rect 33800 262600 35300 262800
rect 33800 262300 34000 262600
rect 34300 262300 34800 262600
rect 35100 262300 35300 262600
rect 33800 262100 35300 262300
rect 33800 261800 34000 262100
rect 34300 261800 34800 262100
rect 35100 261800 35300 262100
rect 33800 261600 35300 261800
rect 33800 261300 34000 261600
rect 34300 261300 34800 261600
rect 35100 261300 35300 261600
rect 33800 261100 35300 261300
rect 33800 260800 34000 261100
rect 34300 260800 34800 261100
rect 35100 260800 35300 261100
rect 33800 242000 35300 260800
rect 37100 276140 38500 276300
rect 37100 275900 37660 276140
rect 37900 275900 38500 276140
rect 37100 273010 38500 275900
rect 37100 272770 37180 273010
rect 37420 272770 37660 273010
rect 37900 272770 38140 273010
rect 38380 272770 38500 273010
rect 37100 272450 38500 272770
rect 37100 272210 37180 272450
rect 37420 272210 37660 272450
rect 37900 272210 38140 272450
rect 38380 272210 38500 272450
rect 37100 269440 38500 272210
rect 37100 269200 37660 269440
rect 37900 269200 38500 269440
rect 37100 268600 38500 269200
rect 37100 268300 37300 268600
rect 37600 268300 38000 268600
rect 38300 268300 38500 268600
rect 37100 268100 38500 268300
rect 37100 267800 37300 268100
rect 37600 267800 38000 268100
rect 38300 267800 38500 268100
rect 37100 267600 38500 267800
rect 37100 267300 37300 267600
rect 37600 267300 38000 267600
rect 38300 267300 38500 267600
rect 37100 267100 38500 267300
rect 37100 266800 37300 267100
rect 37600 266800 38000 267100
rect 38300 266800 38500 267100
rect 37100 266600 38500 266800
rect 37100 266300 37300 266600
rect 37600 266300 38000 266600
rect 38300 266300 38500 266600
rect 37100 266100 38500 266300
rect 37100 265800 37300 266100
rect 37600 265800 38000 266100
rect 38300 265800 38500 266100
rect 37100 265600 38500 265800
rect 37100 265300 37300 265600
rect 37600 265300 38000 265600
rect 38300 265300 38500 265600
rect 37100 265100 38500 265300
rect 37100 264800 37300 265100
rect 37600 264800 38000 265100
rect 38300 264800 38500 265100
rect 37100 264600 38500 264800
rect 37100 264300 37300 264600
rect 37600 264300 38000 264600
rect 38300 264300 38500 264600
rect 37100 264100 38500 264300
rect 37100 263800 37300 264100
rect 37600 263800 38000 264100
rect 38300 263800 38500 264100
rect 37100 263600 38500 263800
rect 37100 263300 37300 263600
rect 37600 263300 38000 263600
rect 38300 263300 38500 263600
rect 37100 263100 38500 263300
rect 37100 262800 37300 263100
rect 37600 262800 38000 263100
rect 38300 262800 38500 263100
rect 37100 262600 38500 262800
rect 37100 262300 37300 262600
rect 37600 262300 38000 262600
rect 38300 262300 38500 262600
rect 37100 262100 38500 262300
rect 37100 261800 37300 262100
rect 37600 261800 38000 262100
rect 38300 261800 38500 262100
rect 37100 261600 38500 261800
rect 37100 261300 37300 261600
rect 37600 261300 38000 261600
rect 38300 261300 38500 261600
rect 37100 261100 38500 261300
rect 37100 260800 37300 261100
rect 37600 260800 38000 261100
rect 38300 260800 38500 261100
rect 37100 260600 38500 260800
rect 40400 276140 41800 276300
rect 40400 275900 40980 276140
rect 41220 275900 41800 276140
rect 40400 273010 41800 275900
rect 40400 272770 40500 273010
rect 40740 272770 40980 273010
rect 41220 272770 41460 273010
rect 41700 272770 41800 273010
rect 40400 272450 41800 272770
rect 40400 272210 40500 272450
rect 40740 272210 40980 272450
rect 41220 272210 41460 272450
rect 41700 272210 41800 272450
rect 40400 269440 41800 272210
rect 40400 269200 40980 269440
rect 41220 269200 41800 269440
rect 40400 268600 41800 269200
rect 40400 268300 40600 268600
rect 40900 268300 41300 268600
rect 41600 268300 41800 268600
rect 40400 268100 41800 268300
rect 40400 267800 40600 268100
rect 40900 267800 41300 268100
rect 41600 267800 41800 268100
rect 40400 267600 41800 267800
rect 40400 267300 40600 267600
rect 40900 267300 41300 267600
rect 41600 267300 41800 267600
rect 40400 267100 41800 267300
rect 40400 266800 40600 267100
rect 40900 266800 41300 267100
rect 41600 266800 41800 267100
rect 40400 266600 41800 266800
rect 40400 266300 40600 266600
rect 40900 266300 41300 266600
rect 41600 266300 41800 266600
rect 40400 266100 41800 266300
rect 40400 265800 40600 266100
rect 40900 265800 41300 266100
rect 41600 265800 41800 266100
rect 40400 265600 41800 265800
rect 40400 265300 40600 265600
rect 40900 265300 41300 265600
rect 41600 265300 41800 265600
rect 40400 265100 41800 265300
rect 40400 264800 40600 265100
rect 40900 264800 41300 265100
rect 41600 264800 41800 265100
rect 40400 264600 41800 264800
rect 40400 264300 40600 264600
rect 40900 264300 41300 264600
rect 41600 264300 41800 264600
rect 40400 264100 41800 264300
rect 40400 263800 40600 264100
rect 40900 263800 41300 264100
rect 41600 263800 41800 264100
rect 40400 263600 41800 263800
rect 40400 263300 40600 263600
rect 40900 263300 41300 263600
rect 41600 263300 41800 263600
rect 40400 263100 41800 263300
rect 40400 262800 40600 263100
rect 40900 262800 41300 263100
rect 41600 262800 41800 263100
rect 40400 262600 41800 262800
rect 40400 262300 40600 262600
rect 40900 262300 41300 262600
rect 41600 262300 41800 262600
rect 40400 262100 41800 262300
rect 40400 261800 40600 262100
rect 40900 261800 41300 262100
rect 41600 261800 41800 262100
rect 40400 261600 41800 261800
rect 40400 261300 40600 261600
rect 40900 261300 41300 261600
rect 41600 261300 41800 261600
rect 40400 261100 41800 261300
rect 40400 260800 40600 261100
rect 40900 260800 41300 261100
rect 41600 260800 41800 261100
rect 40400 260600 41800 260800
rect 33800 241700 33900 242000
rect 34200 241700 34400 242000
rect 34700 241700 34900 242000
rect 35200 241700 35300 242000
rect 33800 241200 35300 241700
rect 33800 240900 33900 241200
rect 34200 240900 34400 241200
rect 34700 240900 34900 241200
rect 35200 240900 35300 241200
rect 33800 240800 35300 240900
rect 59200 252400 74200 286000
rect 59200 252100 59500 252400
rect 59800 252100 60100 252400
rect 60400 252100 60700 252400
rect 61000 252100 61400 252400
rect 61700 252100 62000 252400
rect 62300 252100 62600 252400
rect 62900 252100 63200 252400
rect 63500 252100 63800 252400
rect 64100 252100 64400 252400
rect 64700 252100 65100 252400
rect 65400 252100 65700 252400
rect 66000 252100 66300 252400
rect 66600 252100 66900 252400
rect 67200 252100 67500 252400
rect 67800 252100 68100 252400
rect 68400 252100 68700 252400
rect 69000 252100 69300 252400
rect 69600 252100 69900 252400
rect 70200 252100 70600 252400
rect 70900 252100 71300 252400
rect 71600 252100 72000 252400
rect 72300 252100 72800 252400
rect 73100 252100 73500 252400
rect 73800 252100 74200 252400
rect 59200 251700 74200 252100
rect 59200 251400 59500 251700
rect 59800 251400 60100 251700
rect 60400 251400 60700 251700
rect 61000 251400 61400 251700
rect 61700 251400 62000 251700
rect 62300 251400 62600 251700
rect 62900 251400 63200 251700
rect 63500 251400 63800 251700
rect 64100 251400 64400 251700
rect 64700 251400 65100 251700
rect 65400 251400 65700 251700
rect 66000 251400 66300 251700
rect 66600 251400 66900 251700
rect 67200 251400 67500 251700
rect 67800 251400 68100 251700
rect 68400 251400 68700 251700
rect 69000 251400 69300 251700
rect 69600 251400 69900 251700
rect 70200 251400 70600 251700
rect 70900 251400 71300 251700
rect 71600 251400 72000 251700
rect 72300 251400 72800 251700
rect 73100 251400 73500 251700
rect 73800 251400 74200 251700
rect 59200 218800 74200 251400
rect 59200 218400 60000 218800
rect 60400 218400 60800 218800
rect 61200 218400 61600 218800
rect 62000 218400 62400 218800
rect 62800 218400 63200 218800
rect 63600 218400 64000 218800
rect 64400 218400 69000 218800
rect 69400 218400 69800 218800
rect 70200 218400 70600 218800
rect 71000 218400 71400 218800
rect 71800 218400 72200 218800
rect 72600 218400 73000 218800
rect 73400 218400 74200 218800
rect 59200 218000 74200 218400
rect 59200 217600 60000 218000
rect 60400 217600 60800 218000
rect 61200 217600 61600 218000
rect 62000 217600 62400 218000
rect 62800 217600 63200 218000
rect 63600 217600 64000 218000
rect 64400 217600 69000 218000
rect 69400 217600 69800 218000
rect 70200 217600 70600 218000
rect 71000 217600 71400 218000
rect 71800 217600 72200 218000
rect 72600 217600 73000 218000
rect 73400 217600 74200 218000
rect 59200 217200 74200 217600
rect 59200 216800 60000 217200
rect 60400 216800 60800 217200
rect 61200 216800 61600 217200
rect 62000 216800 62400 217200
rect 62800 216800 63200 217200
rect 63600 216800 64000 217200
rect 64400 216800 69000 217200
rect 69400 216800 69800 217200
rect 70200 216800 70600 217200
rect 71000 216800 71400 217200
rect 71800 216800 72200 217200
rect 72600 216800 73000 217200
rect 73400 216800 74200 217200
rect 59200 216400 74200 216800
rect 59200 216000 60000 216400
rect 60400 216000 60800 216400
rect 61200 216000 61600 216400
rect 62000 216000 62400 216400
rect 62800 216000 63200 216400
rect 63600 216000 64000 216400
rect 64400 216000 69000 216400
rect 69400 216000 69800 216400
rect 70200 216000 70600 216400
rect 71000 216000 71400 216400
rect 71800 216000 72200 216400
rect 72600 216000 73000 216400
rect 73400 216000 74200 216400
rect 59200 215600 74200 216000
rect 59200 215200 60000 215600
rect 60400 215200 60800 215600
rect 61200 215200 61600 215600
rect 62000 215200 62400 215600
rect 62800 215200 63200 215600
rect 63600 215200 64000 215600
rect 64400 215200 69000 215600
rect 69400 215200 69800 215600
rect 70200 215200 70600 215600
rect 71000 215200 71400 215600
rect 71800 215200 72200 215600
rect 72600 215200 73000 215600
rect 73400 215200 74200 215600
rect 59200 214800 74200 215200
rect 59200 214400 60000 214800
rect 60400 214400 60800 214800
rect 61200 214400 61600 214800
rect 62000 214400 62400 214800
rect 62800 214400 63200 214800
rect 63600 214400 64000 214800
rect 64400 214400 69000 214800
rect 69400 214400 69800 214800
rect 70200 214400 70600 214800
rect 71000 214400 71400 214800
rect 71800 214400 72200 214800
rect 72600 214400 73000 214800
rect 73400 214400 74200 214800
rect 59200 210200 74200 214400
rect 59200 210000 69000 210200
rect 59200 209600 60000 210000
rect 60400 209600 60800 210000
rect 61200 209600 61600 210000
rect 62000 209600 62400 210000
rect 62800 209600 63200 210000
rect 63600 209600 64000 210000
rect 64400 209800 69000 210000
rect 69400 209800 69800 210200
rect 70200 209800 70600 210200
rect 71000 209800 71400 210200
rect 71800 209800 72200 210200
rect 72600 209800 73000 210200
rect 73400 209800 74200 210200
rect 64400 209600 74200 209800
rect 59200 209400 74200 209600
rect 59200 209200 69000 209400
rect 59200 208800 60000 209200
rect 60400 208800 60800 209200
rect 61200 208800 61600 209200
rect 62000 208800 62400 209200
rect 62800 208800 63200 209200
rect 63600 208800 64000 209200
rect 64400 209000 69000 209200
rect 69400 209000 69800 209400
rect 70200 209000 70600 209400
rect 71000 209000 71400 209400
rect 71800 209000 72200 209400
rect 72600 209000 73000 209400
rect 73400 209000 74200 209400
rect 64400 208800 74200 209000
rect 59200 208600 74200 208800
rect 59200 208400 69000 208600
rect 59200 208000 60000 208400
rect 60400 208000 60800 208400
rect 61200 208000 61600 208400
rect 62000 208000 62400 208400
rect 62800 208000 63200 208400
rect 63600 208000 64000 208400
rect 64400 208200 69000 208400
rect 69400 208200 69800 208600
rect 70200 208200 70600 208600
rect 71000 208200 71400 208600
rect 71800 208200 72200 208600
rect 72600 208200 73000 208600
rect 73400 208200 74200 208600
rect 64400 208000 74200 208200
rect 59200 207800 74200 208000
rect 59200 207600 69000 207800
rect 59200 207200 60000 207600
rect 60400 207200 60800 207600
rect 61200 207200 61600 207600
rect 62000 207200 62400 207600
rect 62800 207200 63200 207600
rect 63600 207200 64000 207600
rect 64400 207400 69000 207600
rect 69400 207400 69800 207800
rect 70200 207400 70600 207800
rect 71000 207400 71400 207800
rect 71800 207400 72200 207800
rect 72600 207400 73000 207800
rect 73400 207400 74200 207800
rect 64400 207200 74200 207400
rect 59200 207000 74200 207200
rect 59200 206800 69000 207000
rect 59200 206400 60000 206800
rect 60400 206400 60800 206800
rect 61200 206400 61600 206800
rect 62000 206400 62400 206800
rect 62800 206400 63200 206800
rect 63600 206400 64000 206800
rect 64400 206600 69000 206800
rect 69400 206600 69800 207000
rect 70200 206600 70600 207000
rect 71000 206600 71400 207000
rect 71800 206600 72200 207000
rect 72600 206600 73000 207000
rect 73400 206600 74200 207000
rect 64400 206400 74200 206600
rect 59200 206200 74200 206400
rect 59200 206000 69000 206200
rect 59200 205600 60000 206000
rect 60400 205600 60800 206000
rect 61200 205600 61600 206000
rect 62000 205600 62400 206000
rect 62800 205600 63200 206000
rect 63600 205600 64000 206000
rect 64400 205800 69000 206000
rect 69400 205800 69800 206200
rect 70200 205800 70600 206200
rect 71000 205800 71400 206200
rect 71800 205800 72200 206200
rect 72600 205800 73000 206200
rect 73400 205800 74200 206200
rect 64400 205600 74200 205800
rect 59200 204800 74200 205600
rect 283200 219400 292200 338500
rect 545700 288900 574640 289100
rect 545700 288600 545900 288900
rect 546200 288600 546400 288900
rect 546700 288600 546900 288900
rect 547200 288600 547400 288900
rect 547700 288600 547900 288900
rect 548200 288600 548400 288900
rect 548700 288600 569200 288900
rect 569500 288600 569800 288900
rect 570100 288700 574640 288900
rect 570100 288600 572800 288700
rect 545700 288400 572800 288600
rect 573100 288400 573300 288700
rect 573600 288400 573800 288700
rect 574100 288400 574300 288700
rect 574600 288400 574640 288700
rect 545700 288100 545900 288400
rect 546200 288100 546400 288400
rect 546700 288100 546900 288400
rect 547200 288100 547400 288400
rect 547700 288100 547900 288400
rect 548200 288100 548400 288400
rect 548700 288100 569200 288400
rect 569500 288100 569800 288400
rect 570100 288200 574640 288400
rect 570100 288100 572800 288200
rect 545700 287900 572800 288100
rect 573100 287900 573300 288200
rect 573600 287900 573800 288200
rect 574100 287900 574300 288200
rect 574600 287900 574640 288200
rect 545700 287600 545900 287900
rect 546200 287600 546400 287900
rect 546700 287600 546900 287900
rect 547200 287600 547400 287900
rect 547700 287600 547900 287900
rect 548200 287600 548400 287900
rect 548700 287600 569200 287900
rect 569500 287600 569800 287900
rect 570100 287600 574640 287900
rect 545700 287400 574640 287600
rect 283200 219000 285400 219400
rect 285800 219000 286200 219400
rect 286600 219000 287000 219400
rect 287400 219000 287800 219400
rect 288200 219000 288600 219400
rect 289000 219000 289400 219400
rect 289800 219000 292200 219400
rect 283200 218600 292200 219000
rect 283200 218200 285400 218600
rect 285800 218200 286200 218600
rect 286600 218200 287000 218600
rect 287400 218200 287800 218600
rect 288200 218200 288600 218600
rect 289000 218200 289400 218600
rect 289800 218200 292200 218600
rect 283200 217800 292200 218200
rect 283200 217400 285400 217800
rect 285800 217400 286200 217800
rect 286600 217400 287000 217800
rect 287400 217400 287800 217800
rect 288200 217400 288600 217800
rect 289000 217400 289400 217800
rect 289800 217400 292200 217800
rect 283200 217000 292200 217400
rect 283200 216600 285400 217000
rect 285800 216600 286200 217000
rect 286600 216600 287000 217000
rect 287400 216600 287800 217000
rect 288200 216600 288600 217000
rect 289000 216600 289400 217000
rect 289800 216600 292200 217000
rect 283200 216200 292200 216600
rect 283200 215800 285400 216200
rect 285800 215800 286200 216200
rect 286600 215800 287000 216200
rect 287400 215800 287800 216200
rect 288200 215800 288600 216200
rect 289000 215800 289400 216200
rect 289800 215800 292200 216200
rect 283200 215400 292200 215800
rect 283200 215000 285400 215400
rect 285800 215000 286200 215400
rect 286600 215000 287000 215400
rect 287400 215000 287800 215400
rect 288200 215000 288600 215400
rect 289000 215000 289400 215400
rect 289800 215000 292200 215400
rect 283200 214600 292200 215000
rect 283200 214200 285200 214600
rect 285600 214200 286000 214600
rect 286400 214200 286800 214600
rect 287200 214200 287600 214600
rect 288000 214200 288400 214600
rect 288800 214200 289200 214600
rect 289600 214200 292200 214600
rect 283200 213800 292200 214200
rect 283200 213400 285200 213800
rect 285600 213400 286000 213800
rect 286400 213400 286800 213800
rect 287200 213400 287600 213800
rect 288000 213400 288400 213800
rect 288800 213400 289200 213800
rect 289600 213400 292200 213800
rect 283200 213000 292200 213400
rect 283200 212600 285200 213000
rect 285600 212600 286000 213000
rect 286400 212600 286800 213000
rect 287200 212600 287600 213000
rect 288000 212600 288400 213000
rect 288800 212600 289200 213000
rect 289600 212600 292200 213000
rect 283200 212200 292200 212600
rect 283200 211800 285200 212200
rect 285600 211800 286000 212200
rect 286400 211800 286800 212200
rect 287200 211800 287600 212200
rect 288000 211800 288400 212200
rect 288800 211800 289200 212200
rect 289600 211800 292200 212200
rect 283200 211400 292200 211800
rect 283200 211000 285200 211400
rect 285600 211000 286000 211400
rect 286400 211000 286800 211400
rect 287200 211000 287600 211400
rect 288000 211000 288400 211400
rect 288800 211000 289200 211400
rect 289600 211000 292200 211400
rect 283200 210600 292200 211000
rect 283200 210200 285200 210600
rect 285600 210200 286000 210600
rect 286400 210200 286800 210600
rect 287200 210200 287600 210600
rect 288000 210200 288400 210600
rect 288800 210200 289200 210600
rect 289600 210200 292200 210600
rect 283200 209800 292200 210200
rect 283200 209400 285200 209800
rect 285600 209400 286000 209800
rect 286400 209400 286800 209800
rect 287200 209400 287600 209800
rect 288000 209400 288400 209800
rect 288800 209400 289200 209800
rect 289600 209400 292200 209800
rect 283200 209000 292200 209400
rect 283200 208600 285200 209000
rect 285600 208600 286000 209000
rect 286400 208600 286800 209000
rect 287200 208600 287600 209000
rect 288000 208600 288400 209000
rect 288800 208600 289200 209000
rect 289600 208600 292200 209000
rect 283200 208200 292200 208600
rect 283200 207800 285200 208200
rect 285600 207800 286000 208200
rect 286400 207800 286800 208200
rect 287200 207800 287600 208200
rect 288000 207800 288400 208200
rect 288800 207800 289200 208200
rect 289600 207800 292200 208200
rect 283200 207400 292200 207800
rect 283200 207000 285200 207400
rect 285600 207000 286000 207400
rect 286400 207000 286800 207400
rect 287200 207000 287600 207400
rect 288000 207000 288400 207400
rect 288800 207000 289200 207400
rect 289600 207000 292200 207400
rect 283200 206600 292200 207000
rect 283200 206200 285200 206600
rect 285600 206200 286000 206600
rect 286400 206200 286800 206600
rect 287200 206200 287600 206600
rect 288000 206200 288400 206600
rect 288800 206200 289200 206600
rect 289600 206200 292200 206600
rect 283200 205800 292200 206200
rect 283200 205400 285200 205800
rect 285600 205400 286000 205800
rect 286400 205400 286800 205800
rect 287200 205400 287600 205800
rect 288000 205400 288400 205800
rect 288800 205400 289200 205800
rect 289600 205400 292200 205800
rect 283200 204800 292200 205400
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use OTA_MULT_GM  OTA_MULT_GM_0
timestamp 1683391037
transform 1 0 544600 0 1 677936
box -10044 -14658 10212 17116
use OTA_fingers_031123_NON_FLAT  OTA_fingers_031123_NON_FLAT_0
timestamp 1683391037
transform 1 0 42740 0 1 684710
box -5940 -310 9780 16550
use analog_mux  analog_mux_0
timestamp 1684864136
transform 1 0 281327 0 1 350114
box -327 -10514 13727 4150
use constant_gm_fingers  constant_gm_fingers_0
timestamp 1683407140
transform 1 0 43810 0 1 682900
box -2700 -20100 4420 1140
use diode_connected_nmos  diode_connected_nmos_0
timestamp 1683391037
transform 1 0 23260 0 1 691860
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_1
timestamp 1683391037
transform 1 0 12860 0 1 691860
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_2
timestamp 1683391037
transform 1 0 75260 0 1 691860
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_3
timestamp 1683391037
transform 1 0 64860 0 1 691860
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_4
timestamp 1683391037
transform 1 0 563860 0 1 691660
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_5
timestamp 1683391037
transform 1 0 573060 0 1 691660
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_6
timestamp 1683391037
transform 0 1 572140 -1 0 684834
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_7
timestamp 1683391037
transform 0 1 572160 -1 0 677354
box -60 -60 1254 10360
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_0
timestamp 1683391037
transform 0 -1 37792 1 0 273375
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_1
timestamp 1683391037
transform 0 -1 37792 1 0 271835
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_2
timestamp 1683391037
transform 0 -1 37792 1 0 270285
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_3
timestamp 1683391037
transform 0 -1 37792 1 0 274925
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_4
timestamp 1683391037
transform 1 0 538336 0 1 274670
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_5
timestamp 1683391037
transform 1 0 539856 0 1 274670
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_6
timestamp 1683391037
transform 1 0 541366 0 1 274676
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_7
timestamp 1683391037
transform 1 0 542876 0 1 274676
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_0
timestamp 1683391037
transform 0 1 549214 -1 0 289928
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_1
timestamp 1683391037
transform 0 1 549214 -1 0 291398
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_2
timestamp 1683391037
transform 0 1 532154 -1 0 289928
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_3
timestamp 1683391037
transform 0 1 532154 -1 0 291398
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_4
timestamp 1683391037
transform 1 0 12444 0 1 278195
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_5
timestamp 1683391037
transform 1 0 13904 0 1 278195
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_6
timestamp 1683391037
transform 1 0 12444 0 1 267125
box -739 -1598 739 1598
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_7
timestamp 1683391037
transform 1 0 13904 0 1 267125
box -739 -1598 739 1598
<< labels >>
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 550 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 556 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 556 nsew signal bidirectional
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 704 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 703 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 701 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 700 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 707 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 706 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 705 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 53 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 54 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 55 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 56 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 58 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 59 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 60 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 61 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 62 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 63 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 64 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 65 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 66 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 67 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 68 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 69 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 70 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 71 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 72 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 73 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 74 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 75 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 76 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 77 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 78 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 79 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 80 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 81 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 82 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 83 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 85 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 86 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 87 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 88 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 89 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 90 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 91 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 92 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 93 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 94 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 95 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 96 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 97 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 98 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 99 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 100 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 101 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 102 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 103 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 104 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 105 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 106 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 107 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 108 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 109 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 110 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 112 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 113 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 114 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 115 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 116 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 117 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 118 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 119 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 120 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 121 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 122 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 123 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 124 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 125 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 126 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 127 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 128 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 129 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 130 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 131 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 132 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 133 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 134 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 135 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 136 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 137 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 139 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 140 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 141 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 142 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 143 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 144 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 145 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 146 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 147 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 148 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 149 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 150 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 151 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 152 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 153 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 154 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 155 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 156 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 157 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 158 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 159 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 160 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 161 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 162 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 163 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 164 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 165 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 166 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 167 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 168 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 169 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 170 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 171 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 172 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 173 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 174 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 175 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 176 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 177 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 178 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 179 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 180 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 181 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 182 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 183 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 184 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 185 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 186 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 187 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 188 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 189 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 190 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 191 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 192 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 193 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 194 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 195 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 196 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 197 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 198 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 199 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 200 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 201 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 202 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 203 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 204 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 205 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 206 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 207 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 208 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 209 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 210 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 211 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 212 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 213 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 214 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 215 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 216 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 217 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 218 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 219 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 220 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 221 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 222 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 223 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 224 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 225 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 226 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 227 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 228 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 229 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 230 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 231 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 232 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 233 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 234 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 235 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 236 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 237 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 238 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 239 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 240 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 241 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 242 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 243 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 244 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 245 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 246 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 247 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 248 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 249 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 250 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 251 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 252 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 253 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 254 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 255 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 256 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 257 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 258 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 259 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 260 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 261 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 262 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 263 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 264 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 265 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 266 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 267 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 268 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 269 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 270 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 271 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 272 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 273 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 274 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 275 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 276 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 277 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 278 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 279 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 280 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 281 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 282 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 283 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 284 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 285 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 286 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 287 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 288 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 289 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 290 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 291 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 292 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 293 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 294 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 295 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 296 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 297 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 298 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 299 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 300 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 301 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 302 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 303 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 304 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 305 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 306 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 307 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 308 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 309 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 310 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 311 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 312 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 313 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 314 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 315 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 316 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 317 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 318 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 319 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 320 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 321 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 322 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 323 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 324 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 325 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 326 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 327 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 328 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 329 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 330 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 331 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 332 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 333 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 334 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 335 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 336 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 337 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 338 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 339 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 340 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 341 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 342 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 343 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 344 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 345 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 346 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 347 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 348 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 349 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 350 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 351 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 352 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 353 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 354 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 355 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 356 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 357 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 358 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 359 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 360 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 361 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 362 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 363 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 364 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 365 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 366 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 367 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 368 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 369 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 370 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 371 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 372 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 373 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 374 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 375 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 376 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 377 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 378 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 379 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 380 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 381 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 382 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 383 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 384 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 385 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 386 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 387 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 388 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 389 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 390 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 391 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 392 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 393 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 394 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 395 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 396 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 397 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 398 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 399 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 400 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 401 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 402 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 403 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 404 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 405 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 406 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 407 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 408 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 409 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 410 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 411 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 412 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 413 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 414 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 415 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 416 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 417 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 418 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 419 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 420 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 421 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 422 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 423 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 424 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 425 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 426 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 427 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 428 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 429 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 430 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 431 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 432 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 433 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 434 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 435 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 436 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 437 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 438 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 439 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 440 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 441 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 442 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 443 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 444 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 445 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 446 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 447 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 448 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 449 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 450 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 451 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 452 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 453 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 454 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 455 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 456 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 457 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 458 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 459 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 460 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 461 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 462 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 463 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 464 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 465 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 466 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 467 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 468 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 469 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 470 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 471 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 472 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 473 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 474 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 475 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 476 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 477 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 478 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 479 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 480 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 481 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 482 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 483 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 484 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 485 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 486 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 487 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 488 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 489 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 490 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 491 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 492 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 493 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 494 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 495 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 496 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 497 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 498 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 499 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 500 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 501 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 502 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 503 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 504 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 505 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 506 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 507 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 508 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 509 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 510 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 511 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 512 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 513 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 514 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 515 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 516 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 517 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 518 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 519 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 520 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 521 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 522 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 523 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 524 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 525 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 526 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 527 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 528 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 529 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 530 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 531 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 532 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 533 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 534 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 535 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 536 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 537 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 538 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 539 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 540 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 541 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 542 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 543 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 544 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 545 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 546 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 547 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 548 nsew signal tristate
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 551 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 551 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 552 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 552 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 553 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 553 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 555 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 555 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 557 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 558 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 559 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 560 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 561 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 562 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 563 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 564 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 565 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 566 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 567 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 568 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 569 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 570 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 571 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 572 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 573 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 574 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 575 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 576 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 577 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 578 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 579 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 580 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 581 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 582 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 583 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 584 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 585 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 586 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 587 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 588 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 589 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 590 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 591 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 592 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 593 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 594 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 595 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 596 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 597 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 598 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 599 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 600 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 601 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 602 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 603 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 604 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 605 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 606 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 607 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 608 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 609 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 610 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 611 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 612 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 613 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 614 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 615 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 616 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 617 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 618 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 619 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 620 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 621 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 622 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 623 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 624 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 625 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 626 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 627 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 628 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 629 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 630 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 631 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 632 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 633 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 634 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 635 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 636 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 637 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 638 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 639 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 640 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 641 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 642 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 643 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 644 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 645 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 646 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 647 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 648 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 649 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 650 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 651 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 652 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 653 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 654 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 655 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 656 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 657 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 658 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 659 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 660 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 661 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 662 nsew signal input
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 554 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 554 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 553 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 553 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 551 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 551 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 550 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 549 nsew signal bidirectional
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 549 nsew signal bidirectional
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 138 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 111 nsew signal tristate
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 84 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 57 nsew signal input
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 52 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 51 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 50 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 49 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 48 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 47 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
