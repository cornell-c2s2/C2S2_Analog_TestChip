magic
tech sky130A
magscale 1 2
timestamp 1683929354
<< nwell >>
rect 1500 -990 1620 -970
rect 1820 -990 1940 -970
rect 2120 -990 2240 -970
rect 2440 -990 2560 -970
rect 2760 -990 2880 -970
<< locali >>
rect 1200 -990 1280 -930
rect 1520 -990 1600 -930
rect 1840 -990 1920 -930
rect 2140 -990 2220 -930
rect 2460 -990 2540 -930
rect 2780 -990 2860 -930
<< viali >>
rect 1200 -1070 1280 -990
rect 1520 -1070 1600 -990
rect 1840 -1070 1920 -990
rect 2140 -1070 2220 -990
rect 2460 -1070 2540 -990
rect 2780 -1070 2860 -990
<< metal1 >>
rect 970 260 3096 320
rect 970 -800 1030 260
rect 1100 -50 1110 160
rect 1170 -50 1180 160
rect 1290 -50 1300 160
rect 1360 -50 1370 160
rect 1480 -50 1490 160
rect 1550 -50 1560 160
rect 1670 -50 1680 160
rect 1740 -50 1750 160
rect 1870 -50 1880 160
rect 1940 -50 1950 160
rect 2060 -50 2070 160
rect 2130 -50 2140 160
rect 2250 -50 2260 160
rect 2320 -50 2330 160
rect 2440 -50 2450 160
rect 2510 -50 2520 160
rect 2630 -50 2640 160
rect 2700 -50 2710 160
rect 2820 -50 2830 160
rect 2890 -50 2900 160
rect 1190 -720 1200 -510
rect 1260 -720 1270 -510
rect 1380 -720 1390 -510
rect 1450 -720 1460 -510
rect 1580 -720 1590 -510
rect 1650 -720 1660 -510
rect 1770 -720 1780 -510
rect 1840 -720 1850 -510
rect 1960 -720 1970 -510
rect 2030 -720 2040 -510
rect 2150 -720 2160 -510
rect 2220 -720 2230 -510
rect 2340 -720 2350 -510
rect 2410 -720 2420 -510
rect 2540 -720 2550 -510
rect 2610 -720 2620 -510
rect 2730 -720 2740 -510
rect 2800 -720 2810 -510
rect 2920 -720 2930 -510
rect 2990 -720 3000 -510
rect 3036 -800 3096 260
rect 970 -860 3096 -800
rect 3210 260 4390 320
rect 3210 -800 3270 260
rect 3340 -40 3350 170
rect 3410 -40 3420 170
rect 3530 -40 3540 170
rect 3600 -40 3610 170
rect 3720 -40 3730 170
rect 3790 -40 3800 170
rect 3910 -40 3920 170
rect 3980 -40 3990 170
rect 4110 -40 4120 170
rect 4180 -40 4190 170
rect 3430 -730 3440 -520
rect 3500 -730 3510 -520
rect 3620 -730 3630 -520
rect 3690 -730 3700 -520
rect 3820 -740 3830 -530
rect 3890 -740 3900 -530
rect 4010 -740 4020 -530
rect 4080 -740 4090 -530
rect 4200 -740 4210 -530
rect 4270 -740 4280 -530
rect 4330 -800 4390 260
rect 3210 -860 4390 -800
rect 1188 -990 1292 -984
rect 1188 -1070 1200 -990
rect 1280 -1070 1292 -990
rect 1188 -1076 1292 -1070
rect 1508 -990 1612 -984
rect 1508 -1070 1520 -990
rect 1600 -1070 1612 -990
rect 1508 -1076 1612 -1070
rect 1828 -990 1932 -984
rect 1828 -1070 1840 -990
rect 1920 -1070 1932 -990
rect 1828 -1076 1932 -1070
rect 2128 -990 2232 -984
rect 2128 -1070 2140 -990
rect 2220 -1070 2232 -990
rect 2128 -1076 2232 -1070
rect 2448 -990 2552 -984
rect 2448 -1070 2460 -990
rect 2540 -1070 2552 -990
rect 2448 -1076 2552 -1070
rect 2768 -990 2872 -984
rect 2768 -1070 2780 -990
rect 2860 -1070 2872 -990
rect 2768 -1076 2872 -1070
<< via1 >>
rect 1110 -50 1170 160
rect 1300 -50 1360 160
rect 1490 -50 1550 160
rect 1680 -50 1740 160
rect 1880 -50 1940 160
rect 2070 -50 2130 160
rect 2260 -50 2320 160
rect 2450 -50 2510 160
rect 2640 -50 2700 160
rect 2830 -50 2890 160
rect 1200 -720 1260 -510
rect 1390 -720 1450 -510
rect 1590 -720 1650 -510
rect 1780 -720 1840 -510
rect 1970 -720 2030 -510
rect 2160 -720 2220 -510
rect 2350 -720 2410 -510
rect 2550 -720 2610 -510
rect 2740 -720 2800 -510
rect 2930 -720 2990 -510
rect 3350 -40 3410 170
rect 3540 -40 3600 170
rect 3730 -40 3790 170
rect 3920 -40 3980 170
rect 4120 -40 4180 170
rect 3440 -730 3500 -520
rect 3630 -730 3690 -520
rect 3830 -740 3890 -530
rect 4020 -740 4080 -530
rect 4210 -740 4270 -530
rect 1200 -1070 1280 -990
rect 1520 -1070 1600 -990
rect 1840 -1070 1920 -990
rect 2140 -1070 2220 -990
rect 2460 -1070 2540 -990
rect 2780 -1070 2860 -990
<< metal2 >>
rect 920 170 4438 184
rect 920 160 3350 170
rect 920 -50 1110 160
rect 1170 -50 1300 160
rect 1360 -50 1490 160
rect 1550 -50 1680 160
rect 1740 -50 1880 160
rect 1940 -50 2070 160
rect 2130 -50 2260 160
rect 2320 -50 2450 160
rect 2510 -50 2640 160
rect 2700 -50 2830 160
rect 2890 -40 3350 160
rect 3410 -40 3540 170
rect 3600 -40 3730 170
rect 3790 -40 3920 170
rect 3980 -40 4120 170
rect 4180 -40 4438 170
rect 2890 -50 4438 -40
rect 920 -70 4438 -50
rect 930 -490 4438 -488
rect 920 -510 4438 -490
rect 920 -720 1200 -510
rect 1260 -720 1390 -510
rect 1450 -720 1590 -510
rect 1650 -720 1780 -510
rect 1840 -720 1970 -510
rect 2030 -720 2160 -510
rect 2220 -720 2350 -510
rect 2410 -720 2550 -510
rect 2610 -720 2740 -510
rect 2800 -720 2930 -510
rect 2990 -520 4438 -510
rect 2990 -720 3440 -520
rect 920 -730 3440 -720
rect 3500 -730 3630 -520
rect 3690 -530 4438 -520
rect 3690 -730 3830 -530
rect 920 -740 3830 -730
rect 3890 -740 4020 -530
rect 4080 -740 4210 -530
rect 4270 -740 4438 -530
rect 930 -742 4438 -740
rect 3830 -750 3890 -742
rect 4020 -750 4080 -742
rect 4210 -750 4270 -742
rect 1200 -990 1280 -980
rect 1200 -1080 1280 -1070
rect 1520 -990 1600 -980
rect 1520 -1080 1600 -1070
rect 1840 -990 1920 -980
rect 1840 -1080 1920 -1070
rect 2140 -990 2220 -980
rect 2140 -1080 2220 -1070
rect 2460 -990 2540 -980
rect 2460 -1080 2540 -1070
rect 2780 -990 2860 -980
rect 2780 -1080 2860 -1070
<< via2 >>
rect 1200 -1070 1280 -990
rect 1520 -1070 1600 -990
rect 1840 -1070 1920 -990
rect 2140 -1070 2220 -990
rect 2460 -1070 2540 -990
rect 2780 -1070 2860 -990
<< metal3 >>
rect 1140 -990 3060 -970
rect 1140 -1070 1200 -990
rect 1280 -1070 1520 -990
rect 1600 -1070 1840 -990
rect 1920 -1070 2140 -990
rect 2220 -1070 2460 -990
rect 2540 -1070 2780 -990
rect 2860 -1070 3060 -990
rect 1140 -1090 3060 -1070
use sky130_fd_pr__pfet_01v8_BDZ9JN  XM1
timestamp 1683919673
transform 1 0 2049 0 1 -271
box -1079 -719 1079 719
use sky130_fd_pr__nfet_01v8_KBNS5F  sky130_fd_pr__nfet_01v8_KBNS5F_0
timestamp 1683919673
transform 1 0 3809 0 1 -270
box -599 -710 599 710
<< end >>
