magic
tech sky130A
magscale 1 2
timestamp 1676063568
<< xpolycontact >>
rect -573 23000 573 23432
rect -573 -23432 573 -23000
<< xpolyres >>
rect -573 -23000 573 23000
<< viali >>
rect -557 23017 557 23414
rect -557 -23414 557 -23017
<< metal1 >>
rect -569 23414 569 23420
rect -569 23017 -557 23414
rect 557 23017 569 23414
rect -569 23011 569 23017
rect -569 -23017 569 -23011
rect -569 -23414 -557 -23017
rect 557 -23414 569 -23017
rect -569 -23420 569 -23414
<< res5p73 >>
rect -575 -23002 575 23002
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 230 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 80.344k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
