magic
tech sky130A
magscale 1 2
timestamp 1683908447
<< pwell >>
rect 541314 677258 547888 678108
rect 541312 663278 547884 664522
<< metal1 >>
rect 65040 702260 65940 702300
rect 23380 702180 24340 702200
rect 23380 702060 23400 702180
rect 23520 702060 23600 702180
rect 23720 702060 23800 702180
rect 23920 702060 24000 702180
rect 24120 702060 24200 702180
rect 24320 702060 24340 702180
rect 23380 702040 24340 702060
rect 65040 702080 65060 702260
rect 65240 702080 65400 702260
rect 65580 702080 65740 702260
rect 65920 702080 65940 702260
rect 573240 702240 574140 702280
rect 65040 702040 65940 702080
rect 563800 702120 565120 702160
rect 563800 702020 563840 702120
rect 563940 702020 563980 702120
rect 564080 702020 564120 702120
rect 564220 702020 564260 702120
rect 564360 702020 564400 702120
rect 564500 702020 564540 702120
rect 564640 702020 564680 702120
rect 564780 702020 564820 702120
rect 564920 702020 564960 702120
rect 565060 702020 565120 702120
rect 563800 701980 565120 702020
rect 563800 701880 563840 701980
rect 563940 701880 563980 701980
rect 564080 701880 564120 701980
rect 564220 701880 564260 701980
rect 564360 701880 564400 701980
rect 564500 701880 564540 701980
rect 564640 701880 564680 701980
rect 564780 701880 564820 701980
rect 564920 701880 564960 701980
rect 565060 701880 565120 701980
rect 563800 701840 565120 701880
rect 573240 702140 573280 702240
rect 573380 702140 573420 702240
rect 573520 702140 573560 702240
rect 573660 702140 573700 702240
rect 573800 702140 573840 702240
rect 573940 702140 573980 702240
rect 574080 702140 574140 702240
rect 573240 701980 574140 702140
rect 573240 701880 573280 701980
rect 573380 701880 573420 701980
rect 573520 701880 573560 701980
rect 573660 701880 573700 701980
rect 573800 701880 573840 701980
rect 573940 701880 573980 701980
rect 574080 701880 574140 701980
rect 573240 701840 574140 701880
rect 565040 699740 573080 700240
rect 24440 693020 24600 693060
rect 24440 692900 24460 693020
rect 24580 692900 24600 693020
rect 24440 692840 24600 692900
rect 24440 692720 24460 692840
rect 24580 692720 24600 692840
rect 24440 692660 24600 692720
rect 24440 692540 24460 692660
rect 24580 692540 24600 692660
rect 64680 693000 64880 693040
rect 64680 692860 64720 693000
rect 64860 692860 64880 693000
rect 64680 692800 64880 692860
rect 64680 692660 64720 692800
rect 64860 692660 64880 692800
rect 64680 692620 64880 692660
rect 66040 693000 66240 693040
rect 66040 692860 66060 693000
rect 66200 692860 66240 693000
rect 66040 692800 66240 692860
rect 66040 692660 66060 692800
rect 66200 692660 66240 692800
rect 66040 692620 66240 692660
rect 75080 693000 75280 693040
rect 75080 692860 75120 693000
rect 75260 692860 75280 693000
rect 75080 692800 75280 692860
rect 75080 692660 75120 692800
rect 75260 692660 75280 692800
rect 75080 692620 75280 692660
rect 24440 692480 24600 692540
rect 24440 692360 24460 692480
rect 24580 692360 24600 692480
rect 24440 692300 24600 692360
rect 24440 692180 24460 692300
rect 24580 692180 24600 692300
rect 12800 691900 14120 691980
rect 12800 691700 12900 691900
rect 13100 691700 13200 691900
rect 13400 691700 13500 691900
rect 13700 691700 13800 691900
rect 14000 691700 14120 691900
rect 75220 691820 76500 691980
rect 12800 691600 14120 691700
rect 566260 691100 571840 691320
rect 566260 690900 566300 691100
rect 566500 690900 566700 691100
rect 566900 690900 567100 691100
rect 567300 690900 567500 691100
rect 567700 690900 567900 691100
rect 568100 690900 568300 691100
rect 568500 690900 568700 691100
rect 568900 690900 569100 691100
rect 569300 690900 569500 691100
rect 569700 690900 569900 691100
rect 570100 690900 570300 691100
rect 570500 690900 570700 691100
rect 570900 690900 571100 691100
rect 571300 690900 571500 691100
rect 571700 690900 571840 691100
rect 566260 690700 571840 690900
rect 566260 690500 566300 690700
rect 566500 690500 566700 690700
rect 566900 690500 567100 690700
rect 567300 690500 567500 690700
rect 567700 690500 567900 690700
rect 568100 690500 568300 690700
rect 568500 690500 568700 690700
rect 568900 690500 569100 690700
rect 569300 690500 569500 690700
rect 569700 690500 569900 690700
rect 570100 690500 570300 690700
rect 570500 690500 570700 690700
rect 570900 690500 571100 690700
rect 571300 690500 571500 690700
rect 571700 690500 571840 690700
rect 47100 690300 47400 690400
rect 47100 690200 47200 690300
rect 47300 690200 47400 690300
rect 47100 690010 47400 690200
rect 43870 689830 43950 690010
rect 45350 690000 47400 690010
rect 45350 689830 47200 690000
rect 47100 689800 47200 689830
rect 47300 689800 47400 690000
rect 47100 689600 47400 689800
rect 47100 689500 47200 689600
rect 47300 689500 47400 689600
rect 47100 689400 47400 689500
rect 566260 690300 571840 690500
rect 566260 690100 566300 690300
rect 566500 690100 566700 690300
rect 566900 690100 567100 690300
rect 567300 690100 567500 690300
rect 567700 690100 567900 690300
rect 568100 690100 568300 690300
rect 568500 690100 568700 690300
rect 568900 690100 569100 690300
rect 569300 690100 569500 690300
rect 569700 690100 569900 690300
rect 570100 690100 570300 690300
rect 570500 690100 570700 690300
rect 570900 690100 571100 690300
rect 571300 690100 571500 690300
rect 571700 690100 571840 690300
rect 566260 689900 571840 690100
rect 566260 689700 566300 689900
rect 566500 689700 566700 689900
rect 566900 689700 567100 689900
rect 567300 689700 567500 689900
rect 567700 689700 567900 689900
rect 568100 689700 568300 689900
rect 568500 689700 568700 689900
rect 568900 689700 569100 689900
rect 569300 689700 569500 689900
rect 569700 689700 569900 689900
rect 570100 689700 570300 689900
rect 570500 689700 570700 689900
rect 570900 689700 571100 689900
rect 571300 689700 571500 689900
rect 571700 689700 571840 689900
rect 566260 689520 571840 689700
rect 566260 689500 571820 689520
rect 566260 689300 566300 689500
rect 566500 689300 566700 689500
rect 566900 689300 567100 689500
rect 567300 689300 567500 689500
rect 567700 689300 567900 689500
rect 568100 689300 568300 689500
rect 568500 689300 568700 689500
rect 568900 689300 569100 689500
rect 569300 689300 569500 689500
rect 569700 689300 569900 689500
rect 570100 689300 570300 689500
rect 570500 689300 570700 689500
rect 570900 689300 571100 689500
rect 571300 689300 571500 689500
rect 571700 689300 571820 689500
rect 41900 688700 42200 688800
rect 41900 688600 42000 688700
rect 42100 688600 42200 688700
rect 41900 688500 42200 688600
rect 41900 688300 42000 688500
rect 42100 688490 42200 688500
rect 42100 688310 43870 688490
rect 42100 688300 42200 688310
rect 41900 688200 42200 688300
rect 41900 688100 42000 688200
rect 42100 688100 42200 688200
rect 41900 688000 42200 688100
rect 566260 685080 571820 689300
rect 548820 684860 571820 685080
rect 582320 684600 582660 684660
rect 548820 684360 554960 684580
rect 554420 682300 554960 684360
rect 582320 684520 582360 684600
rect 582440 684520 582540 684600
rect 582620 684520 582660 684600
rect 582320 684440 582660 684520
rect 582320 684360 582360 684440
rect 582440 684360 582540 684440
rect 582620 684360 582660 684440
rect 582320 684280 582660 684360
rect 582320 684200 582360 684280
rect 582440 684200 582540 684280
rect 582620 684200 582660 684280
rect 582320 684100 582660 684200
rect 582320 684020 582360 684100
rect 582440 684020 582540 684100
rect 582620 684020 582660 684100
rect 582320 683940 582660 684020
rect 582320 683860 582360 683940
rect 582440 683860 582540 683940
rect 582620 683860 582660 683940
rect 582320 683740 582660 683860
rect 554420 682200 563740 682300
rect 554420 682000 561700 682200
rect 561900 682000 562100 682200
rect 562300 682000 562500 682200
rect 562700 682000 562900 682200
rect 563100 682000 563300 682200
rect 563500 682000 563740 682200
rect 554420 681800 563740 682000
rect 554420 681600 561700 681800
rect 561900 681600 562100 681800
rect 562300 681600 562500 681800
rect 562700 681600 562900 681800
rect 563100 681600 563300 681800
rect 563500 681600 563740 681800
rect 554420 681400 563740 681600
rect 554420 681200 561700 681400
rect 561900 681200 562100 681400
rect 562300 681200 562500 681400
rect 562700 681200 562900 681400
rect 563100 681200 563300 681400
rect 563500 681200 563740 681400
rect 554420 681000 563740 681200
rect 554420 680800 561700 681000
rect 561900 680800 562100 681000
rect 562300 680800 562500 681000
rect 562700 680800 562900 681000
rect 563100 680800 563300 681000
rect 563500 680800 563740 681000
rect 554420 680600 563740 680800
rect 554420 680400 561700 680600
rect 561900 680400 562100 680600
rect 562300 680400 562500 680600
rect 562700 680400 562900 680600
rect 563100 680400 563300 680600
rect 563500 680400 563740 680600
rect 554420 680200 563740 680400
rect 554420 680000 561700 680200
rect 561900 680000 562100 680200
rect 562300 680000 562500 680200
rect 562700 680000 562900 680200
rect 563100 680000 563300 680200
rect 563500 680000 563740 680200
rect 554420 679800 563740 680000
rect 554420 679600 561700 679800
rect 561900 679600 562100 679800
rect 562300 679600 562500 679800
rect 562700 679600 562900 679800
rect 563100 679600 563300 679800
rect 563500 679600 563740 679800
rect 554420 679400 563740 679600
rect 554420 679200 561700 679400
rect 561900 679200 562100 679400
rect 562300 679200 562500 679400
rect 562700 679200 562900 679400
rect 563100 679200 563300 679400
rect 563500 679200 563740 679400
rect 554420 679000 563740 679200
rect 554420 678800 561700 679000
rect 561900 678800 562100 679000
rect 562300 678800 562500 679000
rect 562700 678800 562900 679000
rect 563100 678800 563300 679000
rect 563500 678800 563740 679000
rect 554420 678600 563740 678800
rect 554420 678400 561700 678600
rect 561900 678400 562100 678600
rect 562300 678400 562500 678600
rect 562700 678400 562900 678600
rect 563100 678400 563300 678600
rect 563500 678400 563740 678600
rect 554420 678340 563740 678400
rect 571800 677350 572390 683650
rect 571800 677300 572280 677350
rect 571800 677100 571900 677300
rect 572100 677100 572280 677300
rect 571800 677000 572280 677100
rect 571800 676800 571900 677000
rect 572100 676800 572280 677000
rect 571800 676700 572280 676800
rect 571800 676500 571900 676700
rect 572100 676500 572280 676700
rect 571800 676400 572280 676500
rect 571800 676200 571900 676400
rect 572100 676200 572280 676400
rect 571800 676100 572280 676200
rect 32600 663300 48300 663400
rect 32600 663000 32800 663300
rect 33100 663000 33300 663300
rect 33600 663000 33800 663300
rect 34100 663000 34300 663300
rect 34600 663000 34800 663300
rect 35100 663000 35300 663300
rect 35600 663000 35800 663300
rect 36100 663000 36300 663300
rect 36600 663000 36800 663300
rect 37100 663000 37300 663300
rect 37600 663000 37800 663300
rect 38100 663000 38300 663300
rect 38600 663000 38800 663300
rect 39100 663000 39300 663300
rect 39600 663000 39800 663300
rect 40100 663000 40300 663300
rect 40600 663000 48300 663300
rect 32600 662800 48300 663000
<< via1 >>
rect 23400 702060 23520 702180
rect 23600 702060 23720 702180
rect 23800 702060 23920 702180
rect 24000 702060 24120 702180
rect 24200 702060 24320 702180
rect 65060 702080 65240 702260
rect 65400 702080 65580 702260
rect 65740 702080 65920 702260
rect 563840 702020 563940 702120
rect 563980 702020 564080 702120
rect 564120 702020 564220 702120
rect 564260 702020 564360 702120
rect 564400 702020 564500 702120
rect 564540 702020 564640 702120
rect 564680 702020 564780 702120
rect 564820 702020 564920 702120
rect 564960 702020 565060 702120
rect 563840 701880 563940 701980
rect 563980 701880 564080 701980
rect 564120 701880 564220 701980
rect 564260 701880 564360 701980
rect 564400 701880 564500 701980
rect 564540 701880 564640 701980
rect 564680 701880 564780 701980
rect 564820 701880 564920 701980
rect 564960 701880 565060 701980
rect 573280 702140 573380 702240
rect 573420 702140 573520 702240
rect 573560 702140 573660 702240
rect 573700 702140 573800 702240
rect 573840 702140 573940 702240
rect 573980 702140 574080 702240
rect 573280 701880 573380 701980
rect 573420 701880 573520 701980
rect 573560 701880 573660 701980
rect 573700 701880 573800 701980
rect 573840 701880 573940 701980
rect 573980 701880 574080 701980
rect 24460 692900 24580 693020
rect 24460 692720 24580 692840
rect 24460 692540 24580 692660
rect 64720 692860 64860 693000
rect 64720 692660 64860 692800
rect 66060 692860 66200 693000
rect 66060 692660 66200 692800
rect 75120 692860 75260 693000
rect 75120 692660 75260 692800
rect 24460 692360 24580 692480
rect 24460 692180 24580 692300
rect 12900 691700 13100 691900
rect 13200 691700 13400 691900
rect 13500 691700 13700 691900
rect 13800 691700 14000 691900
rect 566300 690900 566500 691100
rect 566700 690900 566900 691100
rect 567100 690900 567300 691100
rect 567500 690900 567700 691100
rect 567900 690900 568100 691100
rect 568300 690900 568500 691100
rect 568700 690900 568900 691100
rect 569100 690900 569300 691100
rect 569500 690900 569700 691100
rect 569900 690900 570100 691100
rect 570300 690900 570500 691100
rect 570700 690900 570900 691100
rect 571100 690900 571300 691100
rect 571500 690900 571700 691100
rect 566300 690500 566500 690700
rect 566700 690500 566900 690700
rect 567100 690500 567300 690700
rect 567500 690500 567700 690700
rect 567900 690500 568100 690700
rect 568300 690500 568500 690700
rect 568700 690500 568900 690700
rect 569100 690500 569300 690700
rect 569500 690500 569700 690700
rect 569900 690500 570100 690700
rect 570300 690500 570500 690700
rect 570700 690500 570900 690700
rect 571100 690500 571300 690700
rect 571500 690500 571700 690700
rect 47200 690200 47300 690300
rect 47200 689800 47300 690000
rect 47200 689500 47300 689600
rect 566300 690100 566500 690300
rect 566700 690100 566900 690300
rect 567100 690100 567300 690300
rect 567500 690100 567700 690300
rect 567900 690100 568100 690300
rect 568300 690100 568500 690300
rect 568700 690100 568900 690300
rect 569100 690100 569300 690300
rect 569500 690100 569700 690300
rect 569900 690100 570100 690300
rect 570300 690100 570500 690300
rect 570700 690100 570900 690300
rect 571100 690100 571300 690300
rect 571500 690100 571700 690300
rect 566300 689700 566500 689900
rect 566700 689700 566900 689900
rect 567100 689700 567300 689900
rect 567500 689700 567700 689900
rect 567900 689700 568100 689900
rect 568300 689700 568500 689900
rect 568700 689700 568900 689900
rect 569100 689700 569300 689900
rect 569500 689700 569700 689900
rect 569900 689700 570100 689900
rect 570300 689700 570500 689900
rect 570700 689700 570900 689900
rect 571100 689700 571300 689900
rect 571500 689700 571700 689900
rect 566300 689300 566500 689500
rect 566700 689300 566900 689500
rect 567100 689300 567300 689500
rect 567500 689300 567700 689500
rect 567900 689300 568100 689500
rect 568300 689300 568500 689500
rect 568700 689300 568900 689500
rect 569100 689300 569300 689500
rect 569500 689300 569700 689500
rect 569900 689300 570100 689500
rect 570300 689300 570500 689500
rect 570700 689300 570900 689500
rect 571100 689300 571300 689500
rect 571500 689300 571700 689500
rect 42000 688600 42100 688700
rect 42000 688300 42100 688500
rect 42000 688100 42100 688200
rect 582360 684520 582440 684600
rect 582540 684520 582620 684600
rect 582360 684360 582440 684440
rect 582540 684360 582620 684440
rect 582360 684200 582440 684280
rect 582540 684200 582620 684280
rect 582360 684020 582440 684100
rect 582540 684020 582620 684100
rect 582360 683860 582440 683940
rect 582540 683860 582620 683940
rect 561700 682000 561900 682200
rect 562100 682000 562300 682200
rect 562500 682000 562700 682200
rect 562900 682000 563100 682200
rect 563300 682000 563500 682200
rect 561700 681600 561900 681800
rect 562100 681600 562300 681800
rect 562500 681600 562700 681800
rect 562900 681600 563100 681800
rect 563300 681600 563500 681800
rect 561700 681200 561900 681400
rect 562100 681200 562300 681400
rect 562500 681200 562700 681400
rect 562900 681200 563100 681400
rect 563300 681200 563500 681400
rect 561700 680800 561900 681000
rect 562100 680800 562300 681000
rect 562500 680800 562700 681000
rect 562900 680800 563100 681000
rect 563300 680800 563500 681000
rect 561700 680400 561900 680600
rect 562100 680400 562300 680600
rect 562500 680400 562700 680600
rect 562900 680400 563100 680600
rect 563300 680400 563500 680600
rect 561700 680000 561900 680200
rect 562100 680000 562300 680200
rect 562500 680000 562700 680200
rect 562900 680000 563100 680200
rect 563300 680000 563500 680200
rect 561700 679600 561900 679800
rect 562100 679600 562300 679800
rect 562500 679600 562700 679800
rect 562900 679600 563100 679800
rect 563300 679600 563500 679800
rect 561700 679200 561900 679400
rect 562100 679200 562300 679400
rect 562500 679200 562700 679400
rect 562900 679200 563100 679400
rect 563300 679200 563500 679400
rect 561700 678800 561900 679000
rect 562100 678800 562300 679000
rect 562500 678800 562700 679000
rect 562900 678800 563100 679000
rect 563300 678800 563500 679000
rect 561700 678400 561900 678600
rect 562100 678400 562300 678600
rect 562500 678400 562700 678600
rect 562900 678400 563100 678600
rect 563300 678400 563500 678600
rect 571900 677100 572100 677300
rect 571900 676800 572100 677000
rect 571900 676500 572100 676700
rect 571900 676200 572100 676400
rect 32800 663000 33100 663300
rect 33300 663000 33600 663300
rect 33800 663000 34100 663300
rect 34300 663000 34600 663300
rect 34800 663000 35100 663300
rect 35300 663000 35600 663300
rect 35800 663000 36100 663300
rect 36300 663000 36600 663300
rect 36800 663000 37100 663300
rect 37300 663000 37600 663300
rect 37800 663000 38100 663300
rect 38300 663000 38600 663300
rect 38800 663000 39100 663300
rect 39300 663000 39600 663300
rect 39800 663000 40100 663300
rect 40300 663000 40600 663300
<< metal2 >>
rect 65060 702260 65240 702270
rect 23400 702180 23520 702190
rect 23400 702050 23520 702060
rect 23600 702180 23720 702190
rect 23600 702050 23720 702060
rect 23800 702180 23920 702190
rect 23800 702050 23920 702060
rect 24000 702180 24120 702190
rect 24000 702050 24120 702060
rect 24200 702180 24320 702190
rect 65060 702070 65240 702080
rect 65400 702260 65580 702270
rect 65400 702070 65580 702080
rect 65740 702260 65920 702270
rect 573280 702240 573380 702250
rect 65740 702070 65920 702080
rect 563800 702120 565120 702160
rect 573280 702130 573380 702140
rect 573420 702240 573520 702250
rect 573420 702130 573520 702140
rect 573560 702240 573660 702250
rect 573560 702130 573660 702140
rect 573700 702240 573800 702250
rect 573700 702130 573800 702140
rect 573840 702240 573940 702250
rect 573840 702130 573940 702140
rect 573980 702240 574080 702250
rect 573980 702130 574080 702140
rect 24200 702050 24320 702060
rect 563800 702020 563840 702120
rect 563940 702020 563980 702120
rect 564080 702020 564120 702120
rect 564220 702020 564260 702120
rect 564360 702020 564400 702120
rect 564500 702020 564540 702120
rect 564640 702020 564680 702120
rect 564780 702020 564820 702120
rect 564920 702020 564960 702120
rect 565060 702020 565120 702120
rect 563800 701980 565120 702020
rect 563800 701880 563840 701980
rect 563940 701880 563980 701980
rect 564080 701880 564120 701980
rect 564220 701880 564260 701980
rect 564360 701880 564400 701980
rect 564500 701880 564540 701980
rect 564640 701880 564680 701980
rect 564780 701880 564820 701980
rect 564920 701880 564960 701980
rect 565060 701880 565120 701980
rect 563800 701840 565120 701880
rect 573280 701980 573380 701990
rect 573280 701870 573380 701880
rect 573420 701980 573520 701990
rect 573420 701870 573520 701880
rect 573560 701980 573660 701990
rect 573560 701870 573660 701880
rect 573700 701980 573800 701990
rect 573700 701870 573800 701880
rect 573840 701980 573940 701990
rect 573840 701870 573940 701880
rect 573980 701980 574080 701990
rect 573980 701870 574080 701880
rect 24460 693020 24580 693030
rect 24460 692890 24580 692900
rect 64720 693000 64860 693010
rect 64720 692850 64860 692860
rect 66060 693000 66200 693010
rect 66060 692850 66200 692860
rect 75120 693000 75260 693010
rect 75120 692850 75260 692860
rect 24460 692840 24580 692850
rect 24460 692710 24580 692720
rect 64720 692800 64860 692810
rect 24460 692660 24580 692670
rect 64720 692650 64860 692660
rect 66060 692800 66200 692810
rect 66060 692650 66200 692660
rect 75120 692800 75260 692810
rect 75120 692650 75260 692660
rect 24460 692530 24580 692540
rect 24460 692480 24580 692490
rect 24460 692350 24580 692360
rect 24460 692300 24580 692310
rect 24460 692170 24580 692180
rect 12900 691900 13100 691910
rect 12900 691690 13100 691700
rect 13200 691900 13400 691910
rect 13200 691690 13400 691700
rect 13500 691900 13700 691910
rect 13500 691690 13700 691700
rect 13800 691900 14000 691910
rect 13800 691690 14000 691700
rect 566290 690900 566300 691100
rect 566500 690900 566510 691100
rect 566690 690900 566700 691100
rect 566900 690900 566910 691100
rect 567090 690900 567100 691100
rect 567300 690900 567310 691100
rect 567490 690900 567500 691100
rect 567700 690900 567710 691100
rect 567890 690900 567900 691100
rect 568100 690900 568110 691100
rect 568290 690900 568300 691100
rect 568500 690900 568510 691100
rect 568690 690900 568700 691100
rect 568900 690900 568910 691100
rect 569090 690900 569100 691100
rect 569300 690900 569310 691100
rect 569490 690900 569500 691100
rect 569700 690900 569710 691100
rect 569890 690900 569900 691100
rect 570100 690900 570110 691100
rect 570290 690900 570300 691100
rect 570500 690900 570510 691100
rect 570690 690900 570700 691100
rect 570900 690900 570910 691100
rect 571090 690900 571100 691100
rect 571300 690900 571310 691100
rect 571490 690900 571500 691100
rect 571700 690900 571710 691100
rect 566290 690500 566300 690700
rect 566500 690500 566510 690700
rect 566690 690500 566700 690700
rect 566900 690500 566910 690700
rect 567090 690500 567100 690700
rect 567300 690500 567310 690700
rect 567490 690500 567500 690700
rect 567700 690500 567710 690700
rect 567890 690500 567900 690700
rect 568100 690500 568110 690700
rect 568290 690500 568300 690700
rect 568500 690500 568510 690700
rect 568690 690500 568700 690700
rect 568900 690500 568910 690700
rect 569090 690500 569100 690700
rect 569300 690500 569310 690700
rect 569490 690500 569500 690700
rect 569700 690500 569710 690700
rect 569890 690500 569900 690700
rect 570100 690500 570110 690700
rect 570290 690500 570300 690700
rect 570500 690500 570510 690700
rect 570690 690500 570700 690700
rect 570900 690500 570910 690700
rect 571090 690500 571100 690700
rect 571300 690500 571310 690700
rect 571490 690500 571500 690700
rect 571700 690500 571710 690700
rect 47200 690300 47300 690310
rect 47200 690190 47300 690200
rect 566290 690100 566300 690300
rect 566500 690100 566510 690300
rect 566690 690100 566700 690300
rect 566900 690100 566910 690300
rect 567090 690100 567100 690300
rect 567300 690100 567310 690300
rect 567490 690100 567500 690300
rect 567700 690100 567710 690300
rect 567890 690100 567900 690300
rect 568100 690100 568110 690300
rect 568290 690100 568300 690300
rect 568500 690100 568510 690300
rect 568690 690100 568700 690300
rect 568900 690100 568910 690300
rect 569090 690100 569100 690300
rect 569300 690100 569310 690300
rect 569490 690100 569500 690300
rect 569700 690100 569710 690300
rect 569890 690100 569900 690300
rect 570100 690100 570110 690300
rect 570290 690100 570300 690300
rect 570500 690100 570510 690300
rect 570690 690100 570700 690300
rect 570900 690100 570910 690300
rect 571090 690100 571100 690300
rect 571300 690100 571310 690300
rect 571490 690100 571500 690300
rect 571700 690100 571710 690300
rect 47200 690000 47300 690010
rect 47200 689790 47300 689800
rect 566290 689700 566300 689900
rect 566500 689700 566510 689900
rect 566690 689700 566700 689900
rect 566900 689700 566910 689900
rect 567090 689700 567100 689900
rect 567300 689700 567310 689900
rect 567490 689700 567500 689900
rect 567700 689700 567710 689900
rect 567890 689700 567900 689900
rect 568100 689700 568110 689900
rect 568290 689700 568300 689900
rect 568500 689700 568510 689900
rect 568690 689700 568700 689900
rect 568900 689700 568910 689900
rect 569090 689700 569100 689900
rect 569300 689700 569310 689900
rect 569490 689700 569500 689900
rect 569700 689700 569710 689900
rect 569890 689700 569900 689900
rect 570100 689700 570110 689900
rect 570290 689700 570300 689900
rect 570500 689700 570510 689900
rect 570690 689700 570700 689900
rect 570900 689700 570910 689900
rect 571090 689700 571100 689900
rect 571300 689700 571310 689900
rect 571490 689700 571500 689900
rect 571700 689700 571710 689900
rect 47200 689600 47300 689610
rect 47200 689490 47300 689500
rect 566290 689300 566300 689500
rect 566500 689300 566510 689500
rect 566690 689300 566700 689500
rect 566900 689300 566910 689500
rect 567090 689300 567100 689500
rect 567300 689300 567310 689500
rect 567490 689300 567500 689500
rect 567700 689300 567710 689500
rect 567890 689300 567900 689500
rect 568100 689300 568110 689500
rect 568290 689300 568300 689500
rect 568500 689300 568510 689500
rect 568690 689300 568700 689500
rect 568900 689300 568910 689500
rect 569090 689300 569100 689500
rect 569300 689300 569310 689500
rect 569490 689300 569500 689500
rect 569700 689300 569710 689500
rect 569890 689300 569900 689500
rect 570100 689300 570110 689500
rect 570290 689300 570300 689500
rect 570500 689300 570510 689500
rect 570690 689300 570700 689500
rect 570900 689300 570910 689500
rect 571090 689300 571100 689500
rect 571300 689300 571310 689500
rect 571490 689300 571500 689500
rect 571700 689300 571710 689500
rect 42000 688700 42100 688710
rect 42000 688590 42100 688600
rect 42000 688500 42100 688510
rect 42000 688290 42100 688300
rect 42000 688200 42100 688210
rect 42000 688090 42100 688100
rect 42240 683120 42640 684610
rect 42240 683040 42260 683120
rect 42340 683040 42400 683120
rect 42480 683040 42540 683120
rect 42620 683040 42640 683120
rect 42240 683020 42640 683040
rect 46640 683120 47040 684610
rect 582360 684600 582440 684610
rect 582360 684510 582440 684520
rect 582540 684600 582620 684610
rect 582540 684510 582620 684520
rect 582360 684440 582440 684450
rect 582360 684350 582440 684360
rect 582540 684440 582620 684450
rect 582540 684350 582620 684360
rect 582360 684280 582440 684290
rect 582360 684190 582440 684200
rect 582540 684280 582620 684290
rect 582540 684190 582620 684200
rect 582360 684100 582440 684110
rect 582360 684010 582440 684020
rect 582540 684100 582620 684110
rect 582540 684010 582620 684020
rect 582360 683940 582440 683950
rect 582360 683850 582440 683860
rect 582540 683940 582620 683950
rect 582540 683850 582620 683860
rect 46640 683040 46660 683120
rect 46740 683040 46800 683120
rect 46880 683040 46940 683120
rect 47020 683040 47040 683120
rect 46640 683020 47040 683040
rect 561700 682200 561900 682210
rect 561700 681990 561900 682000
rect 562100 682200 562300 682210
rect 562100 681990 562300 682000
rect 562500 682200 562700 682210
rect 562500 681990 562700 682000
rect 562900 682200 563100 682210
rect 562900 681990 563100 682000
rect 563300 682200 563500 682210
rect 563300 681990 563500 682000
rect 561700 681800 561900 681810
rect 561700 681590 561900 681600
rect 562100 681800 562300 681810
rect 562100 681590 562300 681600
rect 562500 681800 562700 681810
rect 562500 681590 562700 681600
rect 562900 681800 563100 681810
rect 562900 681590 563100 681600
rect 563300 681800 563500 681810
rect 563300 681590 563500 681600
rect 561700 681400 561900 681410
rect 561700 681190 561900 681200
rect 562100 681400 562300 681410
rect 562100 681190 562300 681200
rect 562500 681400 562700 681410
rect 562500 681190 562700 681200
rect 562900 681400 563100 681410
rect 562900 681190 563100 681200
rect 563300 681400 563500 681410
rect 563300 681190 563500 681200
rect 561700 681000 561900 681010
rect 561700 680790 561900 680800
rect 562100 681000 562300 681010
rect 562100 680790 562300 680800
rect 562500 681000 562700 681010
rect 562500 680790 562700 680800
rect 562900 681000 563100 681010
rect 562900 680790 563100 680800
rect 563300 681000 563500 681010
rect 563300 680790 563500 680800
rect 561700 680600 561900 680610
rect 561700 680390 561900 680400
rect 562100 680600 562300 680610
rect 562100 680390 562300 680400
rect 562500 680600 562700 680610
rect 562500 680390 562700 680400
rect 562900 680600 563100 680610
rect 562900 680390 563100 680400
rect 563300 680600 563500 680610
rect 563300 680390 563500 680400
rect 561700 680200 561900 680210
rect 561700 679990 561900 680000
rect 562100 680200 562300 680210
rect 562100 679990 562300 680000
rect 562500 680200 562700 680210
rect 562500 679990 562700 680000
rect 562900 680200 563100 680210
rect 562900 679990 563100 680000
rect 563300 680200 563500 680210
rect 563300 679990 563500 680000
rect 561700 679800 561900 679810
rect 561700 679590 561900 679600
rect 562100 679800 562300 679810
rect 562100 679590 562300 679600
rect 562500 679800 562700 679810
rect 562500 679590 562700 679600
rect 562900 679800 563100 679810
rect 562900 679590 563100 679600
rect 563300 679800 563500 679810
rect 563300 679590 563500 679600
rect 561700 679400 561900 679410
rect 561700 679190 561900 679200
rect 562100 679400 562300 679410
rect 562100 679190 562300 679200
rect 562500 679400 562700 679410
rect 562500 679190 562700 679200
rect 562900 679400 563100 679410
rect 562900 679190 563100 679200
rect 563300 679400 563500 679410
rect 563300 679190 563500 679200
rect 561700 679000 561900 679010
rect 561700 678790 561900 678800
rect 562100 679000 562300 679010
rect 562100 678790 562300 678800
rect 562500 679000 562700 679010
rect 562500 678790 562700 678800
rect 562900 679000 563100 679010
rect 562900 678790 563100 678800
rect 563300 679000 563500 679010
rect 563300 678790 563500 678800
rect 561700 678600 561900 678610
rect 561700 678390 561900 678400
rect 562100 678600 562300 678610
rect 562100 678390 562300 678400
rect 562500 678600 562700 678610
rect 562500 678390 562700 678400
rect 562900 678600 563100 678610
rect 562900 678390 563100 678400
rect 563300 678600 563500 678610
rect 563300 678390 563500 678400
rect 571900 677300 572100 677310
rect 571900 677090 572100 677100
rect 571900 677000 572100 677010
rect 571900 676790 572100 676800
rect 571900 676700 572100 676710
rect 571900 676490 572100 676500
rect 571900 676400 572100 676410
rect 571900 676190 572100 676200
rect 32800 663300 33100 663310
rect 32800 662990 33100 663000
rect 33300 663300 33600 663310
rect 33300 662990 33600 663000
rect 33800 663300 34100 663310
rect 33800 662990 34100 663000
rect 34300 663300 34600 663310
rect 34300 662990 34600 663000
rect 34800 663300 35100 663310
rect 34800 662990 35100 663000
rect 35300 663300 35600 663310
rect 35300 662990 35600 663000
rect 35800 663300 36100 663310
rect 35800 662990 36100 663000
rect 36300 663300 36600 663310
rect 36300 662990 36600 663000
rect 36800 663300 37100 663310
rect 36800 662990 37100 663000
rect 37300 663300 37600 663310
rect 37300 662990 37600 663000
rect 37800 663300 38100 663310
rect 37800 662990 38100 663000
rect 38300 663300 38600 663310
rect 38300 662990 38600 663000
rect 38800 663300 39100 663310
rect 38800 662990 39100 663000
rect 39300 663300 39600 663310
rect 39300 662990 39600 663000
rect 39800 663300 40100 663310
rect 39800 662990 40100 663000
rect 40300 663300 40600 663310
rect 40300 662990 40600 663000
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 23400 702060 23520 702180
rect 23600 702060 23720 702180
rect 23800 702060 23920 702180
rect 24000 702060 24120 702180
rect 24200 702060 24320 702180
rect 65060 702080 65240 702260
rect 65400 702080 65580 702260
rect 65740 702080 65920 702260
rect 573280 702140 573380 702240
rect 573420 702140 573520 702240
rect 573560 702140 573660 702240
rect 573700 702140 573800 702240
rect 573840 702140 573940 702240
rect 573980 702140 574080 702240
rect 563840 702020 563940 702120
rect 563980 702020 564080 702120
rect 564120 702020 564220 702120
rect 564260 702020 564360 702120
rect 564400 702020 564500 702120
rect 564540 702020 564640 702120
rect 564680 702020 564780 702120
rect 564820 702020 564920 702120
rect 564960 702020 565060 702120
rect 563840 701880 563940 701980
rect 563980 701880 564080 701980
rect 564120 701880 564220 701980
rect 564260 701880 564360 701980
rect 564400 701880 564500 701980
rect 564540 701880 564640 701980
rect 564680 701880 564780 701980
rect 564820 701880 564920 701980
rect 564960 701880 565060 701980
rect 573280 701880 573380 701980
rect 573420 701880 573520 701980
rect 573560 701880 573660 701980
rect 573700 701880 573800 701980
rect 573840 701880 573940 701980
rect 573980 701880 574080 701980
rect 24460 692900 24580 693020
rect 64720 692860 64860 693000
rect 66060 692860 66200 693000
rect 75120 692860 75260 693000
rect 24460 692720 24580 692840
rect 24460 692540 24580 692660
rect 64720 692660 64860 692800
rect 66060 692660 66200 692800
rect 75120 692660 75260 692800
rect 24460 692360 24580 692480
rect 24460 692180 24580 692300
rect 12900 691700 13100 691900
rect 13200 691700 13400 691900
rect 13500 691700 13700 691900
rect 13800 691700 14000 691900
rect 566300 690900 566500 691100
rect 566700 690900 566900 691100
rect 567100 690900 567300 691100
rect 567500 690900 567700 691100
rect 567900 690900 568100 691100
rect 568300 690900 568500 691100
rect 568700 690900 568900 691100
rect 569100 690900 569300 691100
rect 569500 690900 569700 691100
rect 569900 690900 570100 691100
rect 570300 690900 570500 691100
rect 570700 690900 570900 691100
rect 571100 690900 571300 691100
rect 571500 690900 571700 691100
rect 566300 690500 566500 690700
rect 566700 690500 566900 690700
rect 567100 690500 567300 690700
rect 567500 690500 567700 690700
rect 567900 690500 568100 690700
rect 568300 690500 568500 690700
rect 568700 690500 568900 690700
rect 569100 690500 569300 690700
rect 569500 690500 569700 690700
rect 569900 690500 570100 690700
rect 570300 690500 570500 690700
rect 570700 690500 570900 690700
rect 571100 690500 571300 690700
rect 571500 690500 571700 690700
rect 47200 690200 47300 690300
rect 566300 690100 566500 690300
rect 566700 690100 566900 690300
rect 567100 690100 567300 690300
rect 567500 690100 567700 690300
rect 567900 690100 568100 690300
rect 568300 690100 568500 690300
rect 568700 690100 568900 690300
rect 569100 690100 569300 690300
rect 569500 690100 569700 690300
rect 569900 690100 570100 690300
rect 570300 690100 570500 690300
rect 570700 690100 570900 690300
rect 571100 690100 571300 690300
rect 571500 690100 571700 690300
rect 47200 689800 47300 690000
rect 566300 689700 566500 689900
rect 566700 689700 566900 689900
rect 567100 689700 567300 689900
rect 567500 689700 567700 689900
rect 567900 689700 568100 689900
rect 568300 689700 568500 689900
rect 568700 689700 568900 689900
rect 569100 689700 569300 689900
rect 569500 689700 569700 689900
rect 569900 689700 570100 689900
rect 570300 689700 570500 689900
rect 570700 689700 570900 689900
rect 571100 689700 571300 689900
rect 571500 689700 571700 689900
rect 47200 689500 47300 689600
rect 566300 689300 566500 689500
rect 566700 689300 566900 689500
rect 567100 689300 567300 689500
rect 567500 689300 567700 689500
rect 567900 689300 568100 689500
rect 568300 689300 568500 689500
rect 568700 689300 568900 689500
rect 569100 689300 569300 689500
rect 569500 689300 569700 689500
rect 569900 689300 570100 689500
rect 570300 689300 570500 689500
rect 570700 689300 570900 689500
rect 571100 689300 571300 689500
rect 571500 689300 571700 689500
rect 42000 688600 42100 688700
rect 42000 688300 42100 688500
rect 42000 688100 42100 688200
rect 42260 683040 42340 683120
rect 42400 683040 42480 683120
rect 42540 683040 42620 683120
rect 582360 684520 582440 684600
rect 582540 684520 582620 684600
rect 582360 684360 582440 684440
rect 582540 684360 582620 684440
rect 582360 684200 582440 684280
rect 582540 684200 582620 684280
rect 582360 684020 582440 684100
rect 582540 684020 582620 684100
rect 582360 683860 582440 683940
rect 582540 683860 582620 683940
rect 46660 683040 46740 683120
rect 46800 683040 46880 683120
rect 46940 683040 47020 683120
rect 561700 682000 561900 682200
rect 562100 682000 562300 682200
rect 562500 682000 562700 682200
rect 562900 682000 563100 682200
rect 563300 682000 563500 682200
rect 561700 681600 561900 681800
rect 562100 681600 562300 681800
rect 562500 681600 562700 681800
rect 562900 681600 563100 681800
rect 563300 681600 563500 681800
rect 561700 681200 561900 681400
rect 562100 681200 562300 681400
rect 562500 681200 562700 681400
rect 562900 681200 563100 681400
rect 563300 681200 563500 681400
rect 561700 680800 561900 681000
rect 562100 680800 562300 681000
rect 562500 680800 562700 681000
rect 562900 680800 563100 681000
rect 563300 680800 563500 681000
rect 561700 680400 561900 680600
rect 562100 680400 562300 680600
rect 562500 680400 562700 680600
rect 562900 680400 563100 680600
rect 563300 680400 563500 680600
rect 561700 680000 561900 680200
rect 562100 680000 562300 680200
rect 562500 680000 562700 680200
rect 562900 680000 563100 680200
rect 563300 680000 563500 680200
rect 561700 679600 561900 679800
rect 562100 679600 562300 679800
rect 562500 679600 562700 679800
rect 562900 679600 563100 679800
rect 563300 679600 563500 679800
rect 561700 679200 561900 679400
rect 562100 679200 562300 679400
rect 562500 679200 562700 679400
rect 562900 679200 563100 679400
rect 563300 679200 563500 679400
rect 561700 678800 561900 679000
rect 562100 678800 562300 679000
rect 562500 678800 562700 679000
rect 562900 678800 563100 679000
rect 563300 678800 563500 679000
rect 561700 678400 561900 678600
rect 562100 678400 562300 678600
rect 562500 678400 562700 678600
rect 562900 678400 563100 678600
rect 563300 678400 563500 678600
rect 571900 677100 572100 677300
rect 571900 676800 572100 677000
rect 571900 676500 572100 676700
rect 571900 676200 572100 676400
rect 32800 663000 33100 663300
rect 33300 663000 33600 663300
rect 33800 663000 34100 663300
rect 34300 663000 34600 663300
rect 34800 663000 35100 663300
rect 35300 663000 35600 663300
rect 35800 663000 36100 663300
rect 36300 663000 36600 663300
rect 36800 663000 37100 663300
rect 37300 663000 37600 663300
rect 37800 663000 38100 663300
rect 38300 663000 38600 663300
rect 38800 663000 39100 663300
rect 39300 663000 39600 663300
rect 39800 663000 40100 663300
rect 40300 663000 40600 663300
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 703700 470394 704800
rect 510594 704000 515394 704800
rect 520594 704000 525394 704800
rect 566594 704000 571594 704800
rect 16200 702200 21200 702300
rect 16200 702000 16400 702200
rect 16600 702000 16800 702200
rect 17000 702000 17200 702200
rect 17400 702000 17600 702200
rect 17800 702000 18000 702200
rect 18200 702000 18400 702200
rect 18600 702000 18800 702200
rect 19000 702000 19200 702200
rect 19400 702000 19600 702200
rect 19800 702000 20000 702200
rect 20200 702000 20400 702200
rect 20600 702000 20800 702200
rect 21000 702000 21200 702200
rect 65050 702260 65250 702265
rect 23390 702180 23530 702185
rect 23390 702060 23400 702180
rect 23520 702060 23530 702180
rect 23390 702055 23530 702060
rect 23590 702180 23730 702185
rect 23590 702060 23600 702180
rect 23720 702060 23730 702180
rect 23590 702055 23730 702060
rect 23790 702180 23930 702185
rect 23790 702060 23800 702180
rect 23920 702060 23930 702180
rect 23790 702055 23930 702060
rect 23990 702180 24130 702185
rect 23990 702060 24000 702180
rect 24120 702060 24130 702180
rect 23990 702055 24130 702060
rect 24190 702180 24330 702185
rect 24190 702060 24200 702180
rect 24320 702060 24330 702180
rect 65050 702080 65060 702260
rect 65240 702080 65250 702260
rect 65050 702075 65250 702080
rect 65390 702260 65590 702265
rect 65390 702080 65400 702260
rect 65580 702080 65590 702260
rect 65390 702075 65590 702080
rect 65730 702260 65930 702265
rect 65730 702080 65740 702260
rect 65920 702080 65930 702260
rect 65730 702075 65930 702080
rect 68200 702200 73200 702300
rect 24190 702055 24330 702060
rect 16200 701800 21200 702000
rect 16200 701600 16400 701800
rect 16600 701600 16800 701800
rect 17000 701600 17200 701800
rect 17400 701600 17600 701800
rect 17800 701600 18000 701800
rect 18200 701600 18400 701800
rect 18600 701600 18800 701800
rect 19000 701600 19200 701800
rect 19400 701600 19600 701800
rect 19800 701600 20000 701800
rect 20200 701600 20400 701800
rect 20600 701600 20800 701800
rect 21000 701600 21200 701800
rect 16200 701400 21200 701600
rect 16200 701200 16400 701400
rect 16600 701200 16800 701400
rect 17000 701200 17200 701400
rect 17400 701200 17600 701400
rect 17800 701200 18000 701400
rect 18200 701200 18400 701400
rect 18600 701200 18800 701400
rect 19000 701200 19200 701400
rect 19400 701200 19600 701400
rect 19800 701200 20000 701400
rect 20200 701200 20400 701400
rect 20600 701200 20800 701400
rect 21000 701200 21200 701400
rect 16200 701000 21200 701200
rect 16200 700800 16400 701000
rect 16600 700800 16800 701000
rect 17000 700800 17200 701000
rect 17400 700800 17600 701000
rect 17800 700800 18000 701000
rect 18200 700800 18400 701000
rect 18600 700800 18800 701000
rect 19000 700800 19200 701000
rect 19400 700800 19600 701000
rect 19800 700800 20000 701000
rect 20200 700800 20400 701000
rect 20600 700800 20800 701000
rect 21000 700800 21200 701000
rect 16200 700600 21200 700800
rect 16200 700400 16400 700600
rect 16600 700400 16800 700600
rect 17000 700400 17200 700600
rect 17400 700400 17600 700600
rect 17800 700400 18000 700600
rect 18200 700400 18400 700600
rect 18600 700400 18800 700600
rect 19000 700400 19200 700600
rect 19400 700400 19600 700600
rect 19800 700400 20000 700600
rect 20200 700400 20400 700600
rect 20600 700400 20800 700600
rect 21000 700400 21200 700600
rect 16200 700200 21200 700400
rect 16200 700000 16400 700200
rect 16600 700000 16800 700200
rect 17000 700000 17200 700200
rect 17400 700000 17600 700200
rect 17800 700000 18000 700200
rect 18200 700000 18400 700200
rect 18600 700000 18800 700200
rect 19000 700000 19200 700200
rect 19400 700000 19600 700200
rect 19800 700000 20000 700200
rect 20200 700000 20400 700200
rect 20600 700000 20800 700200
rect 21000 700000 21200 700200
rect 16200 699800 21200 700000
rect 68200 702000 68400 702200
rect 68600 702000 68800 702200
rect 69000 702000 69200 702200
rect 69400 702000 69600 702200
rect 69800 702000 70000 702200
rect 70200 702000 70400 702200
rect 70600 702000 70800 702200
rect 71000 702000 71200 702200
rect 71400 702000 71600 702200
rect 71800 702000 72000 702200
rect 72200 702000 72400 702200
rect 72600 702000 72800 702200
rect 73000 702000 73200 702200
rect 68200 701800 73200 702000
rect 68200 701600 68400 701800
rect 68600 701600 68800 701800
rect 69000 701600 69200 701800
rect 69400 701600 69600 701800
rect 69800 701600 70000 701800
rect 70200 701600 70400 701800
rect 70600 701600 70800 701800
rect 71000 701600 71200 701800
rect 71400 701600 71600 701800
rect 71800 701600 72000 701800
rect 72200 701600 72400 701800
rect 72600 701600 72800 701800
rect 73000 701600 73200 701800
rect 68200 701400 73200 701600
rect 68200 701200 68400 701400
rect 68600 701200 68800 701400
rect 69000 701200 69200 701400
rect 69400 701200 69600 701400
rect 69800 701200 70000 701400
rect 70200 701200 70400 701400
rect 70600 701200 70800 701400
rect 71000 701200 71200 701400
rect 71400 701200 71600 701400
rect 71800 701200 72000 701400
rect 72200 701200 72400 701400
rect 72600 701200 72800 701400
rect 73000 701200 73200 701400
rect 68200 701000 73200 701200
rect 68200 700800 68400 701000
rect 68600 700800 68800 701000
rect 69000 700800 69200 701000
rect 69400 700800 69600 701000
rect 69800 700800 70000 701000
rect 70200 700800 70400 701000
rect 70600 700800 70800 701000
rect 71000 700800 71200 701000
rect 71400 700800 71600 701000
rect 71800 700800 72000 701000
rect 72200 700800 72400 701000
rect 72600 700800 72800 701000
rect 73000 700800 73200 701000
rect 68200 700600 73200 700800
rect 68200 700400 68400 700600
rect 68600 700400 68800 700600
rect 69000 700400 69200 700600
rect 69400 700400 69600 700600
rect 69800 700400 70000 700600
rect 70200 700400 70400 700600
rect 70600 700400 70800 700600
rect 71000 700400 71200 700600
rect 71400 700400 71600 700600
rect 71800 700400 72000 700600
rect 72200 700400 72400 700600
rect 72600 700400 72800 700600
rect 73000 700400 73200 700600
rect 68200 700200 73200 700400
rect 68200 700000 68400 700200
rect 68600 700000 68800 700200
rect 69000 700000 69200 700200
rect 69400 700000 69600 700200
rect 69800 700000 70000 700200
rect 70200 700000 70400 700200
rect 70600 700000 70800 700200
rect 71000 700000 71200 700200
rect 71400 700000 71600 700200
rect 71800 700000 72000 700200
rect 72200 700000 72400 700200
rect 72600 700000 72800 700200
rect 73000 700000 73200 700200
rect 68200 699800 73200 700000
rect 12990 698000 13000 698200
rect 13200 698000 13210 698200
rect 13590 698000 13600 698200
rect 13800 698000 13810 698200
rect 23390 698000 23400 698200
rect 23600 698000 23610 698200
rect 23790 698000 23800 698200
rect 24000 698000 24010 698200
rect 24190 698000 24200 698200
rect 24400 698000 24410 698200
rect 64990 698000 65000 698200
rect 65200 698000 65210 698200
rect 65590 698000 65600 698200
rect 65800 698000 65810 698200
rect 75390 698000 75400 698200
rect 75600 698000 75610 698200
rect 75990 698000 76000 698200
rect 76200 698000 76210 698200
rect 12990 697600 13000 697800
rect 13200 697600 13210 697800
rect 13590 697600 13600 697800
rect 13800 697600 13810 697800
rect 23390 697600 23400 697800
rect 23600 697600 23610 697800
rect 23790 697600 23800 697800
rect 24000 697600 24010 697800
rect 24190 697600 24200 697800
rect 24400 697600 24410 697800
rect 64990 697600 65000 697800
rect 65200 697600 65210 697800
rect 65590 697600 65600 697800
rect 65800 697600 65810 697800
rect 75390 697600 75400 697800
rect 75600 697600 75610 697800
rect 75990 697600 76000 697800
rect 76200 697600 76210 697800
rect 23390 697200 23400 697400
rect 23600 697200 23610 697400
rect 23790 697200 23800 697400
rect 24000 697200 24010 697400
rect 24190 697200 24200 697400
rect 24400 697200 24410 697400
rect 64990 697200 65000 697400
rect 65200 697200 65210 697400
rect 65590 697200 65600 697400
rect 65800 697200 65810 697400
rect 75390 697200 75400 697400
rect 75600 697200 75610 697400
rect 75990 697200 76000 697400
rect 76200 697200 76210 697400
rect 12990 697000 13000 697200
rect 13200 697000 13210 697200
rect 13590 697000 13600 697200
rect 13800 697000 13810 697200
rect 23390 696800 23400 697000
rect 23600 696800 23610 697000
rect 23790 696800 23800 697000
rect 24000 696800 24010 697000
rect 24190 696800 24200 697000
rect 24400 696800 24410 697000
rect 64990 696800 65000 697000
rect 65200 696800 65210 697000
rect 65590 696800 65600 697000
rect 65800 696800 65810 697000
rect 75390 696800 75400 697000
rect 75600 696800 75610 697000
rect 75990 696800 76000 697000
rect 76200 696800 76210 697000
rect 12990 696600 13000 696800
rect 13200 696600 13210 696800
rect 13590 696600 13600 696800
rect 13800 696600 13810 696800
rect 23300 696600 24400 696700
rect 23300 696400 23400 696600
rect 23600 696400 23800 696600
rect 24000 696400 24200 696600
rect 24400 696400 24410 696600
rect 64990 696400 65000 696600
rect 65200 696400 65210 696600
rect 65590 696400 65600 696600
rect 65800 696400 65810 696600
rect 75390 696400 75400 696600
rect 75600 696400 75610 696600
rect 75990 696400 76000 696600
rect 76200 696400 76210 696600
rect 24440 693020 39320 693060
rect 24440 692900 24460 693020
rect 24580 693000 39320 693020
rect 24580 692900 38700 693000
rect 24440 692840 38700 692900
rect 38860 692840 39120 693000
rect 39280 692840 39320 693000
rect 24440 692720 24460 692840
rect 24580 692780 39320 692840
rect 24580 692720 38700 692780
rect 24440 692660 38700 692720
rect 24440 692540 24460 692660
rect 24580 692620 38700 692660
rect 38860 692620 39120 692780
rect 39280 692620 39320 692780
rect 49920 693000 64880 693040
rect 49920 692860 49960 693000
rect 50100 692860 50180 693000
rect 50320 692860 50400 693000
rect 50540 692860 64720 693000
rect 64860 692860 64880 693000
rect 49920 692800 64880 692860
rect 49920 692660 49960 692800
rect 50100 692660 50180 692800
rect 50320 692660 50400 692800
rect 50540 692660 64720 692800
rect 64860 692660 64880 692800
rect 49920 692620 64880 692660
rect 66040 693000 75280 693040
rect 66040 692860 66060 693000
rect 66200 692860 75120 693000
rect 75260 692860 75280 693000
rect 66040 692800 75280 692860
rect 66040 692660 66060 692800
rect 66200 692660 75120 692800
rect 75260 692660 75280 692800
rect 66040 692620 75280 692660
rect 24580 692560 39320 692620
rect 24580 692540 38700 692560
rect 24440 692480 38700 692540
rect 24440 692360 24460 692480
rect 24580 692400 38700 692480
rect 38860 692400 39120 692560
rect 39280 692400 39320 692560
rect 24580 692360 39320 692400
rect 24440 692340 39320 692360
rect 24440 692300 38700 692340
rect 24440 692180 24460 692300
rect 24580 692180 38700 692300
rect 38860 692180 39120 692340
rect 39280 692180 39320 692340
rect 24440 692140 39320 692180
rect 12890 691900 13110 691905
rect 12890 691700 12900 691900
rect 13100 691700 13110 691900
rect 12890 691695 13110 691700
rect 13190 691900 13410 691905
rect 13190 691700 13200 691900
rect 13400 691700 13410 691900
rect 13190 691695 13410 691700
rect 13490 691900 13710 691905
rect 13490 691700 13500 691900
rect 13700 691700 13710 691900
rect 13490 691695 13710 691700
rect 13790 691900 14010 691905
rect 13790 691700 13800 691900
rect 14000 691700 14010 691900
rect 13790 691695 14010 691700
rect 46320 691900 62200 692040
rect 46320 691700 58000 691900
rect 58200 691700 58400 691900
rect 58600 691700 58800 691900
rect 59000 691700 59200 691900
rect 59400 691700 59600 691900
rect 59800 691700 60000 691900
rect 60200 691700 60400 691900
rect 60600 691700 60800 691900
rect 61000 691700 61200 691900
rect 61400 691700 61600 691900
rect 61800 691700 62200 691900
rect 46320 691560 62200 691700
rect 465100 690500 470600 703700
rect 510400 701600 525470 704000
rect 510400 701400 515700 701600
rect 515900 701400 516100 701600
rect 516300 701400 516500 701600
rect 516700 701400 516900 701600
rect 517100 701400 517300 701600
rect 517500 701400 517700 701600
rect 517900 701400 518100 701600
rect 518300 701400 518500 701600
rect 518700 701400 518900 701600
rect 519100 701400 519300 701600
rect 519500 701400 519700 701600
rect 519900 701400 520100 701600
rect 520300 701400 520500 701600
rect 520700 701400 525470 701600
rect 510400 701200 525470 701400
rect 510400 701000 515700 701200
rect 515900 701000 516100 701200
rect 516300 701000 516500 701200
rect 516700 701000 516900 701200
rect 517100 701000 517300 701200
rect 517500 701000 517700 701200
rect 517900 701000 518100 701200
rect 518300 701000 518500 701200
rect 518700 701000 518900 701200
rect 519100 701000 519300 701200
rect 519500 701000 519700 701200
rect 519900 701000 520100 701200
rect 520300 701000 520500 701200
rect 520700 701000 525470 701200
rect 510400 700800 525470 701000
rect 510400 700600 515700 700800
rect 515900 700600 516100 700800
rect 516300 700600 516500 700800
rect 516700 700600 516900 700800
rect 517100 700600 517300 700800
rect 517500 700600 517700 700800
rect 517900 700600 518100 700800
rect 518300 700600 518500 700800
rect 518700 700600 518900 700800
rect 519100 700600 519300 700800
rect 519500 700600 519700 700800
rect 519900 700600 520100 700800
rect 520300 700600 520500 700800
rect 520700 700600 525470 700800
rect 510400 700400 525470 700600
rect 510400 700200 515700 700400
rect 515900 700200 516100 700400
rect 516300 700200 516500 700400
rect 516700 700200 516900 700400
rect 517100 700200 517300 700400
rect 517500 700200 517700 700400
rect 517900 700200 518100 700400
rect 518300 700200 518500 700400
rect 518700 700200 518900 700400
rect 519100 700200 519300 700400
rect 519500 700200 519700 700400
rect 519900 700200 520100 700400
rect 520300 700200 520500 700400
rect 520700 700200 525470 700400
rect 510400 700000 525470 700200
rect 510400 699800 515700 700000
rect 515900 699800 516100 700000
rect 516300 699800 516500 700000
rect 516700 699800 516900 700000
rect 517100 699800 517300 700000
rect 517500 699800 517700 700000
rect 517900 699800 518100 700000
rect 518300 699800 518500 700000
rect 518700 699800 518900 700000
rect 519100 699800 519300 700000
rect 519500 699800 519700 700000
rect 519900 699800 520100 700000
rect 520300 699800 520500 700000
rect 520700 699800 525470 700000
rect 510400 699600 525470 699800
rect 510400 699400 515700 699600
rect 515900 699400 516100 699600
rect 516300 699400 516500 699600
rect 516700 699400 516900 699600
rect 517100 699400 517300 699600
rect 517500 699400 517700 699600
rect 517900 699400 518100 699600
rect 518300 699400 518500 699600
rect 518700 699400 518900 699600
rect 519100 699400 519300 699600
rect 519500 699400 519700 699600
rect 519900 699400 520100 699600
rect 520300 699400 520500 699600
rect 520700 699400 525470 699600
rect 510400 699200 525470 699400
rect 510400 699000 515700 699200
rect 515900 699000 516100 699200
rect 516300 699000 516500 699200
rect 516700 699000 516900 699200
rect 517100 699000 517300 699200
rect 517500 699000 517700 699200
rect 517900 699000 518100 699200
rect 518300 699000 518500 699200
rect 518700 699000 518900 699200
rect 519100 699000 519300 699200
rect 519500 699000 519700 699200
rect 519900 699000 520100 699200
rect 520300 699000 520500 699200
rect 520700 699000 525470 699200
rect 510400 698600 525470 699000
rect 560300 702120 565120 702400
rect 560300 702020 563840 702120
rect 563940 702020 563980 702120
rect 564080 702020 564120 702120
rect 564220 702020 564260 702120
rect 564360 702020 564400 702120
rect 564500 702020 564540 702120
rect 564640 702020 564680 702120
rect 564780 702020 564820 702120
rect 564920 702020 564960 702120
rect 565060 702020 565120 702120
rect 560300 701980 565120 702020
rect 560300 701880 563840 701980
rect 563940 701880 563980 701980
rect 564080 701880 564120 701980
rect 564220 701880 564260 701980
rect 564360 701880 564400 701980
rect 564500 701880 564540 701980
rect 564640 701880 564680 701980
rect 564780 701880 564820 701980
rect 564920 701880 564960 701980
rect 565060 701880 565120 701980
rect 560300 701800 565120 701880
rect 566200 702280 572000 704000
rect 566200 702240 574140 702280
rect 566200 702140 573280 702240
rect 573380 702140 573420 702240
rect 573520 702140 573560 702240
rect 573660 702140 573700 702240
rect 573800 702140 573840 702240
rect 573940 702140 573980 702240
rect 574080 702140 574140 702240
rect 566200 701980 574140 702140
rect 566200 701880 573280 701980
rect 573380 701880 573420 701980
rect 573520 701880 573560 701980
rect 573660 701880 573700 701980
rect 573800 701880 573840 701980
rect 573940 701880 573980 701980
rect 574080 701880 574140 701980
rect 566200 701840 574140 701880
rect 560300 697600 561600 701800
rect 566200 698160 572000 701840
rect 515500 697400 561600 697600
rect 515500 697200 515700 697400
rect 515900 697200 516100 697400
rect 516300 697200 516500 697400
rect 516700 697200 516900 697400
rect 517100 697200 517300 697400
rect 517500 697200 517700 697400
rect 517900 697200 518100 697400
rect 518300 697200 518500 697400
rect 518700 697200 518900 697400
rect 519100 697200 519300 697400
rect 519500 697200 519700 697400
rect 519900 697200 520100 697400
rect 520300 697200 520500 697400
rect 520700 697200 561600 697400
rect 515500 697000 561600 697200
rect 515500 696800 515700 697000
rect 515900 696800 516100 697000
rect 516300 696800 516500 697000
rect 516700 696800 516900 697000
rect 517100 696800 517300 697000
rect 517500 696800 517700 697000
rect 517900 696800 518100 697000
rect 518300 696800 518500 697000
rect 518700 696800 518900 697000
rect 519100 696800 519300 697000
rect 519500 696800 519700 697000
rect 519900 696800 520100 697000
rect 520300 696800 520500 697000
rect 520700 696800 561600 697000
rect 515500 696600 561600 696800
rect 515500 696400 515700 696600
rect 515900 696400 516100 696600
rect 516300 696400 516500 696600
rect 516700 696400 516900 696600
rect 517100 696400 517300 696600
rect 517500 696400 517700 696600
rect 517900 696400 518100 696600
rect 518300 696400 518500 696600
rect 518700 696400 518900 696600
rect 519100 696400 519300 696600
rect 519500 696400 519700 696600
rect 519900 696400 520100 696600
rect 520300 696400 520500 696600
rect 520700 696400 561600 696600
rect 515500 696000 561600 696400
rect 563800 696220 572000 698160
rect 566200 691100 572000 696220
rect 573100 698000 574220 698180
rect 573100 697800 573300 698000
rect 573500 697800 573800 698000
rect 574000 697800 574220 698000
rect 573100 697600 574220 697800
rect 573100 697400 573300 697600
rect 573500 697400 573800 697600
rect 574000 697400 574220 697600
rect 573100 697200 574220 697400
rect 573100 697000 573300 697200
rect 573500 697000 573800 697200
rect 574000 697000 574220 697200
rect 573100 696800 574220 697000
rect 573100 696600 573300 696800
rect 573500 696600 573800 696800
rect 574000 696600 574220 696800
rect 573100 696400 574220 696600
rect 573100 696200 573300 696400
rect 573500 696200 573800 696400
rect 574000 696200 574220 696400
rect 573100 696100 574220 696200
rect 566200 690900 566300 691100
rect 566500 690900 566700 691100
rect 566900 690900 567100 691100
rect 567300 690900 567500 691100
rect 567700 690900 567900 691100
rect 568100 690900 568300 691100
rect 568500 690900 568700 691100
rect 568900 690900 569100 691100
rect 569300 690900 569500 691100
rect 569700 690900 569900 691100
rect 570100 690900 570300 691100
rect 570500 690900 570700 691100
rect 570900 690900 571100 691100
rect 571300 690900 571500 691100
rect 571700 690900 572000 691100
rect 566200 690700 572000 690900
rect 566200 690500 566300 690700
rect 566500 690500 566700 690700
rect 566900 690500 567100 690700
rect 567300 690500 567500 690700
rect 567700 690500 567900 690700
rect 568100 690500 568300 690700
rect 568500 690500 568700 690700
rect 568900 690500 569100 690700
rect 569300 690500 569500 690700
rect 569700 690500 569900 690700
rect 570100 690500 570300 690700
rect 570500 690500 570700 690700
rect 570900 690500 571100 690700
rect 571300 690500 571500 690700
rect 571700 690500 572000 690700
rect 465100 690400 534200 690500
rect 47100 690300 73200 690400
rect 47100 690200 47200 690300
rect 47300 690200 73200 690300
rect 47100 690000 68400 690200
rect 68600 690000 68800 690200
rect 69000 690000 69200 690200
rect 69400 690000 69600 690200
rect 69800 690000 70000 690200
rect 70200 690000 70400 690200
rect 70600 690000 70800 690200
rect 71000 690000 71200 690200
rect 71400 690000 71600 690200
rect 71800 690000 72000 690200
rect 72200 690000 72400 690200
rect 72600 690000 72800 690200
rect 73000 690000 73200 690200
rect 47100 689800 47200 690000
rect 47300 689800 73200 690000
rect 47100 689600 68400 689800
rect 68600 689600 68800 689800
rect 69000 689600 69200 689800
rect 69400 689600 69600 689800
rect 69800 689600 70000 689800
rect 70200 689600 70400 689800
rect 70600 689600 70800 689800
rect 71000 689600 71200 689800
rect 71400 689600 71600 689800
rect 71800 689600 72000 689800
rect 72200 689600 72400 689800
rect 72600 689600 72800 689800
rect 73000 689600 73200 689800
rect 47100 689500 47200 689600
rect 47300 689500 73200 689600
rect 47100 689400 73200 689500
rect 465100 690200 532300 690400
rect 532500 690200 532700 690400
rect 532900 690200 533100 690400
rect 533300 690200 533500 690400
rect 533700 690200 533900 690400
rect 534100 690200 534200 690400
rect 465100 690100 534200 690200
rect 465100 689900 532300 690100
rect 532500 689900 532700 690100
rect 532900 689900 533100 690100
rect 533300 689900 533500 690100
rect 533700 689900 533900 690100
rect 534100 689900 534200 690100
rect 465100 689700 534200 689900
rect 465100 689500 532300 689700
rect 532500 689500 532700 689700
rect 532900 689500 533100 689700
rect 533300 689500 533500 689700
rect 533700 689500 533900 689700
rect 534100 689500 534200 689700
rect 465100 689300 534200 689500
rect 465100 689100 532300 689300
rect 532500 689100 532700 689300
rect 532900 689100 533100 689300
rect 533300 689100 533500 689300
rect 533700 689100 533900 689300
rect 534100 689100 534200 689300
rect 566200 690300 572000 690500
rect 566200 690100 566300 690300
rect 566500 690100 566700 690300
rect 566900 690100 567100 690300
rect 567300 690100 567500 690300
rect 567700 690100 567900 690300
rect 568100 690100 568300 690300
rect 568500 690100 568700 690300
rect 568900 690100 569100 690300
rect 569300 690100 569500 690300
rect 569700 690100 569900 690300
rect 570100 690100 570300 690300
rect 570500 690100 570700 690300
rect 570900 690100 571100 690300
rect 571300 690100 571500 690300
rect 571700 690100 572000 690300
rect 566200 689900 572000 690100
rect 566200 689700 566300 689900
rect 566500 689700 566700 689900
rect 566900 689700 567100 689900
rect 567300 689700 567500 689900
rect 567700 689700 567900 689900
rect 568100 689700 568300 689900
rect 568500 689700 568700 689900
rect 568900 689700 569100 689900
rect 569300 689700 569500 689900
rect 569700 689700 569900 689900
rect 570100 689700 570300 689900
rect 570500 689700 570700 689900
rect 570900 689700 571100 689900
rect 571300 689700 571500 689900
rect 571700 689700 572000 689900
rect 566200 689500 572000 689700
rect 566200 689300 566300 689500
rect 566500 689300 566700 689500
rect 566900 689300 567100 689500
rect 567300 689300 567500 689500
rect 567700 689300 567900 689500
rect 568100 689300 568300 689500
rect 568500 689300 568700 689500
rect 568900 689300 569100 689500
rect 569300 689300 569500 689500
rect 569700 689300 569900 689500
rect 570100 689300 570300 689500
rect 570500 689300 570700 689500
rect 570900 689300 571100 689500
rect 571300 689300 571500 689500
rect 571700 689300 572000 689500
rect 566200 689200 572000 689300
rect 465100 688900 534200 689100
rect 16200 688700 42200 688800
rect 16200 688500 16400 688700
rect 16600 688500 16800 688700
rect 17000 688500 17200 688700
rect 17400 688500 17600 688700
rect 17800 688500 18000 688700
rect 18200 688500 18400 688700
rect 18600 688500 18800 688700
rect 19000 688500 19200 688700
rect 19400 688500 19600 688700
rect 19800 688500 20000 688700
rect 20200 688500 20400 688700
rect 20600 688500 20800 688700
rect 21000 688600 42000 688700
rect 42100 688600 42200 688700
rect 465100 688700 532300 688900
rect 532500 688700 532700 688900
rect 532900 688700 533100 688900
rect 533300 688700 533500 688900
rect 533700 688700 533900 688900
rect 534100 688700 534200 688900
rect 465100 688600 534200 688700
rect 21000 688500 42200 688600
rect 16200 688300 42000 688500
rect 42100 688300 42200 688500
rect 16200 688100 16400 688300
rect 16600 688100 16800 688300
rect 17000 688100 17200 688300
rect 17400 688100 17600 688300
rect 17800 688100 18000 688300
rect 18200 688100 18400 688300
rect 18600 688100 18800 688300
rect 19000 688100 19200 688300
rect 19400 688100 19600 688300
rect 19800 688100 20000 688300
rect 20200 688100 20400 688300
rect 20600 688100 20800 688300
rect 21000 688200 42200 688300
rect 21000 688100 42000 688200
rect 42100 688100 42200 688200
rect 16200 688000 42200 688100
rect 36600 687300 47800 687400
rect 36600 687100 36800 687300
rect 37000 687100 37200 687300
rect 37400 687100 37600 687300
rect 37800 687100 38000 687300
rect 38200 687100 47800 687300
rect 36600 687000 47800 687100
rect 549890 687000 549900 687200
rect 550100 687000 550110 687200
rect 550190 687000 550200 687200
rect 550400 687000 550410 687200
rect 550490 687000 550500 687200
rect 550700 687000 550710 687200
rect 550790 687000 550800 687200
rect 551000 687000 551010 687200
rect 551190 687100 551200 687300
rect 551400 687100 551410 687300
rect 551190 686800 551200 687000
rect 551400 686800 551410 687000
rect 551190 686500 551200 686700
rect 551400 686500 551410 686700
rect 551190 686200 551200 686400
rect 551400 686200 551410 686400
rect 549790 685900 549800 686100
rect 550000 685900 550010 686100
rect 550090 685900 550100 686100
rect 550300 685900 550310 686100
rect 550390 685900 550400 686100
rect 550600 685900 550610 686100
rect 550790 685900 550800 686100
rect 551000 685900 551010 686100
rect 0 685300 38400 685400
rect 0 685242 36800 685300
rect -800 685100 36800 685242
rect 37000 685100 37200 685300
rect 37400 685100 37600 685300
rect 37800 685100 38000 685300
rect 38200 685100 38400 685300
rect -800 684900 38400 685100
rect -800 684700 36800 684900
rect 37000 684700 37200 684900
rect 37400 684700 37600 684900
rect 37800 684700 38000 684900
rect 38200 684700 38400 684900
rect -800 684500 38400 684700
rect -800 684300 36800 684500
rect 37000 684300 37200 684500
rect 37400 684300 37600 684500
rect 37800 684300 38000 684500
rect 38200 684300 38400 684500
rect -800 684100 38400 684300
rect -800 683900 36800 684100
rect 37000 683900 37200 684100
rect 37400 683900 37600 684100
rect 37800 683900 38000 684100
rect 38200 683900 38400 684100
rect -800 683700 38400 683900
rect -800 683500 36800 683700
rect 37000 683500 37200 683700
rect 37400 683500 37600 683700
rect 37800 683500 38000 683700
rect 38200 683500 38400 683700
rect -800 683300 38400 683500
rect -800 683100 36800 683300
rect 37000 683100 37200 683300
rect 37400 683100 37600 683300
rect 37800 683100 38000 683300
rect 38200 683100 38400 683300
rect 515500 684800 540560 684940
rect 515500 684600 515700 684800
rect 515900 684600 516100 684800
rect 516300 684600 516500 684800
rect 516700 684600 516900 684800
rect 517100 684600 517300 684800
rect 517500 684600 517700 684800
rect 517900 684600 518100 684800
rect 518300 684600 518500 684800
rect 518700 684600 518900 684800
rect 519100 684600 519300 684800
rect 519500 684600 519700 684800
rect 519900 684600 520100 684800
rect 520300 684600 520500 684800
rect 520700 684600 540560 684800
rect 515500 684400 540560 684600
rect 515500 684200 515700 684400
rect 515900 684200 516100 684400
rect 516300 684200 516500 684400
rect 516700 684200 516900 684400
rect 517100 684200 517300 684400
rect 517500 684200 517700 684400
rect 517900 684200 518100 684400
rect 518300 684200 518500 684400
rect 518700 684200 518900 684400
rect 519100 684200 519300 684400
rect 519500 684200 519700 684400
rect 519900 684200 520100 684400
rect 520300 684200 520500 684400
rect 520700 684200 540560 684400
rect 515500 684000 540560 684200
rect 515500 683800 515700 684000
rect 515900 683800 516100 684000
rect 516300 683800 516500 684000
rect 516700 683800 516900 684000
rect 517100 683800 517300 684000
rect 517500 683800 517700 684000
rect 517900 683800 518100 684000
rect 518300 683800 518500 684000
rect 518700 683800 518900 684000
rect 519100 683800 519300 684000
rect 519500 683800 519700 684000
rect 519900 683800 520100 684000
rect 520300 683800 520500 684000
rect 520700 683800 540560 684000
rect 515500 683600 540560 683800
rect 576600 684700 578700 684900
rect 576600 684400 576800 684700
rect 577100 684400 577300 684700
rect 577600 684400 577800 684700
rect 578100 684400 578300 684700
rect 578600 684400 578700 684700
rect 576600 684200 578700 684400
rect 576600 683900 576800 684200
rect 577100 683900 577300 684200
rect 577600 683900 577800 684200
rect 578100 683900 578300 684200
rect 578600 683900 578700 684200
rect 576600 683600 578700 683900
rect 582320 684600 582660 684660
rect 582320 684520 582360 684600
rect 582440 684520 582540 684600
rect 582620 684520 582660 684600
rect 582320 684440 582660 684520
rect 582320 684360 582360 684440
rect 582440 684360 582540 684440
rect 582620 684360 582660 684440
rect 582320 684280 582660 684360
rect 582320 684200 582360 684280
rect 582440 684200 582540 684280
rect 582620 684200 582660 684280
rect 582320 684100 582660 684200
rect 582320 684020 582360 684100
rect 582440 684020 582540 684100
rect 582620 684020 582660 684100
rect 582320 683940 582660 684020
rect 582320 683860 582360 683940
rect 582440 683860 582540 683940
rect 582620 683860 582660 683940
rect 515500 683400 515700 683600
rect 515900 683400 516100 683600
rect 516300 683400 516500 683600
rect 516700 683400 516900 683600
rect 517100 683400 517300 683600
rect 517500 683400 517700 683600
rect 517900 683400 518100 683600
rect 518300 683400 518500 683600
rect 518700 683400 518900 683600
rect 519100 683400 519300 683600
rect 519500 683400 519700 683600
rect 519900 683400 520100 683600
rect 520300 683400 520500 683600
rect 520700 683400 540560 683600
rect 515500 683200 540560 683400
rect 582320 683200 582660 683860
rect -800 682900 38400 683100
rect 42240 683120 43910 683140
rect 42240 683040 42260 683120
rect 42340 683040 42400 683120
rect 42480 683040 42540 683120
rect 42620 683040 43910 683120
rect 42240 683020 43910 683040
rect 45360 683120 47040 683140
rect 45360 683040 46660 683120
rect 46740 683040 46800 683120
rect 46880 683040 46940 683120
rect 47020 683040 47040 683120
rect 45360 683020 47040 683040
rect -800 682700 36800 682900
rect 37000 682700 37200 682900
rect 37400 682700 37600 682900
rect 37800 682700 38000 682900
rect 38200 682700 38400 682900
rect -800 682500 38400 682700
rect -800 682300 36800 682500
rect 37000 682300 37200 682500
rect 37400 682300 37600 682500
rect 37800 682300 38000 682500
rect 38200 682300 38400 682500
rect 515500 683000 515700 683200
rect 515900 683000 516100 683200
rect 516300 683000 516500 683200
rect 516700 683000 516900 683200
rect 517100 683000 517300 683200
rect 517500 683000 517700 683200
rect 517900 683000 518100 683200
rect 518300 683000 518500 683200
rect 518700 683000 518900 683200
rect 519100 683000 519300 683200
rect 519500 683000 519700 683200
rect 519900 683000 520100 683200
rect 520300 683000 520500 683200
rect 520700 683000 540560 683200
rect 515500 682800 540560 683000
rect 515500 682600 515700 682800
rect 515900 682600 516100 682800
rect 516300 682600 516500 682800
rect 516700 682600 516900 682800
rect 517100 682600 517300 682800
rect 517500 682600 517700 682800
rect 517900 682600 518100 682800
rect 518300 682600 518500 682800
rect 518700 682600 518900 682800
rect 519100 682600 519300 682800
rect 519500 682600 519700 682800
rect 519900 682600 520100 682800
rect 520300 682600 520500 682800
rect 520700 682600 540560 682800
rect 515500 682460 540560 682600
rect 561600 682984 584000 683200
rect 515500 682400 515600 682460
rect -800 682100 38400 682300
rect -800 681900 36800 682100
rect 37000 681900 37200 682100
rect 37400 681900 37600 682100
rect 37800 681900 38000 682100
rect 38200 681900 38400 682100
rect -800 681700 38400 681900
rect 45440 682200 62200 682320
rect 45440 682000 58000 682200
rect 58200 682000 58400 682200
rect 58600 682000 58800 682200
rect 59000 682000 59200 682200
rect 59400 682000 59600 682200
rect 59800 682000 60000 682200
rect 60200 682000 60400 682200
rect 60600 682000 60800 682200
rect 61000 682000 61200 682200
rect 61400 682000 61600 682200
rect 61800 682000 62200 682200
rect 45440 681860 62200 682000
rect 561600 682200 584800 682984
rect 561600 682000 561700 682200
rect 561900 682000 562100 682200
rect 562300 682000 562500 682200
rect 562700 682000 562900 682200
rect 563100 682000 563300 682200
rect 563500 682000 584800 682200
rect -800 681500 36800 681700
rect 37000 681500 37200 681700
rect 37400 681500 37600 681700
rect 37800 681500 38000 681700
rect 38200 681500 38400 681700
rect 561600 681800 584800 682000
rect 561600 681600 561700 681800
rect 561900 681600 562100 681800
rect 562300 681600 562500 681800
rect 562700 681600 562900 681800
rect 563100 681600 563300 681800
rect 563500 681600 584800 681800
rect -800 681300 38400 681500
rect -800 681100 36800 681300
rect 37000 681100 37200 681300
rect 37400 681100 37600 681300
rect 37800 681100 38000 681300
rect 38200 681100 38400 681300
rect -800 680900 38400 681100
rect -800 680700 36800 680900
rect 37000 680700 37200 680900
rect 37400 680700 37600 680900
rect 37800 680700 38000 680900
rect 38200 680700 38400 680900
rect 547600 681400 553100 681500
rect 547600 681200 549800 681400
rect 550000 681200 550200 681400
rect 550400 681200 550600 681400
rect 550800 681200 551000 681400
rect 551200 681200 551400 681400
rect 551600 681200 551800 681400
rect 552000 681200 552200 681400
rect 552400 681200 552600 681400
rect 552800 681200 553100 681400
rect 547600 681000 553100 681200
rect 547600 680800 549800 681000
rect 550000 680800 550200 681000
rect 550400 680800 550600 681000
rect 550800 680800 551000 681000
rect 551200 680800 551400 681000
rect 551600 680800 551800 681000
rect 552000 680800 552200 681000
rect 552400 680800 552600 681000
rect 552800 680800 553100 681000
rect 547600 680700 553100 680800
rect 561600 681400 584800 681600
rect 561600 681200 561700 681400
rect 561900 681200 562100 681400
rect 562300 681200 562500 681400
rect 562700 681200 562900 681400
rect 563100 681200 563300 681400
rect 563500 681200 584800 681400
rect 561600 681000 584800 681200
rect 561600 680800 561700 681000
rect 561900 680800 562100 681000
rect 562300 680800 562500 681000
rect 562700 680800 562900 681000
rect 563100 680800 563300 681000
rect 563500 680800 584800 681000
rect -800 680500 38400 680700
rect -800 680300 36800 680500
rect 37000 680300 37200 680500
rect 37400 680300 37600 680500
rect 37800 680300 38000 680500
rect 38200 680300 38400 680500
rect -800 680242 38400 680300
rect 0 680200 38400 680242
rect 561600 680600 584800 680800
rect 561600 680400 561700 680600
rect 561900 680400 562100 680600
rect 562300 680400 562500 680600
rect 562700 680400 562900 680600
rect 563100 680400 563300 680600
rect 563500 680400 584800 680600
rect 561600 680200 584800 680400
rect 561600 680000 561700 680200
rect 561900 680000 562100 680200
rect 562300 680000 562500 680200
rect 562700 680000 562900 680200
rect 563100 680000 563300 680200
rect 563500 680000 584800 680200
rect 561600 679800 584800 680000
rect 561600 679600 561700 679800
rect 561900 679600 562100 679800
rect 562300 679600 562500 679800
rect 562700 679600 562900 679800
rect 563100 679600 563300 679800
rect 563500 679600 584800 679800
rect 515500 679200 541760 679560
rect 515500 679000 515900 679200
rect 516100 679000 516300 679200
rect 516500 679000 516700 679200
rect 516900 679000 517100 679200
rect 517300 679000 517500 679200
rect 517700 679000 517900 679200
rect 518100 679000 518300 679200
rect 518500 679000 518700 679200
rect 518900 679000 519100 679200
rect 519300 679000 519500 679200
rect 519700 679000 519900 679200
rect 520100 679000 520300 679200
rect 520500 679000 520700 679200
rect 520900 679000 541760 679200
rect 515500 678800 541760 679000
rect 515500 678600 515900 678800
rect 516100 678600 516300 678800
rect 516500 678600 516700 678800
rect 516900 678600 517100 678800
rect 517300 678600 517500 678800
rect 517700 678600 517900 678800
rect 518100 678600 518300 678800
rect 518500 678600 518700 678800
rect 518900 678600 519100 678800
rect 519300 678600 519500 678800
rect 519700 678600 519900 678800
rect 520100 678600 520300 678800
rect 520500 678600 520700 678800
rect 520900 678600 541760 678800
rect 515500 678400 541760 678600
rect 515500 678200 515900 678400
rect 516100 678200 516300 678400
rect 516500 678200 516700 678400
rect 516900 678200 517100 678400
rect 517300 678200 517500 678400
rect 517700 678200 517900 678400
rect 518100 678200 518300 678400
rect 518500 678200 518700 678400
rect 518900 678200 519100 678400
rect 519300 678200 519500 678400
rect 519700 678200 519900 678400
rect 520100 678200 520300 678400
rect 520500 678200 520700 678400
rect 520900 678200 541760 678400
rect 515500 678000 541760 678200
rect 515500 677800 515900 678000
rect 516100 677800 516300 678000
rect 516500 677800 516700 678000
rect 516900 677800 517100 678000
rect 517300 677800 517500 678000
rect 517700 677800 517900 678000
rect 518100 677800 518300 678000
rect 518500 677800 518700 678000
rect 518900 677800 519100 678000
rect 519300 677800 519500 678000
rect 519700 677800 519900 678000
rect 520100 677800 520300 678000
rect 520500 677800 520700 678000
rect 520900 677800 541760 678000
rect 561600 679400 584800 679600
rect 561600 679200 561700 679400
rect 561900 679200 562100 679400
rect 562300 679200 562500 679400
rect 562700 679200 562900 679400
rect 563100 679200 563300 679400
rect 563500 679200 584800 679400
rect 561600 679000 584800 679200
rect 561600 678800 561700 679000
rect 561900 678800 562100 679000
rect 562300 678800 562500 679000
rect 562700 678800 562900 679000
rect 563100 678800 563300 679000
rect 563500 678800 584800 679000
rect 561600 678600 584800 678800
rect 561600 678400 561700 678600
rect 561900 678400 562100 678600
rect 562300 678400 562500 678600
rect 562700 678400 562900 678600
rect 563100 678400 563300 678600
rect 563500 678400 584800 678600
rect 561600 677984 584800 678400
rect 561600 677800 584000 677984
rect 515500 677600 541760 677800
rect 515500 677400 515900 677600
rect 516100 677400 516300 677600
rect 516500 677400 516700 677600
rect 516900 677400 517100 677600
rect 517300 677400 517500 677600
rect 517700 677400 517900 677600
rect 518100 677400 518300 677600
rect 518500 677400 518700 677600
rect 518900 677400 519100 677600
rect 519300 677400 519500 677600
rect 519700 677400 519900 677600
rect 520100 677400 520300 677600
rect 520500 677400 520700 677600
rect 520900 677400 541760 677600
rect 515500 677200 541760 677400
rect 515500 677000 515900 677200
rect 516100 677000 516300 677200
rect 516500 677000 516700 677200
rect 516900 677000 517100 677200
rect 517300 677000 517500 677200
rect 517700 677000 517900 677200
rect 518100 677000 518300 677200
rect 518500 677000 518700 677200
rect 518900 677000 519100 677200
rect 519300 677000 519500 677200
rect 519700 677000 519900 677200
rect 520100 677000 520300 677200
rect 520500 677000 520700 677200
rect 520900 677000 541760 677200
rect 515500 676800 541760 677000
rect 515500 676600 515900 676800
rect 516100 676600 516300 676800
rect 516500 676600 516700 676800
rect 516900 676600 517100 676800
rect 517300 676600 517500 676800
rect 517700 676600 517900 676800
rect 518100 676600 518300 676800
rect 518500 676600 518700 676800
rect 518900 676600 519100 676800
rect 519300 676600 519500 676800
rect 519700 676600 519900 676800
rect 520100 676600 520300 676800
rect 520500 676600 520700 676800
rect 520900 676600 541760 676800
rect 515500 676460 541760 676600
rect 547600 677300 572280 677400
rect 547600 677100 571900 677300
rect 572100 677100 572280 677300
rect 547600 677000 572280 677100
rect 547600 676800 571900 677000
rect 572100 676800 572280 677000
rect 547600 676700 572280 676800
rect 547600 676500 571900 676700
rect 572100 676500 572280 676700
rect 547600 676400 572280 676500
rect 547600 676200 571900 676400
rect 572100 676200 572280 676400
rect 547600 676100 572280 676200
rect 576700 676100 578700 677800
rect 32790 663300 33110 663305
rect 32790 663000 32800 663300
rect 33100 663000 33110 663300
rect 32790 662995 33110 663000
rect 33290 663300 33610 663305
rect 33290 663000 33300 663300
rect 33600 663000 33610 663300
rect 33290 662995 33610 663000
rect 33790 663300 34110 663305
rect 33790 663000 33800 663300
rect 34100 663000 34110 663300
rect 33790 662995 34110 663000
rect 34290 663300 34610 663305
rect 34290 663000 34300 663300
rect 34600 663000 34610 663300
rect 34290 662995 34610 663000
rect 34790 663300 35110 663305
rect 34790 663000 34800 663300
rect 35100 663000 35110 663300
rect 34790 662995 35110 663000
rect 35290 663300 35610 663305
rect 35290 663000 35300 663300
rect 35600 663000 35610 663300
rect 35290 662995 35610 663000
rect 35790 663300 36110 663305
rect 35790 663000 35800 663300
rect 36100 663000 36110 663300
rect 35790 662995 36110 663000
rect 36290 663300 36610 663305
rect 36290 663000 36300 663300
rect 36600 663000 36610 663300
rect 36290 662995 36610 663000
rect 36790 663300 37110 663305
rect 36790 663000 36800 663300
rect 37100 663000 37110 663300
rect 36790 662995 37110 663000
rect 37290 663300 37610 663305
rect 37290 663000 37300 663300
rect 37600 663000 37610 663300
rect 37290 662995 37610 663000
rect 37790 663300 38110 663305
rect 37790 663000 37800 663300
rect 38100 663000 38110 663300
rect 37790 662995 38110 663000
rect 38290 663300 38610 663305
rect 38290 663000 38300 663300
rect 38600 663000 38610 663300
rect 38290 662995 38610 663000
rect 38790 663300 39110 663305
rect 38790 663000 38800 663300
rect 39100 663000 39110 663300
rect 38790 662995 39110 663000
rect 39290 663300 39610 663305
rect 39290 663000 39300 663300
rect 39600 663000 39610 663300
rect 39290 662995 39610 663000
rect 39790 663300 40110 663305
rect 39790 663000 39800 663300
rect 40100 663000 40110 663300
rect 39790 662995 40110 663000
rect 40290 663300 40610 663305
rect 40290 663000 40300 663300
rect 40600 663000 40610 663300
rect 40290 662995 40610 663000
rect 0 648642 4000 648800
rect -800 648600 4000 648642
rect -800 648300 2500 648600
rect 2800 648300 3000 648600
rect 3300 648300 3500 648600
rect 3800 648300 4000 648600
rect -800 648100 4000 648300
rect -800 647800 2500 648100
rect 2800 647800 3000 648100
rect 3300 647800 3500 648100
rect 3800 647800 4000 648100
rect -800 647600 4000 647800
rect -800 647300 2500 647600
rect 2800 647300 3000 647600
rect 3300 647300 3500 647600
rect 3800 647300 4000 647600
rect -800 647100 4000 647300
rect -800 646800 2500 647100
rect 2800 646800 3000 647100
rect 3300 646800 3500 647100
rect 3800 646800 4000 647100
rect -800 646600 4000 646800
rect -800 646300 2500 646600
rect 2800 646300 3000 646600
rect 3300 646300 3500 646600
rect 3800 646300 4000 646600
rect -800 646100 4000 646300
rect -800 645800 2500 646100
rect 2800 645800 3000 646100
rect 3300 645800 3500 646100
rect 3800 645800 4000 646100
rect -800 645600 4000 645800
rect -800 645300 2500 645600
rect 2800 645300 3000 645600
rect 3300 645300 3500 645600
rect 3800 645300 4000 645600
rect -800 645100 4000 645300
rect -800 644800 2500 645100
rect 2800 644800 3000 645100
rect 3300 644800 3500 645100
rect 3800 644800 4000 645100
rect -800 644600 4000 644800
rect -800 644300 2500 644600
rect 2800 644300 3000 644600
rect 3300 644300 3500 644600
rect 3800 644300 4000 644600
rect -800 644100 4000 644300
rect -800 643842 2500 644100
rect 0 643800 2500 643842
rect 2800 643800 3000 644100
rect 3300 643800 3500 644100
rect 3800 643800 4000 644100
rect 0 643600 4000 643800
rect 0 643300 2500 643600
rect 2800 643300 3000 643600
rect 3300 643300 3500 643600
rect 3800 643300 4000 643600
rect 0 643100 4000 643300
rect 0 642800 2500 643100
rect 2800 642800 3000 643100
rect 3300 642800 3500 643100
rect 3800 642800 4000 643100
rect 0 642600 4000 642800
rect 0 642300 2500 642600
rect 2800 642300 3000 642600
rect 3300 642300 3500 642600
rect 3800 642300 4000 642600
rect 0 642100 4000 642300
rect 0 641800 2500 642100
rect 2800 641800 3000 642100
rect 3300 641800 3500 642100
rect 3800 641800 4000 642100
rect 0 641600 4000 641800
rect 0 641300 2500 641600
rect 2800 641300 3000 641600
rect 3300 641300 3500 641600
rect 3800 641300 4000 641600
rect 0 641100 4000 641300
rect 0 640800 2500 641100
rect 2800 640800 3000 641100
rect 3300 640800 3500 641100
rect 3800 640800 4000 641100
rect 0 640600 4000 640800
rect 0 640300 2500 640600
rect 2800 640300 3000 640600
rect 3300 640300 3500 640600
rect 3800 640300 4000 640600
rect 0 640100 4000 640300
rect 0 639800 2500 640100
rect 2800 639800 3000 640100
rect 3300 639800 3500 640100
rect 3800 639800 4000 640100
rect 0 639600 4000 639800
rect 0 639300 2500 639600
rect 2800 639300 3000 639600
rect 3300 639300 3500 639600
rect 3800 639300 4000 639600
rect 0 639100 4000 639300
rect 0 638800 2500 639100
rect 2800 638800 3000 639100
rect 3300 638800 3500 639100
rect 3800 638800 4000 639100
rect 0 638642 4000 638800
rect -800 638600 4000 638642
rect -800 638300 2500 638600
rect 2800 638300 3000 638600
rect 3300 638300 3500 638600
rect 3800 638300 4000 638600
rect -800 638100 4000 638300
rect -800 637800 2500 638100
rect 2800 637800 3000 638100
rect 3300 637800 3500 638100
rect 3800 637800 4000 638100
rect -800 637600 4000 637800
rect -800 637300 2500 637600
rect 2800 637300 3000 637600
rect 3300 637300 3500 637600
rect 3800 637300 4000 637600
rect -800 637100 4000 637300
rect -800 636800 2500 637100
rect 2800 636800 3000 637100
rect 3300 636800 3500 637100
rect 3800 636800 4000 637100
rect -800 636600 4000 636800
rect -800 636300 2500 636600
rect 2800 636300 3000 636600
rect 3300 636300 3500 636600
rect 3800 636300 4000 636600
rect -800 636100 4000 636300
rect -800 635800 2500 636100
rect 2800 635800 3000 636100
rect 3300 635800 3500 636100
rect 3800 635800 4000 636100
rect -800 635600 4000 635800
rect -800 635300 2500 635600
rect 2800 635300 3000 635600
rect 3300 635300 3500 635600
rect 3800 635300 4000 635600
rect -800 635100 4000 635300
rect -800 634800 2500 635100
rect 2800 634800 3000 635100
rect 3300 634800 3500 635100
rect 3800 634800 4000 635100
rect -800 634600 4000 634800
rect -800 634300 2500 634600
rect 2800 634300 3000 634600
rect 3300 634300 3500 634600
rect 3800 634300 4000 634600
rect -800 633842 4000 634300
rect 0 633800 4000 633842
rect 549600 644600 584000 644800
rect 549600 644400 550000 644600
rect 550200 644400 550400 644600
rect 550600 644400 550800 644600
rect 551000 644400 551200 644600
rect 551400 644400 551600 644600
rect 551800 644400 552000 644600
rect 552200 644400 552400 644600
rect 552600 644400 552800 644600
rect 553000 644584 584000 644600
rect 553000 644400 584800 644584
rect 549600 644200 584800 644400
rect 549600 644000 550000 644200
rect 550200 644000 550400 644200
rect 550600 644000 550800 644200
rect 551000 644000 551200 644200
rect 551400 644000 551600 644200
rect 551800 644000 552000 644200
rect 552200 644000 552400 644200
rect 552600 644000 552800 644200
rect 553000 644000 584800 644200
rect 549600 643800 584800 644000
rect 549600 643600 550000 643800
rect 550200 643600 550400 643800
rect 550600 643600 550800 643800
rect 551000 643600 551200 643800
rect 551400 643600 551600 643800
rect 551800 643600 552000 643800
rect 552200 643600 552400 643800
rect 552600 643600 552800 643800
rect 553000 643600 584800 643800
rect 549600 643400 584800 643600
rect 549600 643200 550000 643400
rect 550200 643200 550400 643400
rect 550600 643200 550800 643400
rect 551000 643200 551200 643400
rect 551400 643200 551600 643400
rect 551800 643200 552000 643400
rect 552200 643200 552400 643400
rect 552600 643200 552800 643400
rect 553000 643200 584800 643400
rect 549600 643000 584800 643200
rect 549600 642800 550000 643000
rect 550200 642800 550400 643000
rect 550600 642800 550800 643000
rect 551000 642800 551200 643000
rect 551400 642800 551600 643000
rect 551800 642800 552000 643000
rect 552200 642800 552400 643000
rect 552600 642800 552800 643000
rect 553000 642800 584800 643000
rect 549600 642600 584800 642800
rect 549600 642400 550000 642600
rect 550200 642400 550400 642600
rect 550600 642400 550800 642600
rect 551000 642400 551200 642600
rect 551400 642400 551600 642600
rect 551800 642400 552000 642600
rect 552200 642400 552400 642600
rect 552600 642400 552800 642600
rect 553000 642400 584800 642600
rect 549600 642200 584800 642400
rect 549600 642000 550000 642200
rect 550200 642000 550400 642200
rect 550600 642000 550800 642200
rect 551000 642000 551200 642200
rect 551400 642000 551600 642200
rect 551800 642000 552000 642200
rect 552200 642000 552400 642200
rect 552600 642000 552800 642200
rect 553000 642000 584800 642200
rect 549600 641800 584800 642000
rect 549600 641600 550000 641800
rect 550200 641600 550400 641800
rect 550600 641600 550800 641800
rect 551000 641600 551200 641800
rect 551400 641600 551600 641800
rect 551800 641600 552000 641800
rect 552200 641600 552400 641800
rect 552600 641600 552800 641800
rect 553000 641600 584800 641800
rect 549600 641400 584800 641600
rect 549600 641200 550000 641400
rect 550200 641200 550400 641400
rect 550600 641200 550800 641400
rect 551000 641200 551200 641400
rect 551400 641200 551600 641400
rect 551800 641200 552000 641400
rect 552200 641200 552400 641400
rect 552600 641200 552800 641400
rect 553000 641200 584800 641400
rect 549600 641000 584800 641200
rect 549600 640800 550000 641000
rect 550200 640800 550400 641000
rect 550600 640800 550800 641000
rect 551000 640800 551200 641000
rect 551400 640800 551600 641000
rect 551800 640800 552000 641000
rect 552200 640800 552400 641000
rect 552600 640800 552800 641000
rect 553000 640800 584800 641000
rect 549600 640600 584800 640800
rect 549600 640400 550000 640600
rect 550200 640400 550400 640600
rect 550600 640400 550800 640600
rect 551000 640400 551200 640600
rect 551400 640400 551600 640600
rect 551800 640400 552000 640600
rect 552200 640400 552400 640600
rect 552600 640400 552800 640600
rect 553000 640400 584800 640600
rect 549600 640200 584800 640400
rect 549600 640000 550000 640200
rect 550200 640000 550400 640200
rect 550600 640000 550800 640200
rect 551000 640000 551200 640200
rect 551400 640000 551600 640200
rect 551800 640000 552000 640200
rect 552200 640000 552400 640200
rect 552600 640000 552800 640200
rect 553000 640000 584800 640200
rect 549600 639800 584800 640000
rect 549600 639600 550000 639800
rect 550200 639600 550400 639800
rect 550600 639600 550800 639800
rect 551000 639600 551200 639800
rect 551400 639600 551600 639800
rect 551800 639600 552000 639800
rect 552200 639600 552400 639800
rect 552600 639600 552800 639800
rect 553000 639784 584800 639800
rect 553000 639600 584000 639784
rect 549600 639400 584000 639600
rect 549600 639200 550000 639400
rect 550200 639200 550400 639400
rect 550600 639200 550800 639400
rect 551000 639200 551200 639400
rect 551400 639200 551600 639400
rect 551800 639200 552000 639400
rect 552200 639200 552400 639400
rect 552600 639200 552800 639400
rect 553000 639200 584000 639400
rect 549600 639000 584000 639200
rect 549600 638800 550000 639000
rect 550200 638800 550400 639000
rect 550600 638800 550800 639000
rect 551000 638800 551200 639000
rect 551400 638800 551600 639000
rect 551800 638800 552000 639000
rect 552200 638800 552400 639000
rect 552600 638800 552800 639000
rect 553000 638800 584000 639000
rect 549600 638600 584000 638800
rect 549600 638400 550000 638600
rect 550200 638400 550400 638600
rect 550600 638400 550800 638600
rect 551000 638400 551200 638600
rect 551400 638400 551600 638600
rect 551800 638400 552000 638600
rect 552200 638400 552400 638600
rect 552600 638400 552800 638600
rect 553000 638400 584000 638600
rect 549600 638200 584000 638400
rect 549600 638000 550000 638200
rect 550200 638000 550400 638200
rect 550600 638000 550800 638200
rect 551000 638000 551200 638200
rect 551400 638000 551600 638200
rect 551800 638000 552000 638200
rect 552200 638000 552400 638200
rect 552600 638000 552800 638200
rect 553000 638000 584000 638200
rect 549600 637800 584000 638000
rect 549600 637600 550000 637800
rect 550200 637600 550400 637800
rect 550600 637600 550800 637800
rect 551000 637600 551200 637800
rect 551400 637600 551600 637800
rect 551800 637600 552000 637800
rect 552200 637600 552400 637800
rect 552600 637600 552800 637800
rect 553000 637600 584000 637800
rect 549600 637400 584000 637600
rect 549600 637200 550000 637400
rect 550200 637200 550400 637400
rect 550600 637200 550800 637400
rect 551000 637200 551200 637400
rect 551400 637200 551600 637400
rect 551800 637200 552000 637400
rect 552200 637200 552400 637400
rect 552600 637200 552800 637400
rect 553000 637200 584000 637400
rect 549600 637000 584000 637200
rect 549600 636800 550000 637000
rect 550200 636800 550400 637000
rect 550600 636800 550800 637000
rect 551000 636800 551200 637000
rect 551400 636800 551600 637000
rect 551800 636800 552000 637000
rect 552200 636800 552400 637000
rect 552600 636800 552800 637000
rect 553000 636800 584000 637000
rect 549600 636600 584000 636800
rect 549600 636400 550000 636600
rect 550200 636400 550400 636600
rect 550600 636400 550800 636600
rect 551000 636400 551200 636600
rect 551400 636400 551600 636600
rect 551800 636400 552000 636600
rect 552200 636400 552400 636600
rect 552600 636400 552800 636600
rect 553000 636400 584000 636600
rect 549600 636200 584000 636400
rect 549600 636000 550000 636200
rect 550200 636000 550400 636200
rect 550600 636000 550800 636200
rect 551000 636000 551200 636200
rect 551400 636000 551600 636200
rect 551800 636000 552000 636200
rect 552200 636000 552400 636200
rect 552600 636000 552800 636200
rect 553000 636000 584000 636200
rect 549600 635800 584000 636000
rect 549600 635600 550000 635800
rect 550200 635600 550400 635800
rect 550600 635600 550800 635800
rect 551000 635600 551200 635800
rect 551400 635600 551600 635800
rect 551800 635600 552000 635800
rect 552200 635600 552400 635800
rect 552600 635600 552800 635800
rect 553000 635600 584000 635800
rect 549600 635400 584000 635600
rect 549600 635200 550000 635400
rect 550200 635200 550400 635400
rect 550600 635200 550800 635400
rect 551000 635200 551200 635400
rect 551400 635200 551600 635400
rect 551800 635200 552000 635400
rect 552200 635200 552400 635400
rect 552600 635200 552800 635400
rect 553000 635200 584000 635400
rect 549600 635000 584000 635200
rect 549600 634800 550000 635000
rect 550200 634800 550400 635000
rect 550600 634800 550800 635000
rect 551000 634800 551200 635000
rect 551400 634800 551600 635000
rect 551800 634800 552000 635000
rect 552200 634800 552400 635000
rect 552600 634800 552800 635000
rect 553000 634800 584000 635000
rect 549600 634600 584000 634800
rect 549600 634400 550000 634600
rect 550200 634400 550400 634600
rect 550600 634400 550800 634600
rect 551000 634400 551200 634600
rect 551400 634400 551600 634600
rect 551800 634400 552000 634600
rect 552200 634400 552400 634600
rect 552600 634400 552800 634600
rect 553000 634584 584000 634600
rect 553000 634400 584800 634584
rect 549600 634200 584800 634400
rect 549600 634000 550000 634200
rect 550200 634000 550400 634200
rect 550600 634000 550800 634200
rect 551000 634000 551200 634200
rect 551400 634000 551600 634200
rect 551800 634000 552000 634200
rect 552200 634000 552400 634200
rect 552600 634000 552800 634200
rect 553000 634000 584800 634200
rect 549600 633800 584800 634000
rect 549600 633600 550000 633800
rect 550200 633600 550400 633800
rect 550600 633600 550800 633800
rect 551000 633600 551200 633800
rect 551400 633600 551600 633800
rect 551800 633600 552000 633800
rect 552200 633600 552400 633800
rect 552600 633600 552800 633800
rect 553000 633600 584800 633800
rect 549600 633400 584800 633600
rect 549600 633200 550000 633400
rect 550200 633200 550400 633400
rect 550600 633200 550800 633400
rect 551000 633200 551200 633400
rect 551400 633200 551600 633400
rect 551800 633200 552000 633400
rect 552200 633200 552400 633400
rect 552600 633200 552800 633400
rect 553000 633200 584800 633400
rect 549600 633000 584800 633200
rect 549600 632800 550000 633000
rect 550200 632800 550400 633000
rect 550600 632800 550800 633000
rect 551000 632800 551200 633000
rect 551400 632800 551600 633000
rect 551800 632800 552000 633000
rect 552200 632800 552400 633000
rect 552600 632800 552800 633000
rect 553000 632800 584800 633000
rect 549600 632600 584800 632800
rect 549600 632400 550000 632600
rect 550200 632400 550400 632600
rect 550600 632400 550800 632600
rect 551000 632400 551200 632600
rect 551400 632400 551600 632600
rect 551800 632400 552000 632600
rect 552200 632400 552400 632600
rect 552600 632400 552800 632600
rect 553000 632400 584800 632600
rect 549600 632200 584800 632400
rect 549600 632000 550000 632200
rect 550200 632000 550400 632200
rect 550600 632000 550800 632200
rect 551000 632000 551200 632200
rect 551400 632000 551600 632200
rect 551800 632000 552000 632200
rect 552200 632000 552400 632200
rect 552600 632000 552800 632200
rect 553000 632000 584800 632200
rect 549600 631800 584800 632000
rect 549600 631600 550000 631800
rect 550200 631600 550400 631800
rect 550600 631600 550800 631800
rect 551000 631600 551200 631800
rect 551400 631600 551600 631800
rect 551800 631600 552000 631800
rect 552200 631600 552400 631800
rect 552600 631600 552800 631800
rect 553000 631600 584800 631800
rect 549600 631400 584800 631600
rect 549600 631200 550000 631400
rect 550200 631200 550400 631400
rect 550600 631200 550800 631400
rect 551000 631200 551200 631400
rect 551400 631200 551600 631400
rect 551800 631200 552000 631400
rect 552200 631200 552400 631400
rect 552600 631200 552800 631400
rect 553000 631200 584800 631400
rect 549600 631000 584800 631200
rect 549600 630800 550000 631000
rect 550200 630800 550400 631000
rect 550600 630800 550800 631000
rect 551000 630800 551200 631000
rect 551400 630800 551600 631000
rect 551800 630800 552000 631000
rect 552200 630800 552400 631000
rect 552600 630800 552800 631000
rect 553000 630800 584800 631000
rect 549600 630700 584800 630800
rect 549600 630500 550000 630700
rect 550200 630500 550400 630700
rect 550600 630500 550800 630700
rect 551000 630500 551200 630700
rect 551400 630500 551600 630700
rect 551800 630500 552000 630700
rect 552200 630500 552400 630700
rect 552600 630500 552800 630700
rect 553000 630500 584800 630700
rect 549600 630400 584800 630500
rect 549600 630200 550000 630400
rect 550200 630200 550400 630400
rect 550600 630200 550800 630400
rect 551000 630200 551200 630400
rect 551400 630200 551600 630400
rect 551800 630200 552000 630400
rect 552200 630200 552400 630400
rect 552600 630200 552800 630400
rect 553000 630200 584800 630400
rect 549600 630000 584800 630200
rect 549600 629800 550000 630000
rect 550200 629800 550400 630000
rect 550600 629800 550800 630000
rect 551000 629800 551200 630000
rect 551400 629800 551600 630000
rect 551800 629800 552000 630000
rect 552200 629800 552400 630000
rect 552600 629800 552800 630000
rect 553000 629800 584800 630000
rect 549600 629784 584800 629800
rect 549600 629400 584000 629784
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 0 564242 12020 564300
rect -800 559442 12020 564242
rect 0 554242 12020 559442
rect -800 549442 12020 554242
rect 0 549400 12020 549442
rect 12540 564100 40800 564300
rect 12540 563900 32800 564100
rect 33000 563900 33200 564100
rect 33400 563900 33600 564100
rect 33800 563900 34000 564100
rect 34200 563900 34400 564100
rect 34600 563900 34800 564100
rect 35000 563900 35200 564100
rect 35400 563900 35600 564100
rect 35800 563900 36000 564100
rect 36200 563900 36400 564100
rect 36600 563900 36800 564100
rect 37000 563900 37200 564100
rect 37400 563900 37600 564100
rect 37800 563900 38000 564100
rect 38200 563900 38400 564100
rect 38600 563900 38800 564100
rect 39000 563900 39200 564100
rect 39400 563900 39600 564100
rect 39800 563900 40000 564100
rect 40200 563900 40400 564100
rect 40600 563900 40800 564100
rect 12540 563700 40800 563900
rect 12540 563500 32800 563700
rect 33000 563500 33200 563700
rect 33400 563500 33600 563700
rect 33800 563500 34000 563700
rect 34200 563500 34400 563700
rect 34600 563500 34800 563700
rect 35000 563500 35200 563700
rect 35400 563500 35600 563700
rect 35800 563500 36000 563700
rect 36200 563500 36400 563700
rect 36600 563500 36800 563700
rect 37000 563500 37200 563700
rect 37400 563500 37600 563700
rect 37800 563500 38000 563700
rect 38200 563500 38400 563700
rect 38600 563500 38800 563700
rect 39000 563500 39200 563700
rect 39400 563500 39600 563700
rect 39800 563500 40000 563700
rect 40200 563500 40400 563700
rect 40600 563500 40800 563700
rect 12540 563300 40800 563500
rect 12540 563100 32800 563300
rect 33000 563100 33200 563300
rect 33400 563100 33600 563300
rect 33800 563100 34000 563300
rect 34200 563100 34400 563300
rect 34600 563100 34800 563300
rect 35000 563100 35200 563300
rect 35400 563100 35600 563300
rect 35800 563100 36000 563300
rect 36200 563100 36400 563300
rect 36600 563100 36800 563300
rect 37000 563100 37200 563300
rect 37400 563100 37600 563300
rect 37800 563100 38000 563300
rect 38200 563100 38400 563300
rect 38600 563100 38800 563300
rect 39000 563100 39200 563300
rect 39400 563100 39600 563300
rect 39800 563100 40000 563300
rect 40200 563100 40400 563300
rect 40600 563220 40800 563300
rect 40600 563100 40760 563220
rect 12540 563060 40760 563100
rect 12540 562900 40800 563060
rect 12540 562700 32800 562900
rect 33000 562700 33200 562900
rect 33400 562700 33600 562900
rect 33800 562700 34000 562900
rect 34200 562700 34400 562900
rect 34600 562700 34800 562900
rect 35000 562700 35200 562900
rect 35400 562700 35600 562900
rect 35800 562700 36000 562900
rect 36200 562700 36400 562900
rect 36600 562700 36800 562900
rect 37000 562700 37200 562900
rect 37400 562700 37600 562900
rect 37800 562700 38000 562900
rect 38200 562700 38400 562900
rect 38600 562700 38800 562900
rect 39000 562700 39200 562900
rect 39400 562700 39600 562900
rect 39800 562700 40000 562900
rect 40200 562700 40400 562900
rect 40600 562700 40800 562900
rect 12540 562500 40800 562700
rect 12540 562300 32800 562500
rect 33000 562300 33200 562500
rect 33400 562300 33600 562500
rect 33800 562300 34000 562500
rect 34200 562300 34400 562500
rect 34600 562300 34800 562500
rect 35000 562300 35200 562500
rect 35400 562300 35600 562500
rect 35800 562300 36000 562500
rect 36200 562300 36400 562500
rect 36600 562300 36800 562500
rect 37000 562300 37200 562500
rect 37400 562300 37600 562500
rect 37800 562300 38000 562500
rect 38200 562300 38400 562500
rect 38600 562300 38800 562500
rect 39000 562300 39200 562500
rect 39400 562300 39600 562500
rect 39800 562300 40000 562500
rect 40200 562300 40400 562500
rect 40600 562300 40800 562500
rect 12540 562100 40800 562300
rect 12540 561900 32800 562100
rect 33000 561900 33200 562100
rect 33400 561900 33600 562100
rect 33800 561900 34000 562100
rect 34200 561900 34400 562100
rect 34600 561900 34800 562100
rect 35000 561900 35200 562100
rect 35400 561900 35600 562100
rect 35800 561900 36000 562100
rect 36200 561900 36400 562100
rect 36600 561900 36800 562100
rect 37000 561900 37200 562100
rect 37400 561900 37600 562100
rect 37800 561900 38000 562100
rect 38200 561900 38400 562100
rect 38600 561900 38800 562100
rect 39000 561900 39200 562100
rect 39400 561900 39600 562100
rect 39800 561900 40000 562100
rect 40200 561900 40400 562100
rect 40600 561900 40800 562100
rect 12540 561700 40800 561900
rect 12540 561500 32800 561700
rect 33000 561500 33200 561700
rect 33400 561500 33600 561700
rect 33800 561500 34000 561700
rect 34200 561500 34400 561700
rect 34600 561500 34800 561700
rect 35000 561500 35200 561700
rect 35400 561500 35600 561700
rect 35800 561500 36000 561700
rect 36200 561500 36400 561700
rect 36600 561500 36800 561700
rect 37000 561500 37200 561700
rect 37400 561500 37600 561700
rect 37800 561500 38000 561700
rect 38200 561500 38400 561700
rect 38600 561500 38800 561700
rect 39000 561500 39200 561700
rect 39400 561500 39600 561700
rect 39800 561500 40000 561700
rect 40200 561500 40400 561700
rect 40600 561500 40800 561700
rect 12540 561300 40800 561500
rect 12540 561100 32800 561300
rect 33000 561100 33200 561300
rect 33400 561100 33600 561300
rect 33800 561100 34000 561300
rect 34200 561100 34400 561300
rect 34600 561100 34800 561300
rect 35000 561100 35200 561300
rect 35400 561100 35600 561300
rect 35800 561100 36000 561300
rect 36200 561100 36400 561300
rect 36600 561100 36800 561300
rect 37000 561100 37200 561300
rect 37400 561100 37600 561300
rect 37800 561100 38000 561300
rect 38200 561100 38400 561300
rect 38600 561100 38800 561300
rect 39000 561100 39200 561300
rect 39400 561100 39600 561300
rect 39800 561100 40000 561300
rect 40200 561100 40400 561300
rect 40600 561100 40800 561300
rect 12540 560900 40800 561100
rect 12540 560700 32800 560900
rect 33000 560700 33200 560900
rect 33400 560700 33600 560900
rect 33800 560700 34000 560900
rect 34200 560700 34400 560900
rect 34600 560700 34800 560900
rect 35000 560700 35200 560900
rect 35400 560700 35600 560900
rect 35800 560700 36000 560900
rect 36200 560700 36400 560900
rect 36600 560700 36800 560900
rect 37000 560700 37200 560900
rect 37400 560700 37600 560900
rect 37800 560700 38000 560900
rect 38200 560700 38400 560900
rect 38600 560700 38800 560900
rect 39000 560700 39200 560900
rect 39400 560700 39600 560900
rect 39800 560700 40000 560900
rect 40200 560700 40400 560900
rect 40600 560700 40800 560900
rect 12540 560500 40800 560700
rect 12540 560300 32800 560500
rect 33000 560300 33200 560500
rect 33400 560300 33600 560500
rect 33800 560300 34000 560500
rect 34200 560300 34400 560500
rect 34600 560300 34800 560500
rect 35000 560300 35200 560500
rect 35400 560300 35600 560500
rect 35800 560300 36000 560500
rect 36200 560300 36400 560500
rect 36600 560300 36800 560500
rect 37000 560300 37200 560500
rect 37400 560300 37600 560500
rect 37800 560300 38000 560500
rect 38200 560300 38400 560500
rect 38600 560300 38800 560500
rect 39000 560300 39200 560500
rect 39400 560300 39600 560500
rect 39800 560300 40000 560500
rect 40200 560300 40400 560500
rect 40600 560300 40800 560500
rect 12540 560100 40800 560300
rect 12540 559900 32800 560100
rect 33000 559900 33200 560100
rect 33400 559900 33600 560100
rect 33800 559900 34000 560100
rect 34200 559900 34400 560100
rect 34600 559900 34800 560100
rect 35000 559900 35200 560100
rect 35400 559900 35600 560100
rect 35800 559900 36000 560100
rect 36200 559900 36400 560100
rect 36600 559900 36800 560100
rect 37000 559900 37200 560100
rect 37400 559900 37600 560100
rect 37800 559900 38000 560100
rect 38200 559900 38400 560100
rect 38600 559900 38800 560100
rect 39000 559900 39200 560100
rect 39400 559900 39600 560100
rect 39800 559900 40000 560100
rect 40200 559900 40400 560100
rect 40600 559900 40800 560100
rect 12540 559700 40800 559900
rect 12540 559500 32800 559700
rect 33000 559500 33200 559700
rect 33400 559500 33600 559700
rect 33800 559500 34000 559700
rect 34200 559500 34400 559700
rect 34600 559500 34800 559700
rect 35000 559500 35200 559700
rect 35400 559500 35600 559700
rect 35800 559500 36000 559700
rect 36200 559500 36400 559700
rect 36600 559500 36800 559700
rect 37000 559500 37200 559700
rect 37400 559500 37600 559700
rect 37800 559500 38000 559700
rect 38200 559500 38400 559700
rect 38600 559500 38800 559700
rect 39000 559500 39200 559700
rect 39400 559500 39600 559700
rect 39800 559500 40000 559700
rect 40200 559500 40400 559700
rect 40600 559500 40800 559700
rect 12540 559300 40800 559500
rect 12540 559100 32800 559300
rect 33000 559100 33200 559300
rect 33400 559100 33600 559300
rect 33800 559100 34000 559300
rect 34200 559100 34400 559300
rect 34600 559100 34800 559300
rect 35000 559100 35200 559300
rect 35400 559100 35600 559300
rect 35800 559100 36000 559300
rect 36200 559100 36400 559300
rect 36600 559100 36800 559300
rect 37000 559100 37200 559300
rect 37400 559100 37600 559300
rect 37800 559100 38000 559300
rect 38200 559100 38400 559300
rect 38600 559100 38800 559300
rect 39000 559100 39200 559300
rect 39400 559100 39600 559300
rect 39800 559100 40000 559300
rect 40200 559100 40400 559300
rect 40600 559100 40800 559300
rect 12540 558900 40800 559100
rect 12540 558700 32800 558900
rect 33000 558700 33200 558900
rect 33400 558700 33600 558900
rect 33800 558700 34000 558900
rect 34200 558700 34400 558900
rect 34600 558700 34800 558900
rect 35000 558700 35200 558900
rect 35400 558700 35600 558900
rect 35800 558700 36000 558900
rect 36200 558700 36400 558900
rect 36600 558700 36800 558900
rect 37000 558700 37200 558900
rect 37400 558700 37600 558900
rect 37800 558700 38000 558900
rect 38200 558700 38400 558900
rect 38600 558700 38800 558900
rect 39000 558700 39200 558900
rect 39400 558700 39600 558900
rect 39800 558700 40000 558900
rect 40200 558700 40400 558900
rect 40600 558700 40800 558900
rect 12540 558500 40800 558700
rect 12540 558300 32800 558500
rect 33000 558300 33200 558500
rect 33400 558300 33600 558500
rect 33800 558300 34000 558500
rect 34200 558300 34400 558500
rect 34600 558300 34800 558500
rect 35000 558300 35200 558500
rect 35400 558300 35600 558500
rect 35800 558300 36000 558500
rect 36200 558300 36400 558500
rect 36600 558300 36800 558500
rect 37000 558300 37200 558500
rect 37400 558300 37600 558500
rect 37800 558300 38000 558500
rect 38200 558300 38400 558500
rect 38600 558300 38800 558500
rect 39000 558300 39200 558500
rect 39400 558300 39600 558500
rect 39800 558300 40000 558500
rect 40200 558300 40400 558500
rect 40600 558300 40800 558500
rect 12540 558100 40800 558300
rect 12540 557900 32800 558100
rect 33000 557900 33200 558100
rect 33400 557900 33600 558100
rect 33800 557900 34000 558100
rect 34200 557900 34400 558100
rect 34600 557900 34800 558100
rect 35000 557900 35200 558100
rect 35400 557900 35600 558100
rect 35800 557900 36000 558100
rect 36200 557900 36400 558100
rect 36600 557900 36800 558100
rect 37000 557900 37200 558100
rect 37400 557900 37600 558100
rect 37800 557900 38000 558100
rect 38200 557900 38400 558100
rect 38600 557900 38800 558100
rect 39000 557900 39200 558100
rect 39400 557900 39600 558100
rect 39800 557900 40000 558100
rect 40200 557900 40400 558100
rect 40600 557900 40800 558100
rect 12540 557700 40800 557900
rect 12540 557500 32800 557700
rect 33000 557500 33200 557700
rect 33400 557500 33600 557700
rect 33800 557500 34000 557700
rect 34200 557500 34400 557700
rect 34600 557500 34800 557700
rect 35000 557500 35200 557700
rect 35400 557500 35600 557700
rect 35800 557500 36000 557700
rect 36200 557500 36400 557700
rect 36600 557500 36800 557700
rect 37000 557500 37200 557700
rect 37400 557500 37600 557700
rect 37800 557500 38000 557700
rect 38200 557500 38400 557700
rect 38600 557500 38800 557700
rect 39000 557500 39200 557700
rect 39400 557500 39600 557700
rect 39800 557500 40000 557700
rect 40200 557500 40400 557700
rect 40600 557500 40800 557700
rect 12540 557300 40800 557500
rect 12540 557100 32800 557300
rect 33000 557100 33200 557300
rect 33400 557100 33600 557300
rect 33800 557100 34000 557300
rect 34200 557100 34400 557300
rect 34600 557100 34800 557300
rect 35000 557100 35200 557300
rect 35400 557100 35600 557300
rect 35800 557100 36000 557300
rect 36200 557100 36400 557300
rect 36600 557100 36800 557300
rect 37000 557100 37200 557300
rect 37400 557100 37600 557300
rect 37800 557100 38000 557300
rect 38200 557100 38400 557300
rect 38600 557100 38800 557300
rect 39000 557100 39200 557300
rect 39400 557100 39600 557300
rect 39800 557100 40000 557300
rect 40200 557100 40400 557300
rect 40600 557100 40800 557300
rect 12540 556900 40800 557100
rect 12540 556700 32800 556900
rect 33000 556700 33200 556900
rect 33400 556700 33600 556900
rect 33800 556700 34000 556900
rect 34200 556700 34400 556900
rect 34600 556700 34800 556900
rect 35000 556700 35200 556900
rect 35400 556700 35600 556900
rect 35800 556700 36000 556900
rect 36200 556700 36400 556900
rect 36600 556700 36800 556900
rect 37000 556700 37200 556900
rect 37400 556700 37600 556900
rect 37800 556700 38000 556900
rect 38200 556700 38400 556900
rect 38600 556700 38800 556900
rect 39000 556700 39200 556900
rect 39400 556700 39600 556900
rect 39800 556700 40000 556900
rect 40200 556700 40400 556900
rect 40600 556700 40800 556900
rect 12540 556500 40800 556700
rect 12540 556300 32800 556500
rect 33000 556300 33200 556500
rect 33400 556300 33600 556500
rect 33800 556300 34000 556500
rect 34200 556300 34400 556500
rect 34600 556300 34800 556500
rect 35000 556300 35200 556500
rect 35400 556300 35600 556500
rect 35800 556300 36000 556500
rect 36200 556300 36400 556500
rect 36600 556300 36800 556500
rect 37000 556300 37200 556500
rect 37400 556300 37600 556500
rect 37800 556300 38000 556500
rect 38200 556300 38400 556500
rect 38600 556300 38800 556500
rect 39000 556300 39200 556500
rect 39400 556300 39600 556500
rect 39800 556300 40000 556500
rect 40200 556300 40400 556500
rect 40600 556300 40800 556500
rect 12540 556100 40800 556300
rect 12540 555900 32800 556100
rect 33000 555900 33200 556100
rect 33400 555900 33600 556100
rect 33800 555900 34000 556100
rect 34200 555900 34400 556100
rect 34600 555900 34800 556100
rect 35000 555900 35200 556100
rect 35400 555900 35600 556100
rect 35800 555900 36000 556100
rect 36200 555900 36400 556100
rect 36600 555900 36800 556100
rect 37000 555900 37200 556100
rect 37400 555900 37600 556100
rect 37800 555900 38000 556100
rect 38200 555900 38400 556100
rect 38600 555900 38800 556100
rect 39000 555900 39200 556100
rect 39400 555900 39600 556100
rect 39800 555900 40000 556100
rect 40200 555900 40400 556100
rect 40600 555900 40800 556100
rect 12540 555700 40800 555900
rect 12540 555500 32800 555700
rect 33000 555500 33200 555700
rect 33400 555500 33600 555700
rect 33800 555500 34000 555700
rect 34200 555500 34400 555700
rect 34600 555500 34800 555700
rect 35000 555500 35200 555700
rect 35400 555500 35600 555700
rect 35800 555500 36000 555700
rect 36200 555500 36400 555700
rect 36600 555500 36800 555700
rect 37000 555500 37200 555700
rect 37400 555500 37600 555700
rect 37800 555500 38000 555700
rect 38200 555500 38400 555700
rect 38600 555500 38800 555700
rect 39000 555500 39200 555700
rect 39400 555500 39600 555700
rect 39800 555500 40000 555700
rect 40200 555500 40400 555700
rect 40600 555500 40800 555700
rect 12540 555300 40800 555500
rect 12540 555100 32800 555300
rect 33000 555100 33200 555300
rect 33400 555100 33600 555300
rect 33800 555100 34000 555300
rect 34200 555100 34400 555300
rect 34600 555100 34800 555300
rect 35000 555100 35200 555300
rect 35400 555100 35600 555300
rect 35800 555100 36000 555300
rect 36200 555100 36400 555300
rect 36600 555100 36800 555300
rect 37000 555100 37200 555300
rect 37400 555100 37600 555300
rect 37800 555100 38000 555300
rect 38200 555100 38400 555300
rect 38600 555100 38800 555300
rect 39000 555100 39200 555300
rect 39400 555100 39600 555300
rect 39800 555100 40000 555300
rect 40200 555100 40400 555300
rect 40600 555100 40800 555300
rect 12540 554900 40800 555100
rect 12540 554700 32800 554900
rect 33000 554700 33200 554900
rect 33400 554700 33600 554900
rect 33800 554700 34000 554900
rect 34200 554700 34400 554900
rect 34600 554700 34800 554900
rect 35000 554700 35200 554900
rect 35400 554700 35600 554900
rect 35800 554700 36000 554900
rect 36200 554700 36400 554900
rect 36600 554700 36800 554900
rect 37000 554700 37200 554900
rect 37400 554700 37600 554900
rect 37800 554700 38000 554900
rect 38200 554700 38400 554900
rect 38600 554700 38800 554900
rect 39000 554700 39200 554900
rect 39400 554700 39600 554900
rect 39800 554700 40000 554900
rect 40200 554700 40400 554900
rect 40600 554700 40800 554900
rect 12540 554500 40800 554700
rect 12540 554300 32800 554500
rect 33000 554300 33200 554500
rect 33400 554300 33600 554500
rect 33800 554300 34000 554500
rect 34200 554300 34400 554500
rect 34600 554300 34800 554500
rect 35000 554300 35200 554500
rect 35400 554300 35600 554500
rect 35800 554300 36000 554500
rect 36200 554300 36400 554500
rect 36600 554300 36800 554500
rect 37000 554300 37200 554500
rect 37400 554300 37600 554500
rect 37800 554300 38000 554500
rect 38200 554300 38400 554500
rect 38600 554300 38800 554500
rect 39000 554300 39200 554500
rect 39400 554300 39600 554500
rect 39800 554300 40000 554500
rect 40200 554300 40400 554500
rect 40600 554300 40800 554500
rect 12540 554100 40800 554300
rect 12540 553900 32800 554100
rect 33000 553900 33200 554100
rect 33400 553900 33600 554100
rect 33800 553900 34000 554100
rect 34200 553900 34400 554100
rect 34600 553900 34800 554100
rect 35000 553900 35200 554100
rect 35400 553900 35600 554100
rect 35800 553900 36000 554100
rect 36200 553900 36400 554100
rect 36600 553900 36800 554100
rect 37000 553900 37200 554100
rect 37400 553900 37600 554100
rect 37800 553900 38000 554100
rect 38200 553900 38400 554100
rect 38600 553900 38800 554100
rect 39000 553900 39200 554100
rect 39400 553900 39600 554100
rect 39800 553900 40000 554100
rect 40200 553900 40400 554100
rect 40600 553900 40800 554100
rect 12540 553700 40800 553900
rect 12540 553500 32800 553700
rect 33000 553500 33200 553700
rect 33400 553500 33600 553700
rect 33800 553500 34000 553700
rect 34200 553500 34400 553700
rect 34600 553500 34800 553700
rect 35000 553500 35200 553700
rect 35400 553500 35600 553700
rect 35800 553500 36000 553700
rect 36200 553500 36400 553700
rect 36600 553500 36800 553700
rect 37000 553500 37200 553700
rect 37400 553500 37600 553700
rect 37800 553500 38000 553700
rect 38200 553500 38400 553700
rect 38600 553500 38800 553700
rect 39000 553500 39200 553700
rect 39400 553500 39600 553700
rect 39800 553500 40000 553700
rect 40200 553500 40400 553700
rect 40600 553500 40800 553700
rect 12540 553300 40800 553500
rect 12540 553100 32800 553300
rect 33000 553100 33200 553300
rect 33400 553100 33600 553300
rect 33800 553100 34000 553300
rect 34200 553100 34400 553300
rect 34600 553100 34800 553300
rect 35000 553100 35200 553300
rect 35400 553100 35600 553300
rect 35800 553100 36000 553300
rect 36200 553100 36400 553300
rect 36600 553100 36800 553300
rect 37000 553100 37200 553300
rect 37400 553100 37600 553300
rect 37800 553100 38000 553300
rect 38200 553100 38400 553300
rect 38600 553100 38800 553300
rect 39000 553100 39200 553300
rect 39400 553100 39600 553300
rect 39800 553100 40000 553300
rect 40200 553100 40400 553300
rect 40600 553100 40800 553300
rect 12540 552900 40800 553100
rect 12540 552700 32800 552900
rect 33000 552700 33200 552900
rect 33400 552700 33600 552900
rect 33800 552700 34000 552900
rect 34200 552700 34400 552900
rect 34600 552700 34800 552900
rect 35000 552700 35200 552900
rect 35400 552700 35600 552900
rect 35800 552700 36000 552900
rect 36200 552700 36400 552900
rect 36600 552700 36800 552900
rect 37000 552700 37200 552900
rect 37400 552700 37600 552900
rect 37800 552700 38000 552900
rect 38200 552700 38400 552900
rect 38600 552700 38800 552900
rect 39000 552700 39200 552900
rect 39400 552700 39600 552900
rect 39800 552700 40000 552900
rect 40200 552700 40400 552900
rect 40600 552700 40800 552900
rect 12540 552500 40800 552700
rect 12540 552300 32800 552500
rect 33000 552300 33200 552500
rect 33400 552300 33600 552500
rect 33800 552300 34000 552500
rect 34200 552300 34400 552500
rect 34600 552300 34800 552500
rect 35000 552300 35200 552500
rect 35400 552300 35600 552500
rect 35800 552300 36000 552500
rect 36200 552300 36400 552500
rect 36600 552300 36800 552500
rect 37000 552300 37200 552500
rect 37400 552300 37600 552500
rect 37800 552300 38000 552500
rect 38200 552300 38400 552500
rect 38600 552300 38800 552500
rect 39000 552300 39200 552500
rect 39400 552300 39600 552500
rect 39800 552300 40000 552500
rect 40200 552300 40400 552500
rect 40600 552300 40800 552500
rect 12540 552100 40800 552300
rect 12540 551900 32800 552100
rect 33000 551900 33200 552100
rect 33400 551900 33600 552100
rect 33800 551900 34000 552100
rect 34200 551900 34400 552100
rect 34600 551900 34800 552100
rect 35000 551900 35200 552100
rect 35400 551900 35600 552100
rect 35800 551900 36000 552100
rect 36200 551900 36400 552100
rect 36600 551900 36800 552100
rect 37000 551900 37200 552100
rect 37400 551900 37600 552100
rect 37800 551900 38000 552100
rect 38200 551900 38400 552100
rect 38600 551900 38800 552100
rect 39000 551900 39200 552100
rect 39400 551900 39600 552100
rect 39800 551900 40000 552100
rect 40200 551900 40400 552100
rect 40600 551900 40800 552100
rect 12540 551700 40800 551900
rect 12540 551500 32800 551700
rect 33000 551500 33200 551700
rect 33400 551500 33600 551700
rect 33800 551500 34000 551700
rect 34200 551500 34400 551700
rect 34600 551500 34800 551700
rect 35000 551500 35200 551700
rect 35400 551500 35600 551700
rect 35800 551500 36000 551700
rect 36200 551500 36400 551700
rect 36600 551500 36800 551700
rect 37000 551500 37200 551700
rect 37400 551500 37600 551700
rect 37800 551500 38000 551700
rect 38200 551500 38400 551700
rect 38600 551500 38800 551700
rect 39000 551500 39200 551700
rect 39400 551500 39600 551700
rect 39800 551500 40000 551700
rect 40200 551500 40400 551700
rect 40600 551500 40800 551700
rect 12540 551300 40800 551500
rect 12540 551100 32800 551300
rect 33000 551100 33200 551300
rect 33400 551100 33600 551300
rect 33800 551100 34000 551300
rect 34200 551100 34400 551300
rect 34600 551100 34800 551300
rect 35000 551100 35200 551300
rect 35400 551100 35600 551300
rect 35800 551100 36000 551300
rect 36200 551100 36400 551300
rect 36600 551100 36800 551300
rect 37000 551100 37200 551300
rect 37400 551100 37600 551300
rect 37800 551100 38000 551300
rect 38200 551100 38400 551300
rect 38600 551100 38800 551300
rect 39000 551100 39200 551300
rect 39400 551100 39600 551300
rect 39800 551100 40000 551300
rect 40200 551100 40400 551300
rect 40600 551100 40800 551300
rect 12540 550900 40800 551100
rect 12540 550700 32800 550900
rect 33000 550700 33200 550900
rect 33400 550700 33600 550900
rect 33800 550700 34000 550900
rect 34200 550700 34400 550900
rect 34600 550700 34800 550900
rect 35000 550700 35200 550900
rect 35400 550700 35600 550900
rect 35800 550700 36000 550900
rect 36200 550700 36400 550900
rect 36600 550700 36800 550900
rect 37000 550700 37200 550900
rect 37400 550700 37600 550900
rect 37800 550700 38000 550900
rect 38200 550700 38400 550900
rect 38600 550700 38800 550900
rect 39000 550700 39200 550900
rect 39400 550700 39600 550900
rect 39800 550700 40000 550900
rect 40200 550700 40400 550900
rect 40600 550700 40800 550900
rect 12540 550500 40800 550700
rect 582340 550562 584800 555362
rect 12540 550300 32800 550500
rect 33000 550300 33200 550500
rect 33400 550300 33600 550500
rect 33800 550300 34000 550500
rect 34200 550300 34400 550500
rect 34600 550300 34800 550500
rect 35000 550300 35200 550500
rect 35400 550300 35600 550500
rect 35800 550300 36000 550500
rect 36200 550300 36400 550500
rect 36600 550300 36800 550500
rect 37000 550300 37200 550500
rect 37400 550300 37600 550500
rect 37800 550300 38000 550500
rect 38200 550300 38400 550500
rect 38600 550300 38800 550500
rect 39000 550300 39200 550500
rect 39400 550300 39600 550500
rect 39800 550300 40000 550500
rect 40200 550300 40400 550500
rect 40600 550300 40800 550500
rect 12540 550100 40800 550300
rect 12540 549900 32800 550100
rect 33000 549900 33200 550100
rect 33400 549900 33600 550100
rect 33800 549900 34000 550100
rect 34200 549900 34400 550100
rect 34600 549900 34800 550100
rect 35000 549900 35200 550100
rect 35400 549900 35600 550100
rect 35800 549900 36000 550100
rect 36200 549900 36400 550100
rect 36600 549900 36800 550100
rect 37000 549900 37200 550100
rect 37400 549900 37600 550100
rect 37800 549900 38000 550100
rect 38200 549900 38400 550100
rect 38600 549900 38800 550100
rect 39000 549900 39200 550100
rect 39400 549900 39600 550100
rect 39800 549900 40000 550100
rect 40200 549900 40400 550100
rect 40600 549900 40800 550100
rect 12540 549700 40800 549900
rect 12540 549500 32800 549700
rect 33000 549500 33200 549700
rect 33400 549500 33600 549700
rect 33800 549500 34000 549700
rect 34200 549500 34400 549700
rect 34600 549500 34800 549700
rect 35000 549500 35200 549700
rect 35400 549500 35600 549700
rect 35800 549500 36000 549700
rect 36200 549500 36400 549700
rect 36600 549500 36800 549700
rect 37000 549500 37200 549700
rect 37400 549500 37600 549700
rect 37800 549500 38000 549700
rect 38200 549500 38400 549700
rect 38600 549500 38800 549700
rect 39000 549500 39200 549700
rect 39400 549500 39600 549700
rect 39800 549500 40000 549700
rect 40200 549500 40400 549700
rect 40600 549500 40800 549700
rect 12540 549400 40800 549500
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 12020 549400 12540 564300
<< via3 >>
rect 16400 702000 16600 702200
rect 16800 702000 17000 702200
rect 17200 702000 17400 702200
rect 17600 702000 17800 702200
rect 18000 702000 18200 702200
rect 18400 702000 18600 702200
rect 18800 702000 19000 702200
rect 19200 702000 19400 702200
rect 19600 702000 19800 702200
rect 20000 702000 20200 702200
rect 20400 702000 20600 702200
rect 20800 702000 21000 702200
rect 23400 702060 23520 702180
rect 23600 702060 23720 702180
rect 23800 702060 23920 702180
rect 24000 702060 24120 702180
rect 24200 702060 24320 702180
rect 65060 702080 65240 702260
rect 65400 702080 65580 702260
rect 65740 702080 65920 702260
rect 16400 701600 16600 701800
rect 16800 701600 17000 701800
rect 17200 701600 17400 701800
rect 17600 701600 17800 701800
rect 18000 701600 18200 701800
rect 18400 701600 18600 701800
rect 18800 701600 19000 701800
rect 19200 701600 19400 701800
rect 19600 701600 19800 701800
rect 20000 701600 20200 701800
rect 20400 701600 20600 701800
rect 20800 701600 21000 701800
rect 16400 701200 16600 701400
rect 16800 701200 17000 701400
rect 17200 701200 17400 701400
rect 17600 701200 17800 701400
rect 18000 701200 18200 701400
rect 18400 701200 18600 701400
rect 18800 701200 19000 701400
rect 19200 701200 19400 701400
rect 19600 701200 19800 701400
rect 20000 701200 20200 701400
rect 20400 701200 20600 701400
rect 20800 701200 21000 701400
rect 16400 700800 16600 701000
rect 16800 700800 17000 701000
rect 17200 700800 17400 701000
rect 17600 700800 17800 701000
rect 18000 700800 18200 701000
rect 18400 700800 18600 701000
rect 18800 700800 19000 701000
rect 19200 700800 19400 701000
rect 19600 700800 19800 701000
rect 20000 700800 20200 701000
rect 20400 700800 20600 701000
rect 20800 700800 21000 701000
rect 16400 700400 16600 700600
rect 16800 700400 17000 700600
rect 17200 700400 17400 700600
rect 17600 700400 17800 700600
rect 18000 700400 18200 700600
rect 18400 700400 18600 700600
rect 18800 700400 19000 700600
rect 19200 700400 19400 700600
rect 19600 700400 19800 700600
rect 20000 700400 20200 700600
rect 20400 700400 20600 700600
rect 20800 700400 21000 700600
rect 16400 700000 16600 700200
rect 16800 700000 17000 700200
rect 17200 700000 17400 700200
rect 17600 700000 17800 700200
rect 18000 700000 18200 700200
rect 18400 700000 18600 700200
rect 18800 700000 19000 700200
rect 19200 700000 19400 700200
rect 19600 700000 19800 700200
rect 20000 700000 20200 700200
rect 20400 700000 20600 700200
rect 20800 700000 21000 700200
rect 68400 702000 68600 702200
rect 68800 702000 69000 702200
rect 69200 702000 69400 702200
rect 69600 702000 69800 702200
rect 70000 702000 70200 702200
rect 70400 702000 70600 702200
rect 70800 702000 71000 702200
rect 71200 702000 71400 702200
rect 71600 702000 71800 702200
rect 72000 702000 72200 702200
rect 72400 702000 72600 702200
rect 72800 702000 73000 702200
rect 68400 701600 68600 701800
rect 68800 701600 69000 701800
rect 69200 701600 69400 701800
rect 69600 701600 69800 701800
rect 70000 701600 70200 701800
rect 70400 701600 70600 701800
rect 70800 701600 71000 701800
rect 71200 701600 71400 701800
rect 71600 701600 71800 701800
rect 72000 701600 72200 701800
rect 72400 701600 72600 701800
rect 72800 701600 73000 701800
rect 68400 701200 68600 701400
rect 68800 701200 69000 701400
rect 69200 701200 69400 701400
rect 69600 701200 69800 701400
rect 70000 701200 70200 701400
rect 70400 701200 70600 701400
rect 70800 701200 71000 701400
rect 71200 701200 71400 701400
rect 71600 701200 71800 701400
rect 72000 701200 72200 701400
rect 72400 701200 72600 701400
rect 72800 701200 73000 701400
rect 68400 700800 68600 701000
rect 68800 700800 69000 701000
rect 69200 700800 69400 701000
rect 69600 700800 69800 701000
rect 70000 700800 70200 701000
rect 70400 700800 70600 701000
rect 70800 700800 71000 701000
rect 71200 700800 71400 701000
rect 71600 700800 71800 701000
rect 72000 700800 72200 701000
rect 72400 700800 72600 701000
rect 72800 700800 73000 701000
rect 68400 700400 68600 700600
rect 68800 700400 69000 700600
rect 69200 700400 69400 700600
rect 69600 700400 69800 700600
rect 70000 700400 70200 700600
rect 70400 700400 70600 700600
rect 70800 700400 71000 700600
rect 71200 700400 71400 700600
rect 71600 700400 71800 700600
rect 72000 700400 72200 700600
rect 72400 700400 72600 700600
rect 72800 700400 73000 700600
rect 68400 700000 68600 700200
rect 68800 700000 69000 700200
rect 69200 700000 69400 700200
rect 69600 700000 69800 700200
rect 70000 700000 70200 700200
rect 70400 700000 70600 700200
rect 70800 700000 71000 700200
rect 71200 700000 71400 700200
rect 71600 700000 71800 700200
rect 72000 700000 72200 700200
rect 72400 700000 72600 700200
rect 72800 700000 73000 700200
rect 13000 698000 13200 698200
rect 13600 698000 13800 698200
rect 23400 698000 23600 698200
rect 23800 698000 24000 698200
rect 24200 698000 24400 698200
rect 65000 698000 65200 698200
rect 65600 698000 65800 698200
rect 75400 698000 75600 698200
rect 76000 698000 76200 698200
rect 13000 697600 13200 697800
rect 13600 697600 13800 697800
rect 23400 697600 23600 697800
rect 23800 697600 24000 697800
rect 24200 697600 24400 697800
rect 65000 697600 65200 697800
rect 65600 697600 65800 697800
rect 75400 697600 75600 697800
rect 76000 697600 76200 697800
rect 23400 697200 23600 697400
rect 23800 697200 24000 697400
rect 24200 697200 24400 697400
rect 65000 697200 65200 697400
rect 65600 697200 65800 697400
rect 75400 697200 75600 697400
rect 76000 697200 76200 697400
rect 13000 697000 13200 697200
rect 13600 697000 13800 697200
rect 23400 696800 23600 697000
rect 23800 696800 24000 697000
rect 24200 696800 24400 697000
rect 65000 696800 65200 697000
rect 65600 696800 65800 697000
rect 75400 696800 75600 697000
rect 76000 696800 76200 697000
rect 13000 696600 13200 696800
rect 13600 696600 13800 696800
rect 23400 696400 23600 696600
rect 23800 696400 24000 696600
rect 24200 696400 24400 696600
rect 65000 696400 65200 696600
rect 65600 696400 65800 696600
rect 75400 696400 75600 696600
rect 76000 696400 76200 696600
rect 38700 692840 38860 693000
rect 39120 692840 39280 693000
rect 38700 692620 38860 692780
rect 39120 692620 39280 692780
rect 49960 692860 50100 693000
rect 50180 692860 50320 693000
rect 50400 692860 50540 693000
rect 49960 692660 50100 692800
rect 50180 692660 50320 692800
rect 50400 692660 50540 692800
rect 38700 692400 38860 692560
rect 39120 692400 39280 692560
rect 38700 692180 38860 692340
rect 39120 692180 39280 692340
rect 12900 691700 13100 691900
rect 13200 691700 13400 691900
rect 13500 691700 13700 691900
rect 13800 691700 14000 691900
rect 58000 691700 58200 691900
rect 58400 691700 58600 691900
rect 58800 691700 59000 691900
rect 59200 691700 59400 691900
rect 59600 691700 59800 691900
rect 60000 691700 60200 691900
rect 60400 691700 60600 691900
rect 60800 691700 61000 691900
rect 61200 691700 61400 691900
rect 61600 691700 61800 691900
rect 515700 701400 515900 701600
rect 516100 701400 516300 701600
rect 516500 701400 516700 701600
rect 516900 701400 517100 701600
rect 517300 701400 517500 701600
rect 517700 701400 517900 701600
rect 518100 701400 518300 701600
rect 518500 701400 518700 701600
rect 518900 701400 519100 701600
rect 519300 701400 519500 701600
rect 519700 701400 519900 701600
rect 520100 701400 520300 701600
rect 520500 701400 520700 701600
rect 515700 701000 515900 701200
rect 516100 701000 516300 701200
rect 516500 701000 516700 701200
rect 516900 701000 517100 701200
rect 517300 701000 517500 701200
rect 517700 701000 517900 701200
rect 518100 701000 518300 701200
rect 518500 701000 518700 701200
rect 518900 701000 519100 701200
rect 519300 701000 519500 701200
rect 519700 701000 519900 701200
rect 520100 701000 520300 701200
rect 520500 701000 520700 701200
rect 515700 700600 515900 700800
rect 516100 700600 516300 700800
rect 516500 700600 516700 700800
rect 516900 700600 517100 700800
rect 517300 700600 517500 700800
rect 517700 700600 517900 700800
rect 518100 700600 518300 700800
rect 518500 700600 518700 700800
rect 518900 700600 519100 700800
rect 519300 700600 519500 700800
rect 519700 700600 519900 700800
rect 520100 700600 520300 700800
rect 520500 700600 520700 700800
rect 515700 700200 515900 700400
rect 516100 700200 516300 700400
rect 516500 700200 516700 700400
rect 516900 700200 517100 700400
rect 517300 700200 517500 700400
rect 517700 700200 517900 700400
rect 518100 700200 518300 700400
rect 518500 700200 518700 700400
rect 518900 700200 519100 700400
rect 519300 700200 519500 700400
rect 519700 700200 519900 700400
rect 520100 700200 520300 700400
rect 520500 700200 520700 700400
rect 515700 699800 515900 700000
rect 516100 699800 516300 700000
rect 516500 699800 516700 700000
rect 516900 699800 517100 700000
rect 517300 699800 517500 700000
rect 517700 699800 517900 700000
rect 518100 699800 518300 700000
rect 518500 699800 518700 700000
rect 518900 699800 519100 700000
rect 519300 699800 519500 700000
rect 519700 699800 519900 700000
rect 520100 699800 520300 700000
rect 520500 699800 520700 700000
rect 515700 699400 515900 699600
rect 516100 699400 516300 699600
rect 516500 699400 516700 699600
rect 516900 699400 517100 699600
rect 517300 699400 517500 699600
rect 517700 699400 517900 699600
rect 518100 699400 518300 699600
rect 518500 699400 518700 699600
rect 518900 699400 519100 699600
rect 519300 699400 519500 699600
rect 519700 699400 519900 699600
rect 520100 699400 520300 699600
rect 520500 699400 520700 699600
rect 515700 699000 515900 699200
rect 516100 699000 516300 699200
rect 516500 699000 516700 699200
rect 516900 699000 517100 699200
rect 517300 699000 517500 699200
rect 517700 699000 517900 699200
rect 518100 699000 518300 699200
rect 518500 699000 518700 699200
rect 518900 699000 519100 699200
rect 519300 699000 519500 699200
rect 519700 699000 519900 699200
rect 520100 699000 520300 699200
rect 520500 699000 520700 699200
rect 515700 697200 515900 697400
rect 516100 697200 516300 697400
rect 516500 697200 516700 697400
rect 516900 697200 517100 697400
rect 517300 697200 517500 697400
rect 517700 697200 517900 697400
rect 518100 697200 518300 697400
rect 518500 697200 518700 697400
rect 518900 697200 519100 697400
rect 519300 697200 519500 697400
rect 519700 697200 519900 697400
rect 520100 697200 520300 697400
rect 520500 697200 520700 697400
rect 515700 696800 515900 697000
rect 516100 696800 516300 697000
rect 516500 696800 516700 697000
rect 516900 696800 517100 697000
rect 517300 696800 517500 697000
rect 517700 696800 517900 697000
rect 518100 696800 518300 697000
rect 518500 696800 518700 697000
rect 518900 696800 519100 697000
rect 519300 696800 519500 697000
rect 519700 696800 519900 697000
rect 520100 696800 520300 697000
rect 520500 696800 520700 697000
rect 515700 696400 515900 696600
rect 516100 696400 516300 696600
rect 516500 696400 516700 696600
rect 516900 696400 517100 696600
rect 517300 696400 517500 696600
rect 517700 696400 517900 696600
rect 518100 696400 518300 696600
rect 518500 696400 518700 696600
rect 518900 696400 519100 696600
rect 519300 696400 519500 696600
rect 519700 696400 519900 696600
rect 520100 696400 520300 696600
rect 520500 696400 520700 696600
rect 573300 697800 573500 698000
rect 573800 697800 574000 698000
rect 573300 697400 573500 697600
rect 573800 697400 574000 697600
rect 573300 697000 573500 697200
rect 573800 697000 574000 697200
rect 573300 696600 573500 696800
rect 573800 696600 574000 696800
rect 573300 696200 573500 696400
rect 573800 696200 574000 696400
rect 68400 690000 68600 690200
rect 68800 690000 69000 690200
rect 69200 690000 69400 690200
rect 69600 690000 69800 690200
rect 70000 690000 70200 690200
rect 70400 690000 70600 690200
rect 70800 690000 71000 690200
rect 71200 690000 71400 690200
rect 71600 690000 71800 690200
rect 72000 690000 72200 690200
rect 72400 690000 72600 690200
rect 72800 690000 73000 690200
rect 68400 689600 68600 689800
rect 68800 689600 69000 689800
rect 69200 689600 69400 689800
rect 69600 689600 69800 689800
rect 70000 689600 70200 689800
rect 70400 689600 70600 689800
rect 70800 689600 71000 689800
rect 71200 689600 71400 689800
rect 71600 689600 71800 689800
rect 72000 689600 72200 689800
rect 72400 689600 72600 689800
rect 72800 689600 73000 689800
rect 532300 690200 532500 690400
rect 532700 690200 532900 690400
rect 533100 690200 533300 690400
rect 533500 690200 533700 690400
rect 533900 690200 534100 690400
rect 532300 689900 532500 690100
rect 532700 689900 532900 690100
rect 533100 689900 533300 690100
rect 533500 689900 533700 690100
rect 533900 689900 534100 690100
rect 532300 689500 532500 689700
rect 532700 689500 532900 689700
rect 533100 689500 533300 689700
rect 533500 689500 533700 689700
rect 533900 689500 534100 689700
rect 532300 689100 532500 689300
rect 532700 689100 532900 689300
rect 533100 689100 533300 689300
rect 533500 689100 533700 689300
rect 533900 689100 534100 689300
rect 16400 688500 16600 688700
rect 16800 688500 17000 688700
rect 17200 688500 17400 688700
rect 17600 688500 17800 688700
rect 18000 688500 18200 688700
rect 18400 688500 18600 688700
rect 18800 688500 19000 688700
rect 19200 688500 19400 688700
rect 19600 688500 19800 688700
rect 20000 688500 20200 688700
rect 20400 688500 20600 688700
rect 20800 688500 21000 688700
rect 532300 688700 532500 688900
rect 532700 688700 532900 688900
rect 533100 688700 533300 688900
rect 533500 688700 533700 688900
rect 533900 688700 534100 688900
rect 16400 688100 16600 688300
rect 16800 688100 17000 688300
rect 17200 688100 17400 688300
rect 17600 688100 17800 688300
rect 18000 688100 18200 688300
rect 18400 688100 18600 688300
rect 18800 688100 19000 688300
rect 19200 688100 19400 688300
rect 19600 688100 19800 688300
rect 20000 688100 20200 688300
rect 20400 688100 20600 688300
rect 20800 688100 21000 688300
rect 36800 687100 37000 687300
rect 37200 687100 37400 687300
rect 37600 687100 37800 687300
rect 38000 687100 38200 687300
rect 549900 687000 550100 687200
rect 550200 687000 550400 687200
rect 550500 687000 550700 687200
rect 550800 687000 551000 687200
rect 551200 687100 551400 687300
rect 551200 686800 551400 687000
rect 551200 686500 551400 686700
rect 551200 686200 551400 686400
rect 549800 685900 550000 686100
rect 550100 685900 550300 686100
rect 550400 685900 550600 686100
rect 550800 685900 551000 686100
rect 36800 685100 37000 685300
rect 37200 685100 37400 685300
rect 37600 685100 37800 685300
rect 38000 685100 38200 685300
rect 36800 684700 37000 684900
rect 37200 684700 37400 684900
rect 37600 684700 37800 684900
rect 38000 684700 38200 684900
rect 36800 684300 37000 684500
rect 37200 684300 37400 684500
rect 37600 684300 37800 684500
rect 38000 684300 38200 684500
rect 36800 683900 37000 684100
rect 37200 683900 37400 684100
rect 37600 683900 37800 684100
rect 38000 683900 38200 684100
rect 36800 683500 37000 683700
rect 37200 683500 37400 683700
rect 37600 683500 37800 683700
rect 38000 683500 38200 683700
rect 36800 683100 37000 683300
rect 37200 683100 37400 683300
rect 37600 683100 37800 683300
rect 38000 683100 38200 683300
rect 515700 684600 515900 684800
rect 516100 684600 516300 684800
rect 516500 684600 516700 684800
rect 516900 684600 517100 684800
rect 517300 684600 517500 684800
rect 517700 684600 517900 684800
rect 518100 684600 518300 684800
rect 518500 684600 518700 684800
rect 518900 684600 519100 684800
rect 519300 684600 519500 684800
rect 519700 684600 519900 684800
rect 520100 684600 520300 684800
rect 520500 684600 520700 684800
rect 515700 684200 515900 684400
rect 516100 684200 516300 684400
rect 516500 684200 516700 684400
rect 516900 684200 517100 684400
rect 517300 684200 517500 684400
rect 517700 684200 517900 684400
rect 518100 684200 518300 684400
rect 518500 684200 518700 684400
rect 518900 684200 519100 684400
rect 519300 684200 519500 684400
rect 519700 684200 519900 684400
rect 520100 684200 520300 684400
rect 520500 684200 520700 684400
rect 515700 683800 515900 684000
rect 516100 683800 516300 684000
rect 516500 683800 516700 684000
rect 516900 683800 517100 684000
rect 517300 683800 517500 684000
rect 517700 683800 517900 684000
rect 518100 683800 518300 684000
rect 518500 683800 518700 684000
rect 518900 683800 519100 684000
rect 519300 683800 519500 684000
rect 519700 683800 519900 684000
rect 520100 683800 520300 684000
rect 520500 683800 520700 684000
rect 576800 684400 577100 684700
rect 577300 684400 577600 684700
rect 577800 684400 578100 684700
rect 578300 684400 578600 684700
rect 576800 683900 577100 684200
rect 577300 683900 577600 684200
rect 577800 683900 578100 684200
rect 578300 683900 578600 684200
rect 515700 683400 515900 683600
rect 516100 683400 516300 683600
rect 516500 683400 516700 683600
rect 516900 683400 517100 683600
rect 517300 683400 517500 683600
rect 517700 683400 517900 683600
rect 518100 683400 518300 683600
rect 518500 683400 518700 683600
rect 518900 683400 519100 683600
rect 519300 683400 519500 683600
rect 519700 683400 519900 683600
rect 520100 683400 520300 683600
rect 520500 683400 520700 683600
rect 36800 682700 37000 682900
rect 37200 682700 37400 682900
rect 37600 682700 37800 682900
rect 38000 682700 38200 682900
rect 36800 682300 37000 682500
rect 37200 682300 37400 682500
rect 37600 682300 37800 682500
rect 38000 682300 38200 682500
rect 515700 683000 515900 683200
rect 516100 683000 516300 683200
rect 516500 683000 516700 683200
rect 516900 683000 517100 683200
rect 517300 683000 517500 683200
rect 517700 683000 517900 683200
rect 518100 683000 518300 683200
rect 518500 683000 518700 683200
rect 518900 683000 519100 683200
rect 519300 683000 519500 683200
rect 519700 683000 519900 683200
rect 520100 683000 520300 683200
rect 520500 683000 520700 683200
rect 515700 682600 515900 682800
rect 516100 682600 516300 682800
rect 516500 682600 516700 682800
rect 516900 682600 517100 682800
rect 517300 682600 517500 682800
rect 517700 682600 517900 682800
rect 518100 682600 518300 682800
rect 518500 682600 518700 682800
rect 518900 682600 519100 682800
rect 519300 682600 519500 682800
rect 519700 682600 519900 682800
rect 520100 682600 520300 682800
rect 520500 682600 520700 682800
rect 36800 681900 37000 682100
rect 37200 681900 37400 682100
rect 37600 681900 37800 682100
rect 38000 681900 38200 682100
rect 58000 682000 58200 682200
rect 58400 682000 58600 682200
rect 58800 682000 59000 682200
rect 59200 682000 59400 682200
rect 59600 682000 59800 682200
rect 60000 682000 60200 682200
rect 60400 682000 60600 682200
rect 60800 682000 61000 682200
rect 61200 682000 61400 682200
rect 61600 682000 61800 682200
rect 36800 681500 37000 681700
rect 37200 681500 37400 681700
rect 37600 681500 37800 681700
rect 38000 681500 38200 681700
rect 36800 681100 37000 681300
rect 37200 681100 37400 681300
rect 37600 681100 37800 681300
rect 38000 681100 38200 681300
rect 36800 680700 37000 680900
rect 37200 680700 37400 680900
rect 37600 680700 37800 680900
rect 38000 680700 38200 680900
rect 549800 681200 550000 681400
rect 550200 681200 550400 681400
rect 550600 681200 550800 681400
rect 551000 681200 551200 681400
rect 551400 681200 551600 681400
rect 551800 681200 552000 681400
rect 552200 681200 552400 681400
rect 552600 681200 552800 681400
rect 549800 680800 550000 681000
rect 550200 680800 550400 681000
rect 550600 680800 550800 681000
rect 551000 680800 551200 681000
rect 551400 680800 551600 681000
rect 551800 680800 552000 681000
rect 552200 680800 552400 681000
rect 552600 680800 552800 681000
rect 36800 680300 37000 680500
rect 37200 680300 37400 680500
rect 37600 680300 37800 680500
rect 38000 680300 38200 680500
rect 515900 679000 516100 679200
rect 516300 679000 516500 679200
rect 516700 679000 516900 679200
rect 517100 679000 517300 679200
rect 517500 679000 517700 679200
rect 517900 679000 518100 679200
rect 518300 679000 518500 679200
rect 518700 679000 518900 679200
rect 519100 679000 519300 679200
rect 519500 679000 519700 679200
rect 519900 679000 520100 679200
rect 520300 679000 520500 679200
rect 520700 679000 520900 679200
rect 515900 678600 516100 678800
rect 516300 678600 516500 678800
rect 516700 678600 516900 678800
rect 517100 678600 517300 678800
rect 517500 678600 517700 678800
rect 517900 678600 518100 678800
rect 518300 678600 518500 678800
rect 518700 678600 518900 678800
rect 519100 678600 519300 678800
rect 519500 678600 519700 678800
rect 519900 678600 520100 678800
rect 520300 678600 520500 678800
rect 520700 678600 520900 678800
rect 515900 678200 516100 678400
rect 516300 678200 516500 678400
rect 516700 678200 516900 678400
rect 517100 678200 517300 678400
rect 517500 678200 517700 678400
rect 517900 678200 518100 678400
rect 518300 678200 518500 678400
rect 518700 678200 518900 678400
rect 519100 678200 519300 678400
rect 519500 678200 519700 678400
rect 519900 678200 520100 678400
rect 520300 678200 520500 678400
rect 520700 678200 520900 678400
rect 515900 677800 516100 678000
rect 516300 677800 516500 678000
rect 516700 677800 516900 678000
rect 517100 677800 517300 678000
rect 517500 677800 517700 678000
rect 517900 677800 518100 678000
rect 518300 677800 518500 678000
rect 518700 677800 518900 678000
rect 519100 677800 519300 678000
rect 519500 677800 519700 678000
rect 519900 677800 520100 678000
rect 520300 677800 520500 678000
rect 520700 677800 520900 678000
rect 515900 677400 516100 677600
rect 516300 677400 516500 677600
rect 516700 677400 516900 677600
rect 517100 677400 517300 677600
rect 517500 677400 517700 677600
rect 517900 677400 518100 677600
rect 518300 677400 518500 677600
rect 518700 677400 518900 677600
rect 519100 677400 519300 677600
rect 519500 677400 519700 677600
rect 519900 677400 520100 677600
rect 520300 677400 520500 677600
rect 520700 677400 520900 677600
rect 515900 677000 516100 677200
rect 516300 677000 516500 677200
rect 516700 677000 516900 677200
rect 517100 677000 517300 677200
rect 517500 677000 517700 677200
rect 517900 677000 518100 677200
rect 518300 677000 518500 677200
rect 518700 677000 518900 677200
rect 519100 677000 519300 677200
rect 519500 677000 519700 677200
rect 519900 677000 520100 677200
rect 520300 677000 520500 677200
rect 520700 677000 520900 677200
rect 515900 676600 516100 676800
rect 516300 676600 516500 676800
rect 516700 676600 516900 676800
rect 517100 676600 517300 676800
rect 517500 676600 517700 676800
rect 517900 676600 518100 676800
rect 518300 676600 518500 676800
rect 518700 676600 518900 676800
rect 519100 676600 519300 676800
rect 519500 676600 519700 676800
rect 519900 676600 520100 676800
rect 520300 676600 520500 676800
rect 520700 676600 520900 676800
rect 32800 663000 33100 663300
rect 33300 663000 33600 663300
rect 33800 663000 34100 663300
rect 34300 663000 34600 663300
rect 34800 663000 35100 663300
rect 35300 663000 35600 663300
rect 35800 663000 36100 663300
rect 36300 663000 36600 663300
rect 36800 663000 37100 663300
rect 37300 663000 37600 663300
rect 37800 663000 38100 663300
rect 38300 663000 38600 663300
rect 38800 663000 39100 663300
rect 39300 663000 39600 663300
rect 39800 663000 40100 663300
rect 40300 663000 40600 663300
rect 2500 648300 2800 648600
rect 3000 648300 3300 648600
rect 3500 648300 3800 648600
rect 2500 647800 2800 648100
rect 3000 647800 3300 648100
rect 3500 647800 3800 648100
rect 2500 647300 2800 647600
rect 3000 647300 3300 647600
rect 3500 647300 3800 647600
rect 2500 646800 2800 647100
rect 3000 646800 3300 647100
rect 3500 646800 3800 647100
rect 2500 646300 2800 646600
rect 3000 646300 3300 646600
rect 3500 646300 3800 646600
rect 2500 645800 2800 646100
rect 3000 645800 3300 646100
rect 3500 645800 3800 646100
rect 2500 645300 2800 645600
rect 3000 645300 3300 645600
rect 3500 645300 3800 645600
rect 2500 644800 2800 645100
rect 3000 644800 3300 645100
rect 3500 644800 3800 645100
rect 2500 644300 2800 644600
rect 3000 644300 3300 644600
rect 3500 644300 3800 644600
rect 2500 643800 2800 644100
rect 3000 643800 3300 644100
rect 3500 643800 3800 644100
rect 2500 643300 2800 643600
rect 3000 643300 3300 643600
rect 3500 643300 3800 643600
rect 2500 642800 2800 643100
rect 3000 642800 3300 643100
rect 3500 642800 3800 643100
rect 2500 642300 2800 642600
rect 3000 642300 3300 642600
rect 3500 642300 3800 642600
rect 2500 641800 2800 642100
rect 3000 641800 3300 642100
rect 3500 641800 3800 642100
rect 2500 641300 2800 641600
rect 3000 641300 3300 641600
rect 3500 641300 3800 641600
rect 2500 640800 2800 641100
rect 3000 640800 3300 641100
rect 3500 640800 3800 641100
rect 2500 640300 2800 640600
rect 3000 640300 3300 640600
rect 3500 640300 3800 640600
rect 2500 639800 2800 640100
rect 3000 639800 3300 640100
rect 3500 639800 3800 640100
rect 2500 639300 2800 639600
rect 3000 639300 3300 639600
rect 3500 639300 3800 639600
rect 2500 638800 2800 639100
rect 3000 638800 3300 639100
rect 3500 638800 3800 639100
rect 2500 638300 2800 638600
rect 3000 638300 3300 638600
rect 3500 638300 3800 638600
rect 2500 637800 2800 638100
rect 3000 637800 3300 638100
rect 3500 637800 3800 638100
rect 2500 637300 2800 637600
rect 3000 637300 3300 637600
rect 3500 637300 3800 637600
rect 2500 636800 2800 637100
rect 3000 636800 3300 637100
rect 3500 636800 3800 637100
rect 2500 636300 2800 636600
rect 3000 636300 3300 636600
rect 3500 636300 3800 636600
rect 2500 635800 2800 636100
rect 3000 635800 3300 636100
rect 3500 635800 3800 636100
rect 2500 635300 2800 635600
rect 3000 635300 3300 635600
rect 3500 635300 3800 635600
rect 2500 634800 2800 635100
rect 3000 634800 3300 635100
rect 3500 634800 3800 635100
rect 2500 634300 2800 634600
rect 3000 634300 3300 634600
rect 3500 634300 3800 634600
rect 550000 644400 550200 644600
rect 550400 644400 550600 644600
rect 550800 644400 551000 644600
rect 551200 644400 551400 644600
rect 551600 644400 551800 644600
rect 552000 644400 552200 644600
rect 552400 644400 552600 644600
rect 552800 644400 553000 644600
rect 550000 644000 550200 644200
rect 550400 644000 550600 644200
rect 550800 644000 551000 644200
rect 551200 644000 551400 644200
rect 551600 644000 551800 644200
rect 552000 644000 552200 644200
rect 552400 644000 552600 644200
rect 552800 644000 553000 644200
rect 550000 643600 550200 643800
rect 550400 643600 550600 643800
rect 550800 643600 551000 643800
rect 551200 643600 551400 643800
rect 551600 643600 551800 643800
rect 552000 643600 552200 643800
rect 552400 643600 552600 643800
rect 552800 643600 553000 643800
rect 550000 643200 550200 643400
rect 550400 643200 550600 643400
rect 550800 643200 551000 643400
rect 551200 643200 551400 643400
rect 551600 643200 551800 643400
rect 552000 643200 552200 643400
rect 552400 643200 552600 643400
rect 552800 643200 553000 643400
rect 550000 642800 550200 643000
rect 550400 642800 550600 643000
rect 550800 642800 551000 643000
rect 551200 642800 551400 643000
rect 551600 642800 551800 643000
rect 552000 642800 552200 643000
rect 552400 642800 552600 643000
rect 552800 642800 553000 643000
rect 550000 642400 550200 642600
rect 550400 642400 550600 642600
rect 550800 642400 551000 642600
rect 551200 642400 551400 642600
rect 551600 642400 551800 642600
rect 552000 642400 552200 642600
rect 552400 642400 552600 642600
rect 552800 642400 553000 642600
rect 550000 642000 550200 642200
rect 550400 642000 550600 642200
rect 550800 642000 551000 642200
rect 551200 642000 551400 642200
rect 551600 642000 551800 642200
rect 552000 642000 552200 642200
rect 552400 642000 552600 642200
rect 552800 642000 553000 642200
rect 550000 641600 550200 641800
rect 550400 641600 550600 641800
rect 550800 641600 551000 641800
rect 551200 641600 551400 641800
rect 551600 641600 551800 641800
rect 552000 641600 552200 641800
rect 552400 641600 552600 641800
rect 552800 641600 553000 641800
rect 550000 641200 550200 641400
rect 550400 641200 550600 641400
rect 550800 641200 551000 641400
rect 551200 641200 551400 641400
rect 551600 641200 551800 641400
rect 552000 641200 552200 641400
rect 552400 641200 552600 641400
rect 552800 641200 553000 641400
rect 550000 640800 550200 641000
rect 550400 640800 550600 641000
rect 550800 640800 551000 641000
rect 551200 640800 551400 641000
rect 551600 640800 551800 641000
rect 552000 640800 552200 641000
rect 552400 640800 552600 641000
rect 552800 640800 553000 641000
rect 550000 640400 550200 640600
rect 550400 640400 550600 640600
rect 550800 640400 551000 640600
rect 551200 640400 551400 640600
rect 551600 640400 551800 640600
rect 552000 640400 552200 640600
rect 552400 640400 552600 640600
rect 552800 640400 553000 640600
rect 550000 640000 550200 640200
rect 550400 640000 550600 640200
rect 550800 640000 551000 640200
rect 551200 640000 551400 640200
rect 551600 640000 551800 640200
rect 552000 640000 552200 640200
rect 552400 640000 552600 640200
rect 552800 640000 553000 640200
rect 550000 639600 550200 639800
rect 550400 639600 550600 639800
rect 550800 639600 551000 639800
rect 551200 639600 551400 639800
rect 551600 639600 551800 639800
rect 552000 639600 552200 639800
rect 552400 639600 552600 639800
rect 552800 639600 553000 639800
rect 550000 639200 550200 639400
rect 550400 639200 550600 639400
rect 550800 639200 551000 639400
rect 551200 639200 551400 639400
rect 551600 639200 551800 639400
rect 552000 639200 552200 639400
rect 552400 639200 552600 639400
rect 552800 639200 553000 639400
rect 550000 638800 550200 639000
rect 550400 638800 550600 639000
rect 550800 638800 551000 639000
rect 551200 638800 551400 639000
rect 551600 638800 551800 639000
rect 552000 638800 552200 639000
rect 552400 638800 552600 639000
rect 552800 638800 553000 639000
rect 550000 638400 550200 638600
rect 550400 638400 550600 638600
rect 550800 638400 551000 638600
rect 551200 638400 551400 638600
rect 551600 638400 551800 638600
rect 552000 638400 552200 638600
rect 552400 638400 552600 638600
rect 552800 638400 553000 638600
rect 550000 638000 550200 638200
rect 550400 638000 550600 638200
rect 550800 638000 551000 638200
rect 551200 638000 551400 638200
rect 551600 638000 551800 638200
rect 552000 638000 552200 638200
rect 552400 638000 552600 638200
rect 552800 638000 553000 638200
rect 550000 637600 550200 637800
rect 550400 637600 550600 637800
rect 550800 637600 551000 637800
rect 551200 637600 551400 637800
rect 551600 637600 551800 637800
rect 552000 637600 552200 637800
rect 552400 637600 552600 637800
rect 552800 637600 553000 637800
rect 550000 637200 550200 637400
rect 550400 637200 550600 637400
rect 550800 637200 551000 637400
rect 551200 637200 551400 637400
rect 551600 637200 551800 637400
rect 552000 637200 552200 637400
rect 552400 637200 552600 637400
rect 552800 637200 553000 637400
rect 550000 636800 550200 637000
rect 550400 636800 550600 637000
rect 550800 636800 551000 637000
rect 551200 636800 551400 637000
rect 551600 636800 551800 637000
rect 552000 636800 552200 637000
rect 552400 636800 552600 637000
rect 552800 636800 553000 637000
rect 550000 636400 550200 636600
rect 550400 636400 550600 636600
rect 550800 636400 551000 636600
rect 551200 636400 551400 636600
rect 551600 636400 551800 636600
rect 552000 636400 552200 636600
rect 552400 636400 552600 636600
rect 552800 636400 553000 636600
rect 550000 636000 550200 636200
rect 550400 636000 550600 636200
rect 550800 636000 551000 636200
rect 551200 636000 551400 636200
rect 551600 636000 551800 636200
rect 552000 636000 552200 636200
rect 552400 636000 552600 636200
rect 552800 636000 553000 636200
rect 550000 635600 550200 635800
rect 550400 635600 550600 635800
rect 550800 635600 551000 635800
rect 551200 635600 551400 635800
rect 551600 635600 551800 635800
rect 552000 635600 552200 635800
rect 552400 635600 552600 635800
rect 552800 635600 553000 635800
rect 550000 635200 550200 635400
rect 550400 635200 550600 635400
rect 550800 635200 551000 635400
rect 551200 635200 551400 635400
rect 551600 635200 551800 635400
rect 552000 635200 552200 635400
rect 552400 635200 552600 635400
rect 552800 635200 553000 635400
rect 550000 634800 550200 635000
rect 550400 634800 550600 635000
rect 550800 634800 551000 635000
rect 551200 634800 551400 635000
rect 551600 634800 551800 635000
rect 552000 634800 552200 635000
rect 552400 634800 552600 635000
rect 552800 634800 553000 635000
rect 550000 634400 550200 634600
rect 550400 634400 550600 634600
rect 550800 634400 551000 634600
rect 551200 634400 551400 634600
rect 551600 634400 551800 634600
rect 552000 634400 552200 634600
rect 552400 634400 552600 634600
rect 552800 634400 553000 634600
rect 550000 634000 550200 634200
rect 550400 634000 550600 634200
rect 550800 634000 551000 634200
rect 551200 634000 551400 634200
rect 551600 634000 551800 634200
rect 552000 634000 552200 634200
rect 552400 634000 552600 634200
rect 552800 634000 553000 634200
rect 550000 633600 550200 633800
rect 550400 633600 550600 633800
rect 550800 633600 551000 633800
rect 551200 633600 551400 633800
rect 551600 633600 551800 633800
rect 552000 633600 552200 633800
rect 552400 633600 552600 633800
rect 552800 633600 553000 633800
rect 550000 633200 550200 633400
rect 550400 633200 550600 633400
rect 550800 633200 551000 633400
rect 551200 633200 551400 633400
rect 551600 633200 551800 633400
rect 552000 633200 552200 633400
rect 552400 633200 552600 633400
rect 552800 633200 553000 633400
rect 550000 632800 550200 633000
rect 550400 632800 550600 633000
rect 550800 632800 551000 633000
rect 551200 632800 551400 633000
rect 551600 632800 551800 633000
rect 552000 632800 552200 633000
rect 552400 632800 552600 633000
rect 552800 632800 553000 633000
rect 550000 632400 550200 632600
rect 550400 632400 550600 632600
rect 550800 632400 551000 632600
rect 551200 632400 551400 632600
rect 551600 632400 551800 632600
rect 552000 632400 552200 632600
rect 552400 632400 552600 632600
rect 552800 632400 553000 632600
rect 550000 632000 550200 632200
rect 550400 632000 550600 632200
rect 550800 632000 551000 632200
rect 551200 632000 551400 632200
rect 551600 632000 551800 632200
rect 552000 632000 552200 632200
rect 552400 632000 552600 632200
rect 552800 632000 553000 632200
rect 550000 631600 550200 631800
rect 550400 631600 550600 631800
rect 550800 631600 551000 631800
rect 551200 631600 551400 631800
rect 551600 631600 551800 631800
rect 552000 631600 552200 631800
rect 552400 631600 552600 631800
rect 552800 631600 553000 631800
rect 550000 631200 550200 631400
rect 550400 631200 550600 631400
rect 550800 631200 551000 631400
rect 551200 631200 551400 631400
rect 551600 631200 551800 631400
rect 552000 631200 552200 631400
rect 552400 631200 552600 631400
rect 552800 631200 553000 631400
rect 550000 630800 550200 631000
rect 550400 630800 550600 631000
rect 550800 630800 551000 631000
rect 551200 630800 551400 631000
rect 551600 630800 551800 631000
rect 552000 630800 552200 631000
rect 552400 630800 552600 631000
rect 552800 630800 553000 631000
rect 550000 630500 550200 630700
rect 550400 630500 550600 630700
rect 550800 630500 551000 630700
rect 551200 630500 551400 630700
rect 551600 630500 551800 630700
rect 552000 630500 552200 630700
rect 552400 630500 552600 630700
rect 552800 630500 553000 630700
rect 550000 630200 550200 630400
rect 550400 630200 550600 630400
rect 550800 630200 551000 630400
rect 551200 630200 551400 630400
rect 551600 630200 551800 630400
rect 552000 630200 552200 630400
rect 552400 630200 552600 630400
rect 552800 630200 553000 630400
rect 550000 629800 550200 630000
rect 550400 629800 550600 630000
rect 550800 629800 551000 630000
rect 551200 629800 551400 630000
rect 551600 629800 551800 630000
rect 552000 629800 552200 630000
rect 552400 629800 552600 630000
rect 552800 629800 553000 630000
rect 32800 563900 33000 564100
rect 33200 563900 33400 564100
rect 33600 563900 33800 564100
rect 34000 563900 34200 564100
rect 34400 563900 34600 564100
rect 34800 563900 35000 564100
rect 35200 563900 35400 564100
rect 35600 563900 35800 564100
rect 36000 563900 36200 564100
rect 36400 563900 36600 564100
rect 36800 563900 37000 564100
rect 37200 563900 37400 564100
rect 37600 563900 37800 564100
rect 38000 563900 38200 564100
rect 38400 563900 38600 564100
rect 38800 563900 39000 564100
rect 39200 563900 39400 564100
rect 39600 563900 39800 564100
rect 40000 563900 40200 564100
rect 40400 563900 40600 564100
rect 32800 563500 33000 563700
rect 33200 563500 33400 563700
rect 33600 563500 33800 563700
rect 34000 563500 34200 563700
rect 34400 563500 34600 563700
rect 34800 563500 35000 563700
rect 35200 563500 35400 563700
rect 35600 563500 35800 563700
rect 36000 563500 36200 563700
rect 36400 563500 36600 563700
rect 36800 563500 37000 563700
rect 37200 563500 37400 563700
rect 37600 563500 37800 563700
rect 38000 563500 38200 563700
rect 38400 563500 38600 563700
rect 38800 563500 39000 563700
rect 39200 563500 39400 563700
rect 39600 563500 39800 563700
rect 40000 563500 40200 563700
rect 40400 563500 40600 563700
rect 32800 563100 33000 563300
rect 33200 563100 33400 563300
rect 33600 563100 33800 563300
rect 34000 563100 34200 563300
rect 34400 563100 34600 563300
rect 34800 563100 35000 563300
rect 35200 563100 35400 563300
rect 35600 563100 35800 563300
rect 36000 563100 36200 563300
rect 36400 563100 36600 563300
rect 36800 563100 37000 563300
rect 37200 563100 37400 563300
rect 37600 563100 37800 563300
rect 38000 563100 38200 563300
rect 38400 563100 38600 563300
rect 38800 563100 39000 563300
rect 39200 563100 39400 563300
rect 39600 563100 39800 563300
rect 40000 563100 40200 563300
rect 40400 563100 40600 563300
rect 32800 562700 33000 562900
rect 33200 562700 33400 562900
rect 33600 562700 33800 562900
rect 34000 562700 34200 562900
rect 34400 562700 34600 562900
rect 34800 562700 35000 562900
rect 35200 562700 35400 562900
rect 35600 562700 35800 562900
rect 36000 562700 36200 562900
rect 36400 562700 36600 562900
rect 36800 562700 37000 562900
rect 37200 562700 37400 562900
rect 37600 562700 37800 562900
rect 38000 562700 38200 562900
rect 38400 562700 38600 562900
rect 38800 562700 39000 562900
rect 39200 562700 39400 562900
rect 39600 562700 39800 562900
rect 40000 562700 40200 562900
rect 40400 562700 40600 562900
rect 32800 562300 33000 562500
rect 33200 562300 33400 562500
rect 33600 562300 33800 562500
rect 34000 562300 34200 562500
rect 34400 562300 34600 562500
rect 34800 562300 35000 562500
rect 35200 562300 35400 562500
rect 35600 562300 35800 562500
rect 36000 562300 36200 562500
rect 36400 562300 36600 562500
rect 36800 562300 37000 562500
rect 37200 562300 37400 562500
rect 37600 562300 37800 562500
rect 38000 562300 38200 562500
rect 38400 562300 38600 562500
rect 38800 562300 39000 562500
rect 39200 562300 39400 562500
rect 39600 562300 39800 562500
rect 40000 562300 40200 562500
rect 40400 562300 40600 562500
rect 32800 561900 33000 562100
rect 33200 561900 33400 562100
rect 33600 561900 33800 562100
rect 34000 561900 34200 562100
rect 34400 561900 34600 562100
rect 34800 561900 35000 562100
rect 35200 561900 35400 562100
rect 35600 561900 35800 562100
rect 36000 561900 36200 562100
rect 36400 561900 36600 562100
rect 36800 561900 37000 562100
rect 37200 561900 37400 562100
rect 37600 561900 37800 562100
rect 38000 561900 38200 562100
rect 38400 561900 38600 562100
rect 38800 561900 39000 562100
rect 39200 561900 39400 562100
rect 39600 561900 39800 562100
rect 40000 561900 40200 562100
rect 40400 561900 40600 562100
rect 32800 561500 33000 561700
rect 33200 561500 33400 561700
rect 33600 561500 33800 561700
rect 34000 561500 34200 561700
rect 34400 561500 34600 561700
rect 34800 561500 35000 561700
rect 35200 561500 35400 561700
rect 35600 561500 35800 561700
rect 36000 561500 36200 561700
rect 36400 561500 36600 561700
rect 36800 561500 37000 561700
rect 37200 561500 37400 561700
rect 37600 561500 37800 561700
rect 38000 561500 38200 561700
rect 38400 561500 38600 561700
rect 38800 561500 39000 561700
rect 39200 561500 39400 561700
rect 39600 561500 39800 561700
rect 40000 561500 40200 561700
rect 40400 561500 40600 561700
rect 32800 561100 33000 561300
rect 33200 561100 33400 561300
rect 33600 561100 33800 561300
rect 34000 561100 34200 561300
rect 34400 561100 34600 561300
rect 34800 561100 35000 561300
rect 35200 561100 35400 561300
rect 35600 561100 35800 561300
rect 36000 561100 36200 561300
rect 36400 561100 36600 561300
rect 36800 561100 37000 561300
rect 37200 561100 37400 561300
rect 37600 561100 37800 561300
rect 38000 561100 38200 561300
rect 38400 561100 38600 561300
rect 38800 561100 39000 561300
rect 39200 561100 39400 561300
rect 39600 561100 39800 561300
rect 40000 561100 40200 561300
rect 40400 561100 40600 561300
rect 32800 560700 33000 560900
rect 33200 560700 33400 560900
rect 33600 560700 33800 560900
rect 34000 560700 34200 560900
rect 34400 560700 34600 560900
rect 34800 560700 35000 560900
rect 35200 560700 35400 560900
rect 35600 560700 35800 560900
rect 36000 560700 36200 560900
rect 36400 560700 36600 560900
rect 36800 560700 37000 560900
rect 37200 560700 37400 560900
rect 37600 560700 37800 560900
rect 38000 560700 38200 560900
rect 38400 560700 38600 560900
rect 38800 560700 39000 560900
rect 39200 560700 39400 560900
rect 39600 560700 39800 560900
rect 40000 560700 40200 560900
rect 40400 560700 40600 560900
rect 32800 560300 33000 560500
rect 33200 560300 33400 560500
rect 33600 560300 33800 560500
rect 34000 560300 34200 560500
rect 34400 560300 34600 560500
rect 34800 560300 35000 560500
rect 35200 560300 35400 560500
rect 35600 560300 35800 560500
rect 36000 560300 36200 560500
rect 36400 560300 36600 560500
rect 36800 560300 37000 560500
rect 37200 560300 37400 560500
rect 37600 560300 37800 560500
rect 38000 560300 38200 560500
rect 38400 560300 38600 560500
rect 38800 560300 39000 560500
rect 39200 560300 39400 560500
rect 39600 560300 39800 560500
rect 40000 560300 40200 560500
rect 40400 560300 40600 560500
rect 32800 559900 33000 560100
rect 33200 559900 33400 560100
rect 33600 559900 33800 560100
rect 34000 559900 34200 560100
rect 34400 559900 34600 560100
rect 34800 559900 35000 560100
rect 35200 559900 35400 560100
rect 35600 559900 35800 560100
rect 36000 559900 36200 560100
rect 36400 559900 36600 560100
rect 36800 559900 37000 560100
rect 37200 559900 37400 560100
rect 37600 559900 37800 560100
rect 38000 559900 38200 560100
rect 38400 559900 38600 560100
rect 38800 559900 39000 560100
rect 39200 559900 39400 560100
rect 39600 559900 39800 560100
rect 40000 559900 40200 560100
rect 40400 559900 40600 560100
rect 32800 559500 33000 559700
rect 33200 559500 33400 559700
rect 33600 559500 33800 559700
rect 34000 559500 34200 559700
rect 34400 559500 34600 559700
rect 34800 559500 35000 559700
rect 35200 559500 35400 559700
rect 35600 559500 35800 559700
rect 36000 559500 36200 559700
rect 36400 559500 36600 559700
rect 36800 559500 37000 559700
rect 37200 559500 37400 559700
rect 37600 559500 37800 559700
rect 38000 559500 38200 559700
rect 38400 559500 38600 559700
rect 38800 559500 39000 559700
rect 39200 559500 39400 559700
rect 39600 559500 39800 559700
rect 40000 559500 40200 559700
rect 40400 559500 40600 559700
rect 32800 559100 33000 559300
rect 33200 559100 33400 559300
rect 33600 559100 33800 559300
rect 34000 559100 34200 559300
rect 34400 559100 34600 559300
rect 34800 559100 35000 559300
rect 35200 559100 35400 559300
rect 35600 559100 35800 559300
rect 36000 559100 36200 559300
rect 36400 559100 36600 559300
rect 36800 559100 37000 559300
rect 37200 559100 37400 559300
rect 37600 559100 37800 559300
rect 38000 559100 38200 559300
rect 38400 559100 38600 559300
rect 38800 559100 39000 559300
rect 39200 559100 39400 559300
rect 39600 559100 39800 559300
rect 40000 559100 40200 559300
rect 40400 559100 40600 559300
rect 32800 558700 33000 558900
rect 33200 558700 33400 558900
rect 33600 558700 33800 558900
rect 34000 558700 34200 558900
rect 34400 558700 34600 558900
rect 34800 558700 35000 558900
rect 35200 558700 35400 558900
rect 35600 558700 35800 558900
rect 36000 558700 36200 558900
rect 36400 558700 36600 558900
rect 36800 558700 37000 558900
rect 37200 558700 37400 558900
rect 37600 558700 37800 558900
rect 38000 558700 38200 558900
rect 38400 558700 38600 558900
rect 38800 558700 39000 558900
rect 39200 558700 39400 558900
rect 39600 558700 39800 558900
rect 40000 558700 40200 558900
rect 40400 558700 40600 558900
rect 32800 558300 33000 558500
rect 33200 558300 33400 558500
rect 33600 558300 33800 558500
rect 34000 558300 34200 558500
rect 34400 558300 34600 558500
rect 34800 558300 35000 558500
rect 35200 558300 35400 558500
rect 35600 558300 35800 558500
rect 36000 558300 36200 558500
rect 36400 558300 36600 558500
rect 36800 558300 37000 558500
rect 37200 558300 37400 558500
rect 37600 558300 37800 558500
rect 38000 558300 38200 558500
rect 38400 558300 38600 558500
rect 38800 558300 39000 558500
rect 39200 558300 39400 558500
rect 39600 558300 39800 558500
rect 40000 558300 40200 558500
rect 40400 558300 40600 558500
rect 32800 557900 33000 558100
rect 33200 557900 33400 558100
rect 33600 557900 33800 558100
rect 34000 557900 34200 558100
rect 34400 557900 34600 558100
rect 34800 557900 35000 558100
rect 35200 557900 35400 558100
rect 35600 557900 35800 558100
rect 36000 557900 36200 558100
rect 36400 557900 36600 558100
rect 36800 557900 37000 558100
rect 37200 557900 37400 558100
rect 37600 557900 37800 558100
rect 38000 557900 38200 558100
rect 38400 557900 38600 558100
rect 38800 557900 39000 558100
rect 39200 557900 39400 558100
rect 39600 557900 39800 558100
rect 40000 557900 40200 558100
rect 40400 557900 40600 558100
rect 32800 557500 33000 557700
rect 33200 557500 33400 557700
rect 33600 557500 33800 557700
rect 34000 557500 34200 557700
rect 34400 557500 34600 557700
rect 34800 557500 35000 557700
rect 35200 557500 35400 557700
rect 35600 557500 35800 557700
rect 36000 557500 36200 557700
rect 36400 557500 36600 557700
rect 36800 557500 37000 557700
rect 37200 557500 37400 557700
rect 37600 557500 37800 557700
rect 38000 557500 38200 557700
rect 38400 557500 38600 557700
rect 38800 557500 39000 557700
rect 39200 557500 39400 557700
rect 39600 557500 39800 557700
rect 40000 557500 40200 557700
rect 40400 557500 40600 557700
rect 32800 557100 33000 557300
rect 33200 557100 33400 557300
rect 33600 557100 33800 557300
rect 34000 557100 34200 557300
rect 34400 557100 34600 557300
rect 34800 557100 35000 557300
rect 35200 557100 35400 557300
rect 35600 557100 35800 557300
rect 36000 557100 36200 557300
rect 36400 557100 36600 557300
rect 36800 557100 37000 557300
rect 37200 557100 37400 557300
rect 37600 557100 37800 557300
rect 38000 557100 38200 557300
rect 38400 557100 38600 557300
rect 38800 557100 39000 557300
rect 39200 557100 39400 557300
rect 39600 557100 39800 557300
rect 40000 557100 40200 557300
rect 40400 557100 40600 557300
rect 32800 556700 33000 556900
rect 33200 556700 33400 556900
rect 33600 556700 33800 556900
rect 34000 556700 34200 556900
rect 34400 556700 34600 556900
rect 34800 556700 35000 556900
rect 35200 556700 35400 556900
rect 35600 556700 35800 556900
rect 36000 556700 36200 556900
rect 36400 556700 36600 556900
rect 36800 556700 37000 556900
rect 37200 556700 37400 556900
rect 37600 556700 37800 556900
rect 38000 556700 38200 556900
rect 38400 556700 38600 556900
rect 38800 556700 39000 556900
rect 39200 556700 39400 556900
rect 39600 556700 39800 556900
rect 40000 556700 40200 556900
rect 40400 556700 40600 556900
rect 32800 556300 33000 556500
rect 33200 556300 33400 556500
rect 33600 556300 33800 556500
rect 34000 556300 34200 556500
rect 34400 556300 34600 556500
rect 34800 556300 35000 556500
rect 35200 556300 35400 556500
rect 35600 556300 35800 556500
rect 36000 556300 36200 556500
rect 36400 556300 36600 556500
rect 36800 556300 37000 556500
rect 37200 556300 37400 556500
rect 37600 556300 37800 556500
rect 38000 556300 38200 556500
rect 38400 556300 38600 556500
rect 38800 556300 39000 556500
rect 39200 556300 39400 556500
rect 39600 556300 39800 556500
rect 40000 556300 40200 556500
rect 40400 556300 40600 556500
rect 32800 555900 33000 556100
rect 33200 555900 33400 556100
rect 33600 555900 33800 556100
rect 34000 555900 34200 556100
rect 34400 555900 34600 556100
rect 34800 555900 35000 556100
rect 35200 555900 35400 556100
rect 35600 555900 35800 556100
rect 36000 555900 36200 556100
rect 36400 555900 36600 556100
rect 36800 555900 37000 556100
rect 37200 555900 37400 556100
rect 37600 555900 37800 556100
rect 38000 555900 38200 556100
rect 38400 555900 38600 556100
rect 38800 555900 39000 556100
rect 39200 555900 39400 556100
rect 39600 555900 39800 556100
rect 40000 555900 40200 556100
rect 40400 555900 40600 556100
rect 32800 555500 33000 555700
rect 33200 555500 33400 555700
rect 33600 555500 33800 555700
rect 34000 555500 34200 555700
rect 34400 555500 34600 555700
rect 34800 555500 35000 555700
rect 35200 555500 35400 555700
rect 35600 555500 35800 555700
rect 36000 555500 36200 555700
rect 36400 555500 36600 555700
rect 36800 555500 37000 555700
rect 37200 555500 37400 555700
rect 37600 555500 37800 555700
rect 38000 555500 38200 555700
rect 38400 555500 38600 555700
rect 38800 555500 39000 555700
rect 39200 555500 39400 555700
rect 39600 555500 39800 555700
rect 40000 555500 40200 555700
rect 40400 555500 40600 555700
rect 32800 555100 33000 555300
rect 33200 555100 33400 555300
rect 33600 555100 33800 555300
rect 34000 555100 34200 555300
rect 34400 555100 34600 555300
rect 34800 555100 35000 555300
rect 35200 555100 35400 555300
rect 35600 555100 35800 555300
rect 36000 555100 36200 555300
rect 36400 555100 36600 555300
rect 36800 555100 37000 555300
rect 37200 555100 37400 555300
rect 37600 555100 37800 555300
rect 38000 555100 38200 555300
rect 38400 555100 38600 555300
rect 38800 555100 39000 555300
rect 39200 555100 39400 555300
rect 39600 555100 39800 555300
rect 40000 555100 40200 555300
rect 40400 555100 40600 555300
rect 32800 554700 33000 554900
rect 33200 554700 33400 554900
rect 33600 554700 33800 554900
rect 34000 554700 34200 554900
rect 34400 554700 34600 554900
rect 34800 554700 35000 554900
rect 35200 554700 35400 554900
rect 35600 554700 35800 554900
rect 36000 554700 36200 554900
rect 36400 554700 36600 554900
rect 36800 554700 37000 554900
rect 37200 554700 37400 554900
rect 37600 554700 37800 554900
rect 38000 554700 38200 554900
rect 38400 554700 38600 554900
rect 38800 554700 39000 554900
rect 39200 554700 39400 554900
rect 39600 554700 39800 554900
rect 40000 554700 40200 554900
rect 40400 554700 40600 554900
rect 32800 554300 33000 554500
rect 33200 554300 33400 554500
rect 33600 554300 33800 554500
rect 34000 554300 34200 554500
rect 34400 554300 34600 554500
rect 34800 554300 35000 554500
rect 35200 554300 35400 554500
rect 35600 554300 35800 554500
rect 36000 554300 36200 554500
rect 36400 554300 36600 554500
rect 36800 554300 37000 554500
rect 37200 554300 37400 554500
rect 37600 554300 37800 554500
rect 38000 554300 38200 554500
rect 38400 554300 38600 554500
rect 38800 554300 39000 554500
rect 39200 554300 39400 554500
rect 39600 554300 39800 554500
rect 40000 554300 40200 554500
rect 40400 554300 40600 554500
rect 32800 553900 33000 554100
rect 33200 553900 33400 554100
rect 33600 553900 33800 554100
rect 34000 553900 34200 554100
rect 34400 553900 34600 554100
rect 34800 553900 35000 554100
rect 35200 553900 35400 554100
rect 35600 553900 35800 554100
rect 36000 553900 36200 554100
rect 36400 553900 36600 554100
rect 36800 553900 37000 554100
rect 37200 553900 37400 554100
rect 37600 553900 37800 554100
rect 38000 553900 38200 554100
rect 38400 553900 38600 554100
rect 38800 553900 39000 554100
rect 39200 553900 39400 554100
rect 39600 553900 39800 554100
rect 40000 553900 40200 554100
rect 40400 553900 40600 554100
rect 32800 553500 33000 553700
rect 33200 553500 33400 553700
rect 33600 553500 33800 553700
rect 34000 553500 34200 553700
rect 34400 553500 34600 553700
rect 34800 553500 35000 553700
rect 35200 553500 35400 553700
rect 35600 553500 35800 553700
rect 36000 553500 36200 553700
rect 36400 553500 36600 553700
rect 36800 553500 37000 553700
rect 37200 553500 37400 553700
rect 37600 553500 37800 553700
rect 38000 553500 38200 553700
rect 38400 553500 38600 553700
rect 38800 553500 39000 553700
rect 39200 553500 39400 553700
rect 39600 553500 39800 553700
rect 40000 553500 40200 553700
rect 40400 553500 40600 553700
rect 32800 553100 33000 553300
rect 33200 553100 33400 553300
rect 33600 553100 33800 553300
rect 34000 553100 34200 553300
rect 34400 553100 34600 553300
rect 34800 553100 35000 553300
rect 35200 553100 35400 553300
rect 35600 553100 35800 553300
rect 36000 553100 36200 553300
rect 36400 553100 36600 553300
rect 36800 553100 37000 553300
rect 37200 553100 37400 553300
rect 37600 553100 37800 553300
rect 38000 553100 38200 553300
rect 38400 553100 38600 553300
rect 38800 553100 39000 553300
rect 39200 553100 39400 553300
rect 39600 553100 39800 553300
rect 40000 553100 40200 553300
rect 40400 553100 40600 553300
rect 32800 552700 33000 552900
rect 33200 552700 33400 552900
rect 33600 552700 33800 552900
rect 34000 552700 34200 552900
rect 34400 552700 34600 552900
rect 34800 552700 35000 552900
rect 35200 552700 35400 552900
rect 35600 552700 35800 552900
rect 36000 552700 36200 552900
rect 36400 552700 36600 552900
rect 36800 552700 37000 552900
rect 37200 552700 37400 552900
rect 37600 552700 37800 552900
rect 38000 552700 38200 552900
rect 38400 552700 38600 552900
rect 38800 552700 39000 552900
rect 39200 552700 39400 552900
rect 39600 552700 39800 552900
rect 40000 552700 40200 552900
rect 40400 552700 40600 552900
rect 32800 552300 33000 552500
rect 33200 552300 33400 552500
rect 33600 552300 33800 552500
rect 34000 552300 34200 552500
rect 34400 552300 34600 552500
rect 34800 552300 35000 552500
rect 35200 552300 35400 552500
rect 35600 552300 35800 552500
rect 36000 552300 36200 552500
rect 36400 552300 36600 552500
rect 36800 552300 37000 552500
rect 37200 552300 37400 552500
rect 37600 552300 37800 552500
rect 38000 552300 38200 552500
rect 38400 552300 38600 552500
rect 38800 552300 39000 552500
rect 39200 552300 39400 552500
rect 39600 552300 39800 552500
rect 40000 552300 40200 552500
rect 40400 552300 40600 552500
rect 32800 551900 33000 552100
rect 33200 551900 33400 552100
rect 33600 551900 33800 552100
rect 34000 551900 34200 552100
rect 34400 551900 34600 552100
rect 34800 551900 35000 552100
rect 35200 551900 35400 552100
rect 35600 551900 35800 552100
rect 36000 551900 36200 552100
rect 36400 551900 36600 552100
rect 36800 551900 37000 552100
rect 37200 551900 37400 552100
rect 37600 551900 37800 552100
rect 38000 551900 38200 552100
rect 38400 551900 38600 552100
rect 38800 551900 39000 552100
rect 39200 551900 39400 552100
rect 39600 551900 39800 552100
rect 40000 551900 40200 552100
rect 40400 551900 40600 552100
rect 32800 551500 33000 551700
rect 33200 551500 33400 551700
rect 33600 551500 33800 551700
rect 34000 551500 34200 551700
rect 34400 551500 34600 551700
rect 34800 551500 35000 551700
rect 35200 551500 35400 551700
rect 35600 551500 35800 551700
rect 36000 551500 36200 551700
rect 36400 551500 36600 551700
rect 36800 551500 37000 551700
rect 37200 551500 37400 551700
rect 37600 551500 37800 551700
rect 38000 551500 38200 551700
rect 38400 551500 38600 551700
rect 38800 551500 39000 551700
rect 39200 551500 39400 551700
rect 39600 551500 39800 551700
rect 40000 551500 40200 551700
rect 40400 551500 40600 551700
rect 32800 551100 33000 551300
rect 33200 551100 33400 551300
rect 33600 551100 33800 551300
rect 34000 551100 34200 551300
rect 34400 551100 34600 551300
rect 34800 551100 35000 551300
rect 35200 551100 35400 551300
rect 35600 551100 35800 551300
rect 36000 551100 36200 551300
rect 36400 551100 36600 551300
rect 36800 551100 37000 551300
rect 37200 551100 37400 551300
rect 37600 551100 37800 551300
rect 38000 551100 38200 551300
rect 38400 551100 38600 551300
rect 38800 551100 39000 551300
rect 39200 551100 39400 551300
rect 39600 551100 39800 551300
rect 40000 551100 40200 551300
rect 40400 551100 40600 551300
rect 32800 550700 33000 550900
rect 33200 550700 33400 550900
rect 33600 550700 33800 550900
rect 34000 550700 34200 550900
rect 34400 550700 34600 550900
rect 34800 550700 35000 550900
rect 35200 550700 35400 550900
rect 35600 550700 35800 550900
rect 36000 550700 36200 550900
rect 36400 550700 36600 550900
rect 36800 550700 37000 550900
rect 37200 550700 37400 550900
rect 37600 550700 37800 550900
rect 38000 550700 38200 550900
rect 38400 550700 38600 550900
rect 38800 550700 39000 550900
rect 39200 550700 39400 550900
rect 39600 550700 39800 550900
rect 40000 550700 40200 550900
rect 40400 550700 40600 550900
rect 32800 550300 33000 550500
rect 33200 550300 33400 550500
rect 33600 550300 33800 550500
rect 34000 550300 34200 550500
rect 34400 550300 34600 550500
rect 34800 550300 35000 550500
rect 35200 550300 35400 550500
rect 35600 550300 35800 550500
rect 36000 550300 36200 550500
rect 36400 550300 36600 550500
rect 36800 550300 37000 550500
rect 37200 550300 37400 550500
rect 37600 550300 37800 550500
rect 38000 550300 38200 550500
rect 38400 550300 38600 550500
rect 38800 550300 39000 550500
rect 39200 550300 39400 550500
rect 39600 550300 39800 550500
rect 40000 550300 40200 550500
rect 40400 550300 40600 550500
rect 32800 549900 33000 550100
rect 33200 549900 33400 550100
rect 33600 549900 33800 550100
rect 34000 549900 34200 550100
rect 34400 549900 34600 550100
rect 34800 549900 35000 550100
rect 35200 549900 35400 550100
rect 35600 549900 35800 550100
rect 36000 549900 36200 550100
rect 36400 549900 36600 550100
rect 36800 549900 37000 550100
rect 37200 549900 37400 550100
rect 37600 549900 37800 550100
rect 38000 549900 38200 550100
rect 38400 549900 38600 550100
rect 38800 549900 39000 550100
rect 39200 549900 39400 550100
rect 39600 549900 39800 550100
rect 40000 549900 40200 550100
rect 40400 549900 40600 550100
rect 32800 549500 33000 549700
rect 33200 549500 33400 549700
rect 33600 549500 33800 549700
rect 34000 549500 34200 549700
rect 34400 549500 34600 549700
rect 34800 549500 35000 549700
rect 35200 549500 35400 549700
rect 35600 549500 35800 549700
rect 36000 549500 36200 549700
rect 36400 549500 36600 549700
rect 36800 549500 37000 549700
rect 37200 549500 37400 549700
rect 37600 549500 37800 549700
rect 38000 549500 38200 549700
rect 38400 549500 38600 549700
rect 38800 549500 39000 549700
rect 39200 549500 39400 549700
rect 39600 549500 39800 549700
rect 40000 549500 40200 549700
rect 40400 549500 40600 549700
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 16200 702200 24340 702300
rect 16200 702000 16400 702200
rect 16600 702000 16800 702200
rect 17000 702000 17200 702200
rect 17400 702000 17600 702200
rect 17800 702000 18000 702200
rect 18200 702000 18400 702200
rect 18600 702000 18800 702200
rect 19000 702000 19200 702200
rect 19400 702000 19600 702200
rect 19800 702000 20000 702200
rect 20200 702000 20400 702200
rect 20600 702000 20800 702200
rect 21000 702180 24340 702200
rect 21000 702060 23400 702180
rect 23520 702060 23600 702180
rect 23720 702060 23800 702180
rect 23920 702060 24000 702180
rect 24120 702060 24200 702180
rect 24320 702060 24340 702180
rect 21000 702000 24340 702060
rect 65040 702260 73200 702300
rect 65040 702080 65060 702260
rect 65240 702080 65400 702260
rect 65580 702080 65740 702260
rect 65920 702200 73200 702260
rect 65920 702080 68400 702200
rect 65040 702040 68400 702080
rect 16200 701940 24340 702000
rect 68200 702000 68400 702040
rect 68600 702000 68800 702200
rect 69000 702000 69200 702200
rect 69400 702000 69600 702200
rect 69800 702000 70000 702200
rect 70200 702000 70400 702200
rect 70600 702000 70800 702200
rect 71000 702000 71200 702200
rect 71400 702000 71600 702200
rect 71800 702000 72000 702200
rect 72200 702000 72400 702200
rect 72600 702000 72800 702200
rect 73000 702000 73200 702200
rect 16200 701800 21200 701940
rect 16200 701600 16400 701800
rect 16600 701600 16800 701800
rect 17000 701600 17200 701800
rect 17400 701600 17600 701800
rect 17800 701600 18000 701800
rect 18200 701600 18400 701800
rect 18600 701600 18800 701800
rect 19000 701600 19200 701800
rect 19400 701600 19600 701800
rect 19800 701600 20000 701800
rect 20200 701600 20400 701800
rect 20600 701600 20800 701800
rect 21000 701600 21200 701800
rect 16200 701400 21200 701600
rect 16200 701200 16400 701400
rect 16600 701200 16800 701400
rect 17000 701200 17200 701400
rect 17400 701200 17600 701400
rect 17800 701200 18000 701400
rect 18200 701200 18400 701400
rect 18600 701200 18800 701400
rect 19000 701200 19200 701400
rect 19400 701200 19600 701400
rect 19800 701200 20000 701400
rect 20200 701200 20400 701400
rect 20600 701200 20800 701400
rect 21000 701200 21200 701400
rect 16200 701000 21200 701200
rect 16200 700800 16400 701000
rect 16600 700800 16800 701000
rect 17000 700800 17200 701000
rect 17400 700800 17600 701000
rect 17800 700800 18000 701000
rect 18200 700800 18400 701000
rect 18600 700800 18800 701000
rect 19000 700800 19200 701000
rect 19400 700800 19600 701000
rect 19800 700800 20000 701000
rect 20200 700800 20400 701000
rect 20600 700800 20800 701000
rect 21000 700800 21200 701000
rect 16200 700600 21200 700800
rect 16200 700400 16400 700600
rect 16600 700400 16800 700600
rect 17000 700400 17200 700600
rect 17400 700400 17600 700600
rect 17800 700400 18000 700600
rect 18200 700400 18400 700600
rect 18600 700400 18800 700600
rect 19000 700400 19200 700600
rect 19400 700400 19600 700600
rect 19800 700400 20000 700600
rect 20200 700400 20400 700600
rect 20600 700400 20800 700600
rect 21000 700400 21200 700600
rect 16200 700200 21200 700400
rect 16200 700000 16400 700200
rect 16600 700000 16800 700200
rect 17000 700000 17200 700200
rect 17400 700000 17600 700200
rect 17800 700000 18000 700200
rect 18200 700000 18400 700200
rect 18600 700000 18800 700200
rect 19000 700000 19200 700200
rect 19400 700000 19600 700200
rect 19800 700000 20000 700200
rect 20200 700000 20400 700200
rect 20600 700000 20800 700200
rect 21000 700000 21200 700200
rect 16200 698400 21200 700000
rect 68200 701800 73200 702000
rect 68200 701600 68400 701800
rect 68600 701600 68800 701800
rect 69000 701600 69200 701800
rect 69400 701600 69600 701800
rect 69800 701600 70000 701800
rect 70200 701600 70400 701800
rect 70600 701600 70800 701800
rect 71000 701600 71200 701800
rect 71400 701600 71600 701800
rect 71800 701600 72000 701800
rect 72200 701600 72400 701800
rect 72600 701600 72800 701800
rect 73000 701600 73200 701800
rect 68200 701400 73200 701600
rect 68200 701200 68400 701400
rect 68600 701200 68800 701400
rect 69000 701200 69200 701400
rect 69400 701200 69600 701400
rect 69800 701200 70000 701400
rect 70200 701200 70400 701400
rect 70600 701200 70800 701400
rect 71000 701200 71200 701400
rect 71400 701200 71600 701400
rect 71800 701200 72000 701400
rect 72200 701200 72400 701400
rect 72600 701200 72800 701400
rect 73000 701200 73200 701400
rect 68200 701000 73200 701200
rect 68200 700800 68400 701000
rect 68600 700800 68800 701000
rect 69000 700800 69200 701000
rect 69400 700800 69600 701000
rect 69800 700800 70000 701000
rect 70200 700800 70400 701000
rect 70600 700800 70800 701000
rect 71000 700800 71200 701000
rect 71400 700800 71600 701000
rect 71800 700800 72000 701000
rect 72200 700800 72400 701000
rect 72600 700800 72800 701000
rect 73000 700800 73200 701000
rect 68200 700600 73200 700800
rect 68200 700400 68400 700600
rect 68600 700400 68800 700600
rect 69000 700400 69200 700600
rect 69400 700400 69600 700600
rect 69800 700400 70000 700600
rect 70200 700400 70400 700600
rect 70600 700400 70800 700600
rect 71000 700400 71200 700600
rect 71400 700400 71600 700600
rect 71800 700400 72000 700600
rect 72200 700400 72400 700600
rect 72600 700400 72800 700600
rect 73000 700400 73200 700600
rect 68200 700200 73200 700400
rect 68200 700000 68400 700200
rect 68600 700000 68800 700200
rect 69000 700000 69200 700200
rect 69400 700000 69600 700200
rect 69800 700000 70000 700200
rect 70200 700000 70400 700200
rect 70600 700000 70800 700200
rect 71000 700000 71200 700200
rect 71400 700000 71600 700200
rect 71800 700000 72000 700200
rect 72200 700000 72400 700200
rect 72600 700000 72800 700200
rect 73000 700000 73200 700200
rect 68200 698400 73200 700000
rect 515500 701600 521000 701800
rect 515500 701400 515700 701600
rect 515900 701400 516100 701600
rect 516300 701400 516500 701600
rect 516700 701400 516900 701600
rect 517100 701400 517300 701600
rect 517500 701400 517700 701600
rect 517900 701400 518100 701600
rect 518300 701400 518500 701600
rect 518700 701400 518900 701600
rect 519100 701400 519300 701600
rect 519500 701400 519700 701600
rect 519900 701400 520100 701600
rect 520300 701400 520500 701600
rect 520700 701400 521000 701600
rect 515500 701200 521000 701400
rect 515500 701000 515700 701200
rect 515900 701000 516100 701200
rect 516300 701000 516500 701200
rect 516700 701000 516900 701200
rect 517100 701000 517300 701200
rect 517500 701000 517700 701200
rect 517900 701000 518100 701200
rect 518300 701000 518500 701200
rect 518700 701000 518900 701200
rect 519100 701000 519300 701200
rect 519500 701000 519700 701200
rect 519900 701000 520100 701200
rect 520300 701000 520500 701200
rect 520700 701000 521000 701200
rect 515500 700800 521000 701000
rect 515500 700600 515700 700800
rect 515900 700600 516100 700800
rect 516300 700600 516500 700800
rect 516700 700600 516900 700800
rect 517100 700600 517300 700800
rect 517500 700600 517700 700800
rect 517900 700600 518100 700800
rect 518300 700600 518500 700800
rect 518700 700600 518900 700800
rect 519100 700600 519300 700800
rect 519500 700600 519700 700800
rect 519900 700600 520100 700800
rect 520300 700600 520500 700800
rect 520700 700600 521000 700800
rect 515500 700400 521000 700600
rect 515500 700200 515700 700400
rect 515900 700200 516100 700400
rect 516300 700200 516500 700400
rect 516700 700200 516900 700400
rect 517100 700200 517300 700400
rect 517500 700200 517700 700400
rect 517900 700200 518100 700400
rect 518300 700200 518500 700400
rect 518700 700200 518900 700400
rect 519100 700200 519300 700400
rect 519500 700200 519700 700400
rect 519900 700200 520100 700400
rect 520300 700200 520500 700400
rect 520700 700200 521000 700400
rect 515500 700000 521000 700200
rect 515500 699800 515700 700000
rect 515900 699800 516100 700000
rect 516300 699800 516500 700000
rect 516700 699800 516900 700000
rect 517100 699800 517300 700000
rect 517500 699800 517700 700000
rect 517900 699800 518100 700000
rect 518300 699800 518500 700000
rect 518700 699800 518900 700000
rect 519100 699800 519300 700000
rect 519500 699800 519700 700000
rect 519900 699800 520100 700000
rect 520300 699800 520500 700000
rect 520700 699800 521000 700000
rect 515500 699600 521000 699800
rect 515500 699400 515700 699600
rect 515900 699400 516100 699600
rect 516300 699400 516500 699600
rect 516700 699400 516900 699600
rect 517100 699400 517300 699600
rect 517500 699400 517700 699600
rect 517900 699400 518100 699600
rect 518300 699400 518500 699600
rect 518700 699400 518900 699600
rect 519100 699400 519300 699600
rect 519500 699400 519700 699600
rect 519900 699400 520100 699600
rect 520300 699400 520500 699600
rect 520700 699400 521000 699600
rect 515500 699200 521000 699400
rect 515500 699000 515700 699200
rect 515900 699000 516100 699200
rect 516300 699000 516500 699200
rect 516700 699000 516900 699200
rect 517100 699000 517300 699200
rect 517500 699000 517700 699200
rect 517900 699000 518100 699200
rect 518300 699000 518500 699200
rect 518700 699000 518900 699200
rect 519100 699000 519300 699200
rect 519500 699000 519700 699200
rect 519900 699000 520100 699200
rect 520300 699000 520500 699200
rect 520700 699000 521000 699200
rect 515500 698500 521000 699000
rect 12800 698200 21200 698400
rect 12800 698000 13000 698200
rect 13200 698000 13600 698200
rect 13800 698000 21200 698200
rect 12800 697800 21200 698000
rect 12800 697600 13000 697800
rect 13200 697600 13600 697800
rect 13800 697600 21200 697800
rect 12800 697200 21200 697600
rect 12800 697000 13000 697200
rect 13200 697000 13600 697200
rect 13800 697000 21200 697200
rect 12800 696800 21200 697000
rect 12800 696600 13000 696800
rect 13200 696600 13600 696800
rect 13800 696600 21200 696800
rect 12800 696400 21200 696600
rect 12800 691900 14120 691980
rect 12800 691700 12900 691900
rect 13100 691700 13200 691900
rect 13400 691700 13500 691900
rect 13700 691700 13800 691900
rect 14000 691700 14120 691900
rect 12800 674100 14120 691700
rect 16200 688700 21200 696400
rect 16200 688500 16400 688700
rect 16600 688500 16800 688700
rect 17000 688500 17200 688700
rect 17400 688500 17600 688700
rect 17800 688500 18000 688700
rect 18200 688500 18400 688700
rect 18600 688500 18800 688700
rect 19000 688500 19200 688700
rect 19400 688500 19600 688700
rect 19800 688500 20000 688700
rect 20200 688500 20400 688700
rect 20600 688500 20800 688700
rect 21000 688500 21200 688700
rect 16200 688300 21200 688500
rect 16200 688100 16400 688300
rect 16600 688100 16800 688300
rect 17000 688100 17200 688300
rect 17400 688100 17600 688300
rect 17800 688100 18000 688300
rect 18200 688100 18400 688300
rect 18600 688100 18800 688300
rect 19000 688100 19200 688300
rect 19400 688100 19600 688300
rect 19800 688100 20000 688300
rect 20200 688100 20400 688300
rect 20600 688100 20800 688300
rect 21000 688100 21200 688300
rect 16200 688000 21200 688100
rect 23200 698200 24600 698400
rect 23200 698000 23400 698200
rect 23600 698000 23800 698200
rect 24000 698000 24200 698200
rect 24400 698000 24600 698200
rect 23200 697800 24600 698000
rect 23200 697600 23400 697800
rect 23600 697600 23800 697800
rect 24000 697600 24200 697800
rect 24400 697600 24600 697800
rect 23200 697400 24600 697600
rect 23200 697200 23400 697400
rect 23600 697200 23800 697400
rect 24000 697200 24200 697400
rect 24400 697200 24600 697400
rect 23200 697000 24600 697200
rect 23200 696800 23400 697000
rect 23600 696800 23800 697000
rect 24000 696800 24200 697000
rect 24400 696800 24600 697000
rect 23200 696600 24600 696800
rect 23200 696400 23400 696600
rect 23600 696400 23800 696600
rect 24000 696400 24200 696600
rect 24400 696400 24600 696600
rect 12800 673800 12900 674100
rect 13200 673800 13700 674100
rect 14000 673800 14120 674100
rect 12800 673600 14120 673800
rect 12800 673300 12900 673600
rect 13200 673300 13700 673600
rect 14000 673300 14120 673600
rect 12800 673100 14120 673300
rect 12800 672800 12900 673100
rect 13200 672800 13700 673100
rect 14000 672800 14120 673100
rect 12800 672700 14120 672800
rect 2499 648600 2801 648601
rect 2499 648300 2500 648600
rect 2800 648300 2801 648600
rect 2499 648299 2801 648300
rect 2999 648600 3301 648601
rect 2999 648300 3000 648600
rect 3300 648300 3301 648600
rect 2999 648299 3301 648300
rect 3499 648600 3801 648601
rect 3499 648300 3500 648600
rect 3800 648300 3801 648600
rect 3499 648299 3801 648300
rect 23200 648500 24600 696400
rect 57800 698200 66000 698400
rect 57800 698000 65000 698200
rect 65200 698000 65600 698200
rect 65800 698000 66000 698200
rect 57800 697800 66000 698000
rect 57800 697600 65000 697800
rect 65200 697600 65600 697800
rect 65800 697600 66000 697800
rect 57800 697400 66000 697600
rect 57800 697200 65000 697400
rect 65200 697200 65600 697400
rect 65800 697200 66000 697400
rect 57800 697000 66000 697200
rect 57800 696800 65000 697000
rect 65200 696800 65600 697000
rect 65800 696800 66000 697000
rect 57800 696600 66000 696800
rect 57800 696400 65000 696600
rect 65200 696400 65600 696600
rect 65800 696400 66000 696600
rect 57800 696200 66000 696400
rect 68200 698200 76400 698400
rect 68200 698000 75400 698200
rect 75600 698000 76000 698200
rect 76200 698000 76400 698200
rect 68200 697800 76400 698000
rect 68200 697600 75400 697800
rect 75600 697600 76000 697800
rect 76200 697600 76400 697800
rect 68200 697400 76400 697600
rect 68200 697200 75400 697400
rect 75600 697200 76000 697400
rect 76200 697200 76400 697400
rect 68200 697000 76400 697200
rect 68200 696800 75400 697000
rect 75600 696800 76000 697000
rect 76200 696800 76400 697000
rect 68200 696600 76400 696800
rect 68200 696400 75400 696600
rect 75600 696400 76000 696600
rect 76200 696400 76400 696600
rect 68200 696200 76400 696400
rect 515500 697400 521000 697940
rect 515500 697200 515700 697400
rect 515900 697200 516100 697400
rect 516300 697200 516500 697400
rect 516700 697200 516900 697400
rect 517100 697200 517300 697400
rect 517500 697200 517700 697400
rect 517900 697200 518100 697400
rect 518300 697200 518500 697400
rect 518700 697200 518900 697400
rect 519100 697200 519300 697400
rect 519500 697200 519700 697400
rect 519900 697200 520100 697400
rect 520300 697200 520500 697400
rect 520700 697200 521000 697400
rect 515500 697000 521000 697200
rect 515500 696800 515700 697000
rect 515900 696800 516100 697000
rect 516300 696800 516500 697000
rect 516700 696800 516900 697000
rect 517100 696800 517300 697000
rect 517500 696800 517700 697000
rect 517900 696800 518100 697000
rect 518300 696800 518500 697000
rect 518700 696800 518900 697000
rect 519100 696800 519300 697000
rect 519500 696800 519700 697000
rect 519900 696800 520100 697000
rect 520300 696800 520500 697000
rect 520700 696800 521000 697000
rect 515500 696600 521000 696800
rect 515500 696400 515700 696600
rect 515900 696400 516100 696600
rect 516300 696400 516500 696600
rect 516700 696400 516900 696600
rect 517100 696400 517300 696600
rect 517500 696400 517700 696600
rect 517900 696400 518100 696600
rect 518300 696400 518500 696600
rect 518700 696400 518900 696600
rect 519100 696400 519300 696600
rect 519500 696400 519700 696600
rect 519900 696400 520100 696600
rect 520300 696400 520500 696600
rect 520700 696400 521000 696600
rect 38699 693000 38861 693001
rect 38699 692840 38700 693000
rect 38860 692840 38861 693000
rect 38699 692839 38861 692840
rect 39119 693000 39281 693001
rect 39119 692840 39120 693000
rect 39280 692840 39281 693000
rect 49959 693000 50101 693001
rect 49959 692860 49960 693000
rect 50100 692860 50101 693000
rect 49959 692859 50101 692860
rect 50179 693000 50321 693001
rect 50179 692860 50180 693000
rect 50320 692860 50321 693000
rect 50179 692859 50321 692860
rect 50399 693000 50541 693001
rect 50399 692860 50400 693000
rect 50540 692860 50541 693000
rect 50399 692859 50541 692860
rect 39119 692839 39281 692840
rect 49959 692800 50101 692801
rect 38699 692780 38861 692781
rect 38699 692620 38700 692780
rect 38860 692620 38861 692780
rect 38699 692619 38861 692620
rect 39119 692780 39281 692781
rect 39119 692620 39120 692780
rect 39280 692620 39281 692780
rect 49959 692660 49960 692800
rect 50100 692660 50101 692800
rect 49959 692659 50101 692660
rect 50179 692800 50321 692801
rect 50179 692660 50180 692800
rect 50320 692660 50321 692800
rect 50179 692659 50321 692660
rect 50399 692800 50541 692801
rect 50399 692660 50400 692800
rect 50540 692660 50541 692800
rect 50399 692659 50541 692660
rect 39119 692619 39281 692620
rect 38699 692560 38861 692561
rect 38699 692400 38700 692560
rect 38860 692400 38861 692560
rect 38699 692399 38861 692400
rect 39119 692560 39281 692561
rect 39119 692400 39120 692560
rect 39280 692400 39281 692560
rect 39119 692399 39281 692400
rect 38699 692340 38861 692341
rect 38699 692180 38700 692340
rect 38860 692180 38861 692340
rect 38699 692179 38861 692180
rect 39119 692340 39281 692341
rect 39119 692180 39120 692340
rect 39280 692180 39281 692340
rect 39119 692179 39281 692180
rect 57800 691900 62200 696200
rect 57800 691700 58000 691900
rect 58200 691700 58400 691900
rect 58600 691700 58800 691900
rect 59000 691700 59200 691900
rect 59400 691700 59600 691900
rect 59800 691700 60000 691900
rect 60200 691700 60400 691900
rect 60600 691700 60800 691900
rect 61000 691700 61200 691900
rect 61400 691700 61600 691900
rect 61800 691700 62200 691900
rect 36600 687300 38400 687400
rect 36600 687100 36800 687300
rect 37000 687100 37200 687300
rect 37400 687100 37600 687300
rect 37800 687100 38000 687300
rect 38200 687100 38400 687300
rect 36600 685300 38400 687100
rect 36600 685100 36800 685300
rect 37000 685100 37200 685300
rect 37400 685100 37600 685300
rect 37800 685100 38000 685300
rect 38200 685100 38400 685300
rect 36600 684900 38400 685100
rect 36600 684700 36800 684900
rect 37000 684700 37200 684900
rect 37400 684700 37600 684900
rect 37800 684700 38000 684900
rect 38200 684700 38400 684900
rect 36600 684500 38400 684700
rect 36600 684300 36800 684500
rect 37000 684300 37200 684500
rect 37400 684300 37600 684500
rect 37800 684300 38000 684500
rect 38200 684300 38400 684500
rect 36600 684100 38400 684300
rect 36600 683900 36800 684100
rect 37000 683900 37200 684100
rect 37400 683900 37600 684100
rect 37800 683900 38000 684100
rect 38200 683900 38400 684100
rect 36600 683700 38400 683900
rect 36600 683500 36800 683700
rect 37000 683500 37200 683700
rect 37400 683500 37600 683700
rect 37800 683500 38000 683700
rect 38200 683500 38400 683700
rect 36600 683300 38400 683500
rect 36600 683100 36800 683300
rect 37000 683100 37200 683300
rect 37400 683100 37600 683300
rect 37800 683100 38000 683300
rect 38200 683100 38400 683300
rect 36600 682900 38400 683100
rect 36600 682700 36800 682900
rect 37000 682700 37200 682900
rect 37400 682700 37600 682900
rect 37800 682700 38000 682900
rect 38200 682700 38400 682900
rect 36600 682500 38400 682700
rect 36600 682300 36800 682500
rect 37000 682300 37200 682500
rect 37400 682300 37600 682500
rect 37800 682300 38000 682500
rect 38200 682300 38400 682500
rect 36600 682100 38400 682300
rect 36600 681900 36800 682100
rect 37000 681900 37200 682100
rect 37400 681900 37600 682100
rect 37800 681900 38000 682100
rect 38200 681900 38400 682100
rect 36600 681700 38400 681900
rect 36600 681500 36800 681700
rect 37000 681500 37200 681700
rect 37400 681500 37600 681700
rect 37800 681500 38000 681700
rect 38200 681500 38400 681700
rect 36600 681300 38400 681500
rect 36600 681100 36800 681300
rect 37000 681100 37200 681300
rect 37400 681100 37600 681300
rect 37800 681100 38000 681300
rect 38200 681100 38400 681300
rect 36600 680900 38400 681100
rect 36600 680700 36800 680900
rect 37000 680700 37200 680900
rect 37400 680700 37600 680900
rect 37800 680700 38000 680900
rect 38200 680700 38400 680900
rect 36600 680500 38400 680700
rect 36600 680300 36800 680500
rect 37000 680300 37200 680500
rect 37400 680300 37600 680500
rect 37800 680300 38000 680500
rect 38200 680300 38400 680500
rect 36600 680200 38400 680300
rect 38670 675000 39330 686050
rect 23200 648200 23400 648500
rect 23700 648200 24100 648500
rect 24400 648200 24600 648500
rect 2499 648100 2801 648101
rect 2499 647800 2500 648100
rect 2800 647800 2801 648100
rect 2499 647799 2801 647800
rect 2999 648100 3301 648101
rect 2999 647800 3000 648100
rect 3300 647800 3301 648100
rect 2999 647799 3301 647800
rect 3499 648100 3801 648101
rect 3499 647800 3500 648100
rect 3800 647800 3801 648100
rect 3499 647799 3801 647800
rect 23200 647900 24600 648200
rect 2499 647600 2801 647601
rect 2499 647300 2500 647600
rect 2800 647300 2801 647600
rect 2499 647299 2801 647300
rect 2999 647600 3301 647601
rect 2999 647300 3000 647600
rect 3300 647300 3301 647600
rect 2999 647299 3301 647300
rect 3499 647600 3801 647601
rect 3499 647300 3500 647600
rect 3800 647300 3801 647600
rect 3499 647299 3801 647300
rect 23200 647600 23400 647900
rect 23700 647600 24100 647900
rect 24400 647600 24600 647900
rect 23200 647300 24600 647600
rect 2499 647100 2801 647101
rect 2499 646800 2500 647100
rect 2800 646800 2801 647100
rect 2499 646799 2801 646800
rect 2999 647100 3301 647101
rect 2999 646800 3000 647100
rect 3300 646800 3301 647100
rect 2999 646799 3301 646800
rect 3499 647100 3801 647101
rect 3499 646800 3500 647100
rect 3800 646800 3801 647100
rect 3499 646799 3801 646800
rect 23200 647000 23400 647300
rect 23700 647000 24100 647300
rect 24400 647000 24600 647300
rect 2499 646600 2801 646601
rect 2499 646300 2500 646600
rect 2800 646300 2801 646600
rect 2499 646299 2801 646300
rect 2999 646600 3301 646601
rect 2999 646300 3000 646600
rect 3300 646300 3301 646600
rect 2999 646299 3301 646300
rect 3499 646600 3801 646601
rect 3499 646300 3500 646600
rect 3800 646300 3801 646600
rect 3499 646299 3801 646300
rect 23200 646600 24600 647000
rect 23200 646300 23400 646600
rect 23700 646300 24100 646600
rect 24400 646300 24600 646600
rect 2499 646100 2801 646101
rect 2499 645800 2500 646100
rect 2800 645800 2801 646100
rect 2499 645799 2801 645800
rect 2999 646100 3301 646101
rect 2999 645800 3000 646100
rect 3300 645800 3301 646100
rect 2999 645799 3301 645800
rect 3499 646100 3801 646101
rect 3499 645800 3500 646100
rect 3800 645800 3801 646100
rect 3499 645799 3801 645800
rect 23200 646000 24600 646300
rect 23200 645700 23400 646000
rect 23700 645700 24100 646000
rect 24400 645700 24600 646000
rect 2499 645600 2801 645601
rect 2499 645300 2500 645600
rect 2800 645300 2801 645600
rect 2499 645299 2801 645300
rect 2999 645600 3301 645601
rect 2999 645300 3000 645600
rect 3300 645300 3301 645600
rect 2999 645299 3301 645300
rect 3499 645600 3801 645601
rect 3499 645300 3500 645600
rect 3800 645300 3801 645600
rect 3499 645299 3801 645300
rect 23200 645400 24600 645700
rect 2499 645100 2801 645101
rect 2499 644800 2500 645100
rect 2800 644800 2801 645100
rect 2499 644799 2801 644800
rect 2999 645100 3301 645101
rect 2999 644800 3000 645100
rect 3300 644800 3301 645100
rect 2999 644799 3301 644800
rect 3499 645100 3801 645101
rect 3499 644800 3500 645100
rect 3800 644800 3801 645100
rect 3499 644799 3801 644800
rect 23200 645100 23400 645400
rect 23700 645100 24100 645400
rect 24400 645100 24600 645400
rect 23200 644800 24600 645100
rect 2499 644600 2801 644601
rect 2499 644300 2500 644600
rect 2800 644300 2801 644600
rect 2499 644299 2801 644300
rect 2999 644600 3301 644601
rect 2999 644300 3000 644600
rect 3300 644300 3301 644600
rect 2999 644299 3301 644300
rect 3499 644600 3801 644601
rect 3499 644300 3500 644600
rect 3800 644300 3801 644600
rect 3499 644299 3801 644300
rect 23200 644500 23400 644800
rect 23700 644500 24100 644800
rect 24400 644500 24600 644800
rect 23200 644200 24600 644500
rect 2499 644100 2801 644101
rect 2499 643800 2500 644100
rect 2800 643800 2801 644100
rect 2499 643799 2801 643800
rect 2999 644100 3301 644101
rect 2999 643800 3000 644100
rect 3300 643800 3301 644100
rect 2999 643799 3301 643800
rect 3499 644100 3801 644101
rect 3499 643800 3500 644100
rect 3800 643800 3801 644100
rect 3499 643799 3801 643800
rect 23200 643900 23400 644200
rect 23700 643900 24100 644200
rect 24400 643900 24600 644200
rect 2499 643600 2801 643601
rect 2499 643300 2500 643600
rect 2800 643300 2801 643600
rect 2499 643299 2801 643300
rect 2999 643600 3301 643601
rect 2999 643300 3000 643600
rect 3300 643300 3301 643600
rect 2999 643299 3301 643300
rect 3499 643600 3801 643601
rect 3499 643300 3500 643600
rect 3800 643300 3801 643600
rect 3499 643299 3801 643300
rect 23200 643600 24600 643900
rect 23200 643300 23400 643600
rect 23700 643300 24100 643600
rect 24400 643300 24600 643600
rect 2499 643100 2801 643101
rect 2499 642800 2500 643100
rect 2800 642800 2801 643100
rect 2499 642799 2801 642800
rect 2999 643100 3301 643101
rect 2999 642800 3000 643100
rect 3300 642800 3301 643100
rect 2999 642799 3301 642800
rect 3499 643100 3801 643101
rect 3499 642800 3500 643100
rect 3800 642800 3801 643100
rect 3499 642799 3801 642800
rect 23200 642900 24600 643300
rect 2499 642600 2801 642601
rect 2499 642300 2500 642600
rect 2800 642300 2801 642600
rect 2499 642299 2801 642300
rect 2999 642600 3301 642601
rect 2999 642300 3000 642600
rect 3300 642300 3301 642600
rect 2999 642299 3301 642300
rect 3499 642600 3801 642601
rect 3499 642300 3500 642600
rect 3800 642300 3801 642600
rect 3499 642299 3801 642300
rect 23200 642600 23400 642900
rect 23700 642600 24100 642900
rect 24400 642600 24600 642900
rect 23200 642300 24600 642600
rect 2499 642100 2801 642101
rect 2499 641800 2500 642100
rect 2800 641800 2801 642100
rect 2499 641799 2801 641800
rect 2999 642100 3301 642101
rect 2999 641800 3000 642100
rect 3300 641800 3301 642100
rect 2999 641799 3301 641800
rect 3499 642100 3801 642101
rect 3499 641800 3500 642100
rect 3800 641800 3801 642100
rect 3499 641799 3801 641800
rect 23200 642000 23400 642300
rect 23700 642000 24100 642300
rect 24400 642000 24600 642300
rect 23200 641700 24600 642000
rect 2499 641600 2801 641601
rect 2499 641300 2500 641600
rect 2800 641300 2801 641600
rect 2499 641299 2801 641300
rect 2999 641600 3301 641601
rect 2999 641300 3000 641600
rect 3300 641300 3301 641600
rect 2999 641299 3301 641300
rect 3499 641600 3801 641601
rect 3499 641300 3500 641600
rect 3800 641300 3801 641600
rect 3499 641299 3801 641300
rect 23200 641400 23400 641700
rect 23700 641400 24100 641700
rect 24400 641400 24600 641700
rect 2499 641100 2801 641101
rect 2499 640800 2500 641100
rect 2800 640800 2801 641100
rect 2499 640799 2801 640800
rect 2999 641100 3301 641101
rect 2999 640800 3000 641100
rect 3300 640800 3301 641100
rect 2999 640799 3301 640800
rect 3499 641100 3801 641101
rect 3499 640800 3500 641100
rect 3800 640800 3801 641100
rect 3499 640799 3801 640800
rect 23200 641100 24600 641400
rect 23200 640800 23400 641100
rect 23700 640800 24100 641100
rect 24400 640800 24600 641100
rect 2499 640600 2801 640601
rect 2499 640300 2500 640600
rect 2800 640300 2801 640600
rect 2499 640299 2801 640300
rect 2999 640600 3301 640601
rect 2999 640300 3000 640600
rect 3300 640300 3301 640600
rect 2999 640299 3301 640300
rect 3499 640600 3801 640601
rect 3499 640300 3500 640600
rect 3800 640300 3801 640600
rect 3499 640299 3801 640300
rect 23200 640500 24600 640800
rect 23200 640200 23400 640500
rect 23700 640200 24100 640500
rect 24400 640200 24600 640500
rect 2499 640100 2801 640101
rect 2499 639800 2500 640100
rect 2800 639800 2801 640100
rect 2499 639799 2801 639800
rect 2999 640100 3301 640101
rect 2999 639800 3000 640100
rect 3300 639800 3301 640100
rect 2999 639799 3301 639800
rect 3499 640100 3801 640101
rect 3499 639800 3500 640100
rect 3800 639800 3801 640100
rect 3499 639799 3801 639800
rect 23200 639900 24600 640200
rect 2499 639600 2801 639601
rect 2499 639300 2500 639600
rect 2800 639300 2801 639600
rect 2499 639299 2801 639300
rect 2999 639600 3301 639601
rect 2999 639300 3000 639600
rect 3300 639300 3301 639600
rect 2999 639299 3301 639300
rect 3499 639600 3801 639601
rect 3499 639300 3500 639600
rect 3800 639300 3801 639600
rect 3499 639299 3801 639300
rect 23200 639600 23400 639900
rect 23700 639600 24100 639900
rect 24400 639600 24600 639900
rect 23200 639300 24600 639600
rect 2499 639100 2801 639101
rect 2499 638800 2500 639100
rect 2800 638800 2801 639100
rect 2499 638799 2801 638800
rect 2999 639100 3301 639101
rect 2999 638800 3000 639100
rect 3300 638800 3301 639100
rect 2999 638799 3301 638800
rect 3499 639100 3801 639101
rect 3499 638800 3500 639100
rect 3800 638800 3801 639100
rect 3499 638799 3801 638800
rect 23200 639000 23400 639300
rect 23700 639000 24100 639300
rect 24400 639000 24600 639300
rect 23200 638700 24600 639000
rect 2499 638600 2801 638601
rect 2499 638300 2500 638600
rect 2800 638300 2801 638600
rect 2499 638299 2801 638300
rect 2999 638600 3301 638601
rect 2999 638300 3000 638600
rect 3300 638300 3301 638600
rect 2999 638299 3301 638300
rect 3499 638600 3801 638601
rect 3499 638300 3500 638600
rect 3800 638300 3801 638600
rect 3499 638299 3801 638300
rect 23200 638400 23400 638700
rect 23700 638400 24100 638700
rect 24400 638400 24600 638700
rect 2499 638100 2801 638101
rect 2499 637800 2500 638100
rect 2800 637800 2801 638100
rect 2499 637799 2801 637800
rect 2999 638100 3301 638101
rect 2999 637800 3000 638100
rect 3300 637800 3301 638100
rect 2999 637799 3301 637800
rect 3499 638100 3801 638101
rect 3499 637800 3500 638100
rect 3800 637800 3801 638100
rect 3499 637799 3801 637800
rect 23200 638100 24600 638400
rect 23200 637800 23400 638100
rect 23700 637800 24100 638100
rect 24400 637800 24600 638100
rect 2499 637600 2801 637601
rect 2499 637300 2500 637600
rect 2800 637300 2801 637600
rect 2499 637299 2801 637300
rect 2999 637600 3301 637601
rect 2999 637300 3000 637600
rect 3300 637300 3301 637600
rect 2999 637299 3301 637300
rect 3499 637600 3801 637601
rect 3499 637300 3500 637600
rect 3800 637300 3801 637600
rect 3499 637299 3801 637300
rect 23200 637400 24600 637800
rect 2499 637100 2801 637101
rect 2499 636800 2500 637100
rect 2800 636800 2801 637100
rect 2499 636799 2801 636800
rect 2999 637100 3301 637101
rect 2999 636800 3000 637100
rect 3300 636800 3301 637100
rect 2999 636799 3301 636800
rect 3499 637100 3801 637101
rect 3499 636800 3500 637100
rect 3800 636800 3801 637100
rect 3499 636799 3801 636800
rect 23200 637100 23400 637400
rect 23700 637100 24100 637400
rect 24400 637100 24600 637400
rect 23200 636700 24600 637100
rect 2499 636600 2801 636601
rect 2499 636300 2500 636600
rect 2800 636300 2801 636600
rect 2499 636299 2801 636300
rect 2999 636600 3301 636601
rect 2999 636300 3000 636600
rect 3300 636300 3301 636600
rect 2999 636299 3301 636300
rect 3499 636600 3801 636601
rect 3499 636300 3500 636600
rect 3800 636300 3801 636600
rect 3499 636299 3801 636300
rect 23200 636400 23400 636700
rect 23700 636400 24100 636700
rect 24400 636400 24600 636700
rect 2499 636100 2801 636101
rect 2499 635800 2500 636100
rect 2800 635800 2801 636100
rect 2499 635799 2801 635800
rect 2999 636100 3301 636101
rect 2999 635800 3000 636100
rect 3300 635800 3301 636100
rect 2999 635799 3301 635800
rect 3499 636100 3801 636101
rect 3499 635800 3500 636100
rect 3800 635800 3801 636100
rect 3499 635799 3801 635800
rect 23200 636000 24600 636400
rect 23200 635700 23400 636000
rect 23700 635700 24100 636000
rect 24400 635700 24600 636000
rect 2499 635600 2801 635601
rect 2499 635300 2500 635600
rect 2800 635300 2801 635600
rect 2499 635299 2801 635300
rect 2999 635600 3301 635601
rect 2999 635300 3000 635600
rect 3300 635300 3301 635600
rect 2999 635299 3301 635300
rect 3499 635600 3801 635601
rect 3499 635300 3500 635600
rect 3800 635300 3801 635600
rect 3499 635299 3801 635300
rect 23200 635200 24600 635700
rect 2499 635100 2801 635101
rect 2499 634800 2500 635100
rect 2800 634800 2801 635100
rect 2499 634799 2801 634800
rect 2999 635100 3301 635101
rect 2999 634800 3000 635100
rect 3300 634800 3301 635100
rect 2999 634799 3301 634800
rect 3499 635100 3801 635101
rect 3499 634800 3500 635100
rect 3800 634800 3801 635100
rect 3499 634799 3801 634800
rect 23200 634900 23400 635200
rect 23700 634900 24100 635200
rect 24400 634900 24600 635200
rect 2499 634600 2801 634601
rect 2499 634300 2500 634600
rect 2800 634300 2801 634600
rect 2499 634299 2801 634300
rect 2999 634600 3301 634601
rect 2999 634300 3000 634600
rect 3300 634300 3301 634600
rect 2999 634299 3301 634300
rect 3499 634600 3801 634601
rect 3499 634300 3500 634600
rect 3800 634300 3801 634600
rect 3499 634299 3801 634300
rect 23200 634500 24600 634900
rect 23200 634200 23400 634500
rect 23700 634200 24100 634500
rect 24400 634200 24600 634500
rect 23200 633800 24600 634200
rect 32600 674000 40800 675000
rect 32600 673700 32800 674000
rect 33100 673700 33300 674000
rect 33600 673700 33800 674000
rect 34100 673700 34300 674000
rect 34600 673700 34800 674000
rect 35100 673700 35300 674000
rect 35600 673700 35800 674000
rect 36100 673700 36300 674000
rect 36600 673700 36800 674000
rect 37100 673700 37300 674000
rect 37600 673700 37800 674000
rect 38100 673700 38300 674000
rect 38600 673700 38800 674000
rect 39100 673700 39300 674000
rect 39600 673700 39800 674000
rect 40100 673700 40300 674000
rect 40600 673700 40800 674000
rect 32600 673200 40800 673700
rect 32600 672900 32800 673200
rect 33100 672900 33300 673200
rect 33600 672900 33800 673200
rect 34100 672900 34300 673200
rect 34600 672900 34800 673200
rect 35100 672900 35300 673200
rect 35600 672900 35800 673200
rect 36100 672900 36300 673200
rect 36600 672900 36800 673200
rect 37100 672900 37300 673200
rect 37600 672900 37800 673200
rect 38100 672900 38300 673200
rect 38600 672900 38800 673200
rect 39100 672900 39300 673200
rect 39600 672900 39800 673200
rect 40100 672900 40300 673200
rect 40600 672900 40800 673200
rect 32600 670700 40800 672900
rect 49920 674000 50580 686100
rect 49920 673700 50100 674000
rect 50400 673700 50580 674000
rect 49920 673600 50580 673700
rect 49920 673300 50100 673600
rect 50400 673300 50580 673600
rect 49920 673200 50580 673300
rect 49920 672900 50100 673200
rect 50400 672900 50580 673200
rect 49920 672700 50580 672900
rect 57800 682200 62200 691700
rect 68200 690200 73200 696200
rect 68200 690000 68400 690200
rect 68600 690000 68800 690200
rect 69000 690000 69200 690200
rect 69400 690000 69600 690200
rect 69800 690000 70000 690200
rect 70200 690000 70400 690200
rect 70600 690000 70800 690200
rect 71000 690000 71200 690200
rect 71400 690000 71600 690200
rect 71800 690000 72000 690200
rect 72200 690000 72400 690200
rect 72600 690000 72800 690200
rect 73000 690000 73200 690200
rect 68200 689800 73200 690000
rect 68200 689600 68400 689800
rect 68600 689600 68800 689800
rect 69000 689600 69200 689800
rect 69400 689600 69600 689800
rect 69800 689600 70000 689800
rect 70200 689600 70400 689800
rect 70600 689600 70800 689800
rect 71000 689600 71200 689800
rect 71400 689600 71600 689800
rect 71800 689600 72000 689800
rect 72200 689600 72400 689800
rect 72600 689600 72800 689800
rect 73000 689600 73200 689800
rect 68200 689400 73200 689600
rect 57800 682000 58000 682200
rect 58200 682000 58400 682200
rect 58600 682000 58800 682200
rect 59000 682000 59200 682200
rect 59400 682000 59600 682200
rect 59800 682000 60000 682200
rect 60200 682000 60400 682200
rect 60600 682000 60800 682200
rect 61000 682000 61200 682200
rect 61400 682000 61600 682200
rect 61800 682000 62200 682200
rect 32600 670400 32800 670700
rect 33100 670400 33300 670700
rect 33600 670400 33800 670700
rect 34100 670400 34300 670700
rect 34600 670400 34800 670700
rect 35100 670400 35300 670700
rect 35600 670400 35800 670700
rect 36100 670400 36300 670700
rect 36600 670400 36800 670700
rect 37100 670400 37300 670700
rect 37600 670400 37800 670700
rect 38100 670400 38300 670700
rect 38600 670400 38800 670700
rect 39100 670400 39300 670700
rect 39600 670400 39800 670700
rect 40100 670400 40300 670700
rect 40600 670400 40800 670700
rect 32600 670000 40800 670400
rect 32600 669700 32800 670000
rect 33100 669700 33300 670000
rect 33600 669700 33800 670000
rect 34100 669700 34300 670000
rect 34600 669700 34800 670000
rect 35100 669700 35300 670000
rect 35600 669700 35800 670000
rect 36100 669700 36300 670000
rect 36600 669700 36800 670000
rect 37100 669700 37300 670000
rect 37600 669700 37800 670000
rect 38100 669700 38300 670000
rect 38600 669700 38800 670000
rect 39100 669700 39300 670000
rect 39600 669700 39800 670000
rect 40100 669700 40300 670000
rect 40600 669700 40800 670000
rect 32600 667400 40800 669700
rect 32600 667100 32800 667400
rect 33100 667100 33300 667400
rect 33600 667100 33800 667400
rect 34100 667100 34300 667400
rect 34600 667100 34800 667400
rect 35100 667100 35300 667400
rect 35600 667100 35800 667400
rect 36100 667100 36300 667400
rect 36600 667100 36800 667400
rect 37100 667100 37300 667400
rect 37600 667100 37800 667400
rect 38100 667100 38300 667400
rect 38600 667100 38800 667400
rect 39100 667100 39300 667400
rect 39600 667100 39800 667400
rect 40100 667100 40300 667400
rect 40600 667100 40800 667400
rect 32600 666700 40800 667100
rect 32600 666400 32800 666700
rect 33100 666400 33300 666700
rect 33600 666400 33800 666700
rect 34100 666400 34300 666700
rect 34600 666400 34800 666700
rect 35100 666400 35300 666700
rect 35600 666400 35800 666700
rect 36100 666400 36300 666700
rect 36600 666400 36800 666700
rect 37100 666400 37300 666700
rect 37600 666400 37800 666700
rect 38100 666400 38300 666700
rect 38600 666400 38800 666700
rect 39100 666400 39300 666700
rect 39600 666400 39800 666700
rect 40100 666400 40300 666700
rect 40600 666400 40800 666700
rect 32600 663300 40800 666400
rect 32600 663000 32800 663300
rect 33100 663000 33300 663300
rect 33600 663000 33800 663300
rect 34100 663000 34300 663300
rect 34600 663000 34800 663300
rect 35100 663000 35300 663300
rect 35600 663000 35800 663300
rect 36100 663000 36300 663300
rect 36600 663000 36800 663300
rect 37100 663000 37300 663300
rect 37600 663000 37800 663300
rect 38100 663000 38300 663300
rect 38600 663000 38800 663300
rect 39100 663000 39300 663300
rect 39600 663000 39800 663300
rect 40100 663000 40300 663300
rect 40600 663000 40800 663300
rect 32600 564100 40800 663000
rect 57800 648600 62200 682000
rect 515500 684800 521000 696400
rect 573100 698000 574220 698200
rect 573100 697800 573300 698000
rect 573500 697800 573800 698000
rect 574000 697800 574220 698000
rect 573100 697600 574220 697800
rect 573100 697400 573300 697600
rect 573500 697400 573800 697600
rect 574000 697400 574220 697600
rect 573100 697200 574220 697400
rect 573100 697000 573300 697200
rect 573500 697000 573800 697200
rect 574000 697000 574220 697200
rect 573100 696800 574220 697000
rect 573100 696600 573300 696800
rect 573500 696600 573800 696800
rect 574000 696600 574220 696800
rect 573100 696400 574220 696600
rect 573100 696200 573300 696400
rect 573500 696200 573800 696400
rect 574000 696200 574220 696400
rect 532200 690400 539200 690500
rect 532200 690200 532300 690400
rect 532500 690200 532700 690400
rect 532900 690200 533100 690400
rect 533300 690200 533500 690400
rect 533700 690200 533900 690400
rect 534100 690200 539200 690400
rect 532200 690100 539200 690200
rect 532200 689900 532300 690100
rect 532500 689900 532700 690100
rect 532900 689900 533100 690100
rect 533300 689900 533500 690100
rect 533700 689900 533900 690100
rect 534100 689900 539200 690100
rect 532200 689700 539200 689900
rect 532200 689500 532300 689700
rect 532500 689500 532700 689700
rect 532900 689500 533100 689700
rect 533300 689500 533500 689700
rect 533700 689500 533900 689700
rect 534100 689500 539200 689700
rect 532200 689300 539200 689500
rect 532200 689100 532300 689300
rect 532500 689100 532700 689300
rect 532900 689100 533100 689300
rect 533300 689100 533500 689300
rect 533700 689100 533900 689300
rect 534100 689100 539200 689300
rect 532200 688900 539200 689100
rect 532200 688700 532300 688900
rect 532500 688700 532700 688900
rect 532900 688700 533100 688900
rect 533300 688700 533500 688900
rect 533700 688700 533900 688900
rect 534100 688700 539200 688900
rect 532200 688600 539200 688700
rect 515500 684600 515700 684800
rect 515900 684600 516100 684800
rect 516300 684600 516500 684800
rect 516700 684600 516900 684800
rect 517100 684600 517300 684800
rect 517500 684600 517700 684800
rect 517900 684600 518100 684800
rect 518300 684600 518500 684800
rect 518700 684600 518900 684800
rect 519100 684600 519300 684800
rect 519500 684600 519700 684800
rect 519900 684600 520100 684800
rect 520300 684600 520500 684800
rect 520700 684600 521000 684800
rect 515500 684400 521000 684600
rect 515500 684200 515700 684400
rect 515900 684200 516100 684400
rect 516300 684200 516500 684400
rect 516700 684200 516900 684400
rect 517100 684200 517300 684400
rect 517500 684200 517700 684400
rect 517900 684200 518100 684400
rect 518300 684200 518500 684400
rect 518700 684200 518900 684400
rect 519100 684200 519300 684400
rect 519500 684200 519700 684400
rect 519900 684200 520100 684400
rect 520300 684200 520500 684400
rect 520700 684200 521000 684400
rect 515500 684000 521000 684200
rect 515500 683800 515700 684000
rect 515900 683800 516100 684000
rect 516300 683800 516500 684000
rect 516700 683800 516900 684000
rect 517100 683800 517300 684000
rect 517500 683800 517700 684000
rect 517900 683800 518100 684000
rect 518300 683800 518500 684000
rect 518700 683800 518900 684000
rect 519100 683800 519300 684000
rect 519500 683800 519700 684000
rect 519900 683800 520100 684000
rect 520300 683800 520500 684000
rect 520700 683800 521000 684000
rect 515500 683600 521000 683800
rect 515500 683400 515700 683600
rect 515900 683400 516100 683600
rect 516300 683400 516500 683600
rect 516700 683400 516900 683600
rect 517100 683400 517300 683600
rect 517500 683400 517700 683600
rect 517900 683400 518100 683600
rect 518300 683400 518500 683600
rect 518700 683400 518900 683600
rect 519100 683400 519300 683600
rect 519500 683400 519700 683600
rect 519900 683400 520100 683600
rect 520300 683400 520500 683600
rect 520700 683400 521000 683600
rect 515500 683200 521000 683400
rect 515500 683000 515700 683200
rect 515900 683000 516100 683200
rect 516300 683000 516500 683200
rect 516700 683000 516900 683200
rect 517100 683000 517300 683200
rect 517500 683000 517700 683200
rect 517900 683000 518100 683200
rect 518300 683000 518500 683200
rect 518700 683000 518900 683200
rect 519100 683000 519300 683200
rect 519500 683000 519700 683200
rect 519900 683000 520100 683200
rect 520300 683000 520500 683200
rect 520700 683000 521000 683200
rect 515500 682800 521000 683000
rect 515500 682600 515700 682800
rect 515900 682600 516100 682800
rect 516300 682600 516500 682800
rect 516700 682600 516900 682800
rect 517100 682600 517300 682800
rect 517500 682600 517700 682800
rect 517900 682600 518100 682800
rect 518300 682600 518500 682800
rect 518700 682600 518900 682800
rect 519100 682600 519300 682800
rect 519500 682600 519700 682800
rect 519900 682600 520100 682800
rect 520300 682600 520500 682800
rect 520700 682600 521000 682800
rect 515500 679200 521000 682600
rect 515500 679000 515900 679200
rect 516100 679000 516300 679200
rect 516500 679000 516700 679200
rect 516900 679000 517100 679200
rect 517300 679000 517500 679200
rect 517700 679000 517900 679200
rect 518100 679000 518300 679200
rect 518500 679000 518700 679200
rect 518900 679000 519100 679200
rect 519300 679000 519500 679200
rect 519700 679000 519900 679200
rect 520100 679000 520300 679200
rect 520500 679000 520700 679200
rect 520900 679000 521000 679200
rect 515500 678800 521000 679000
rect 515500 678600 515900 678800
rect 516100 678600 516300 678800
rect 516500 678600 516700 678800
rect 516900 678600 517100 678800
rect 517300 678600 517500 678800
rect 517700 678600 517900 678800
rect 518100 678600 518300 678800
rect 518500 678600 518700 678800
rect 518900 678600 519100 678800
rect 519300 678600 519500 678800
rect 519700 678600 519900 678800
rect 520100 678600 520300 678800
rect 520500 678600 520700 678800
rect 520900 678600 521000 678800
rect 515500 678400 521000 678600
rect 515500 678200 515900 678400
rect 516100 678200 516300 678400
rect 516500 678200 516700 678400
rect 516900 678200 517100 678400
rect 517300 678200 517500 678400
rect 517700 678200 517900 678400
rect 518100 678200 518300 678400
rect 518500 678200 518700 678400
rect 518900 678200 519100 678400
rect 519300 678200 519500 678400
rect 519700 678200 519900 678400
rect 520100 678200 520300 678400
rect 520500 678200 520700 678400
rect 520900 678200 521000 678400
rect 515500 678000 521000 678200
rect 515500 677800 515900 678000
rect 516100 677800 516300 678000
rect 516500 677800 516700 678000
rect 516900 677800 517100 678000
rect 517300 677800 517500 678000
rect 517700 677800 517900 678000
rect 518100 677800 518300 678000
rect 518500 677800 518700 678000
rect 518900 677800 519100 678000
rect 519300 677800 519500 678000
rect 519700 677800 519900 678000
rect 520100 677800 520300 678000
rect 520500 677800 520700 678000
rect 520900 677800 521000 678000
rect 515500 677600 521000 677800
rect 515500 677400 515900 677600
rect 516100 677400 516300 677600
rect 516500 677400 516700 677600
rect 516900 677400 517100 677600
rect 517300 677400 517500 677600
rect 517700 677400 517900 677600
rect 518100 677400 518300 677600
rect 518500 677400 518700 677600
rect 518900 677400 519100 677600
rect 519300 677400 519500 677600
rect 519700 677400 519900 677600
rect 520100 677400 520300 677600
rect 520500 677400 520700 677600
rect 520900 677400 521000 677600
rect 515500 677200 521000 677400
rect 515500 677000 515900 677200
rect 516100 677000 516300 677200
rect 516500 677000 516700 677200
rect 516900 677000 517100 677200
rect 517300 677000 517500 677200
rect 517700 677000 517900 677200
rect 518100 677000 518300 677200
rect 518500 677000 518700 677200
rect 518900 677000 519100 677200
rect 519300 677000 519500 677200
rect 519700 677000 519900 677200
rect 520100 677000 520300 677200
rect 520500 677000 520700 677200
rect 520900 677000 521000 677200
rect 515500 676800 521000 677000
rect 515500 676600 515900 676800
rect 516100 676600 516300 676800
rect 516500 676600 516700 676800
rect 516900 676600 517100 676800
rect 517300 676600 517500 676800
rect 517700 676600 517900 676800
rect 518100 676600 518300 676800
rect 518500 676600 518700 676800
rect 518900 676600 519100 676800
rect 519300 676600 519500 676800
rect 519700 676600 519900 676800
rect 520100 676600 520300 676800
rect 520500 676600 520700 676800
rect 520900 676600 521000 676800
rect 515500 676460 521000 676600
rect 549700 687300 553100 687400
rect 549700 687200 551200 687300
rect 549700 687000 549900 687200
rect 550100 687000 550200 687200
rect 550400 687000 550500 687200
rect 550700 687000 550800 687200
rect 551000 687100 551200 687200
rect 551400 687100 553100 687300
rect 551000 687000 553100 687100
rect 549700 686800 551200 687000
rect 551400 686800 553100 687000
rect 549700 686700 553100 686800
rect 549700 686500 551200 686700
rect 551400 686500 553100 686700
rect 549700 686400 553100 686500
rect 549700 686200 551200 686400
rect 551400 686200 553100 686400
rect 549700 686100 553100 686200
rect 549700 685900 549800 686100
rect 550000 685900 550100 686100
rect 550300 685900 550400 686100
rect 550600 685900 550800 686100
rect 551000 685900 553100 686100
rect 549700 684900 553100 685900
rect 549700 684600 549900 684900
rect 550200 684600 550400 684900
rect 550700 684600 550900 684900
rect 551200 684600 551400 684900
rect 551700 684600 551900 684900
rect 552200 684600 552400 684900
rect 552700 684600 553100 684900
rect 549700 684400 553100 684600
rect 549700 684100 549900 684400
rect 550200 684100 550400 684400
rect 550700 684100 550900 684400
rect 551200 684100 551400 684400
rect 551700 684100 551900 684400
rect 552200 684100 552400 684400
rect 552700 684100 553100 684400
rect 549700 683900 553100 684100
rect 549700 683600 549900 683900
rect 550200 683600 550400 683900
rect 550700 683600 550900 683900
rect 551200 683600 551400 683900
rect 551700 683600 551900 683900
rect 552200 683600 552400 683900
rect 552700 683600 553100 683900
rect 549700 681400 553100 683600
rect 573100 684900 574220 696200
rect 573100 684600 573200 684900
rect 573500 684600 573800 684900
rect 574100 684600 574220 684900
rect 573100 684400 574220 684600
rect 573100 684100 573200 684400
rect 573500 684100 573800 684400
rect 574100 684100 574220 684400
rect 576799 684700 577101 684701
rect 576799 684400 576800 684700
rect 577100 684400 577101 684700
rect 576799 684399 577101 684400
rect 577299 684700 577601 684701
rect 577299 684400 577300 684700
rect 577600 684400 577601 684700
rect 577299 684399 577601 684400
rect 577799 684700 578101 684701
rect 577799 684400 577800 684700
rect 578100 684400 578101 684700
rect 577799 684399 578101 684400
rect 578299 684700 578601 684701
rect 578299 684400 578300 684700
rect 578600 684400 578601 684700
rect 578299 684399 578601 684400
rect 573100 683900 574220 684100
rect 573100 683600 573200 683900
rect 573500 683600 573800 683900
rect 574100 683600 574220 683900
rect 576799 684200 577101 684201
rect 576799 683900 576800 684200
rect 577100 683900 577101 684200
rect 576799 683899 577101 683900
rect 577299 684200 577601 684201
rect 577299 683900 577300 684200
rect 577600 683900 577601 684200
rect 577299 683899 577601 683900
rect 577799 684200 578101 684201
rect 577799 683900 577800 684200
rect 578100 683900 578101 684200
rect 577799 683899 578101 683900
rect 578299 684200 578601 684201
rect 578299 683900 578300 684200
rect 578600 683900 578601 684200
rect 578299 683899 578601 683900
rect 573100 683400 574220 683600
rect 549700 681200 549800 681400
rect 550000 681200 550200 681400
rect 550400 681200 550600 681400
rect 550800 681200 551000 681400
rect 551200 681200 551400 681400
rect 551600 681200 551800 681400
rect 552000 681200 552200 681400
rect 552400 681200 552600 681400
rect 552800 681200 553100 681400
rect 549700 681000 553100 681200
rect 549700 680800 549800 681000
rect 550000 680800 550200 681000
rect 550400 680800 550600 681000
rect 550800 680800 551000 681000
rect 551200 680800 551400 681000
rect 551600 680800 551800 681000
rect 552000 680800 552200 681000
rect 552400 680800 552600 681000
rect 552800 680800 553100 681000
rect 57800 648300 58000 648600
rect 58300 648300 58500 648600
rect 58800 648300 59000 648600
rect 59300 648300 59500 648600
rect 59800 648300 60000 648600
rect 60300 648300 60500 648600
rect 60800 648300 61000 648600
rect 61300 648300 61500 648600
rect 61800 648300 62200 648600
rect 57800 648100 62200 648300
rect 57800 647800 58000 648100
rect 58300 647800 58500 648100
rect 58800 647800 59000 648100
rect 59300 647800 59500 648100
rect 59800 647800 60000 648100
rect 60300 647800 60500 648100
rect 60800 647800 61000 648100
rect 61300 647800 61500 648100
rect 61800 647800 62200 648100
rect 57800 647600 62200 647800
rect 57800 647300 58000 647600
rect 58300 647300 58500 647600
rect 58800 647300 59000 647600
rect 59300 647300 59500 647600
rect 59800 647300 60000 647600
rect 60300 647300 60500 647600
rect 60800 647300 61000 647600
rect 61300 647300 61500 647600
rect 61800 647300 62200 647600
rect 57800 647100 62200 647300
rect 57800 646800 58000 647100
rect 58300 646800 58500 647100
rect 58800 646800 59000 647100
rect 59300 646800 59500 647100
rect 59800 646800 60000 647100
rect 60300 646800 60500 647100
rect 60800 646800 61000 647100
rect 61300 646800 61500 647100
rect 61800 646800 62200 647100
rect 57800 646600 62200 646800
rect 57800 646300 58000 646600
rect 58300 646300 58500 646600
rect 58800 646300 59000 646600
rect 59300 646300 59500 646600
rect 59800 646300 60000 646600
rect 60300 646300 60500 646600
rect 60800 646300 61000 646600
rect 61300 646300 61500 646600
rect 61800 646300 62200 646600
rect 57800 646100 62200 646300
rect 57800 645800 58000 646100
rect 58300 645800 58500 646100
rect 58800 645800 59000 646100
rect 59300 645800 59500 646100
rect 59800 645800 60000 646100
rect 60300 645800 60500 646100
rect 60800 645800 61000 646100
rect 61300 645800 61500 646100
rect 61800 645800 62200 646100
rect 57800 645600 62200 645800
rect 57800 645300 58000 645600
rect 58300 645300 58500 645600
rect 58800 645300 59000 645600
rect 59300 645300 59500 645600
rect 59800 645300 60000 645600
rect 60300 645300 60500 645600
rect 60800 645300 61000 645600
rect 61300 645300 61500 645600
rect 61800 645300 62200 645600
rect 57800 645100 62200 645300
rect 57800 644800 58000 645100
rect 58300 644800 58500 645100
rect 58800 644800 59000 645100
rect 59300 644800 59500 645100
rect 59800 644800 60000 645100
rect 60300 644800 60500 645100
rect 60800 644800 61000 645100
rect 61300 644800 61500 645100
rect 61800 644800 62200 645100
rect 57800 644600 62200 644800
rect 57800 644300 58000 644600
rect 58300 644300 58500 644600
rect 58800 644300 59000 644600
rect 59300 644300 59500 644600
rect 59800 644300 60000 644600
rect 60300 644300 60500 644600
rect 60800 644300 61000 644600
rect 61300 644300 61500 644600
rect 61800 644300 62200 644600
rect 57800 644100 62200 644300
rect 57800 643800 58000 644100
rect 58300 643800 58500 644100
rect 58800 643800 59000 644100
rect 59300 643800 59500 644100
rect 59800 643800 60000 644100
rect 60300 643800 60500 644100
rect 60800 643800 61000 644100
rect 61300 643800 61500 644100
rect 61800 643800 62200 644100
rect 57800 643600 62200 643800
rect 57800 643300 58000 643600
rect 58300 643300 58500 643600
rect 58800 643300 59000 643600
rect 59300 643300 59500 643600
rect 59800 643300 60000 643600
rect 60300 643300 60500 643600
rect 60800 643300 61000 643600
rect 61300 643300 61500 643600
rect 61800 643300 62200 643600
rect 57800 643100 62200 643300
rect 57800 642800 58000 643100
rect 58300 642800 58500 643100
rect 58800 642800 59000 643100
rect 59300 642800 59500 643100
rect 59800 642800 60000 643100
rect 60300 642800 60500 643100
rect 60800 642800 61000 643100
rect 61300 642800 61500 643100
rect 61800 642800 62200 643100
rect 57800 642600 62200 642800
rect 57800 642300 58000 642600
rect 58300 642300 58500 642600
rect 58800 642300 59000 642600
rect 59300 642300 59500 642600
rect 59800 642300 60000 642600
rect 60300 642300 60500 642600
rect 60800 642300 61000 642600
rect 61300 642300 61500 642600
rect 61800 642300 62200 642600
rect 57800 642100 62200 642300
rect 57800 641800 58000 642100
rect 58300 641800 58500 642100
rect 58800 641800 59000 642100
rect 59300 641800 59500 642100
rect 59800 641800 60000 642100
rect 60300 641800 60500 642100
rect 60800 641800 61000 642100
rect 61300 641800 61500 642100
rect 61800 641800 62200 642100
rect 57800 641600 62200 641800
rect 57800 641300 58000 641600
rect 58300 641300 58500 641600
rect 58800 641300 59000 641600
rect 59300 641300 59500 641600
rect 59800 641300 60000 641600
rect 60300 641300 60500 641600
rect 60800 641300 61000 641600
rect 61300 641300 61500 641600
rect 61800 641300 62200 641600
rect 57800 641100 62200 641300
rect 57800 640800 58000 641100
rect 58300 640800 58500 641100
rect 58800 640800 59000 641100
rect 59300 640800 59500 641100
rect 59800 640800 60000 641100
rect 60300 640800 60500 641100
rect 60800 640800 61000 641100
rect 61300 640800 61500 641100
rect 61800 640800 62200 641100
rect 57800 640600 62200 640800
rect 57800 640300 58000 640600
rect 58300 640300 58500 640600
rect 58800 640300 59000 640600
rect 59300 640300 59500 640600
rect 59800 640300 60000 640600
rect 60300 640300 60500 640600
rect 60800 640300 61000 640600
rect 61300 640300 61500 640600
rect 61800 640300 62200 640600
rect 57800 640100 62200 640300
rect 57800 639800 58000 640100
rect 58300 639800 58500 640100
rect 58800 639800 59000 640100
rect 59300 639800 59500 640100
rect 59800 639800 60000 640100
rect 60300 639800 60500 640100
rect 60800 639800 61000 640100
rect 61300 639800 61500 640100
rect 61800 639800 62200 640100
rect 57800 639600 62200 639800
rect 57800 639300 58000 639600
rect 58300 639300 58500 639600
rect 58800 639300 59000 639600
rect 59300 639300 59500 639600
rect 59800 639300 60000 639600
rect 60300 639300 60500 639600
rect 60800 639300 61000 639600
rect 61300 639300 61500 639600
rect 61800 639300 62200 639600
rect 57800 639100 62200 639300
rect 57800 638800 58000 639100
rect 58300 638800 58500 639100
rect 58800 638800 59000 639100
rect 59300 638800 59500 639100
rect 59800 638800 60000 639100
rect 60300 638800 60500 639100
rect 60800 638800 61000 639100
rect 61300 638800 61500 639100
rect 61800 638800 62200 639100
rect 57800 638600 62200 638800
rect 57800 638300 58000 638600
rect 58300 638300 58500 638600
rect 58800 638300 59000 638600
rect 59300 638300 59500 638600
rect 59800 638300 60000 638600
rect 60300 638300 60500 638600
rect 60800 638300 61000 638600
rect 61300 638300 61500 638600
rect 61800 638300 62200 638600
rect 57800 638100 62200 638300
rect 57800 637800 58000 638100
rect 58300 637800 58500 638100
rect 58800 637800 59000 638100
rect 59300 637800 59500 638100
rect 59800 637800 60000 638100
rect 60300 637800 60500 638100
rect 60800 637800 61000 638100
rect 61300 637800 61500 638100
rect 61800 637800 62200 638100
rect 57800 637600 62200 637800
rect 57800 637300 58000 637600
rect 58300 637300 58500 637600
rect 58800 637300 59000 637600
rect 59300 637300 59500 637600
rect 59800 637300 60000 637600
rect 60300 637300 60500 637600
rect 60800 637300 61000 637600
rect 61300 637300 61500 637600
rect 61800 637300 62200 637600
rect 57800 637100 62200 637300
rect 57800 636800 58000 637100
rect 58300 636800 58500 637100
rect 58800 636800 59000 637100
rect 59300 636800 59500 637100
rect 59800 636800 60000 637100
rect 60300 636800 60500 637100
rect 60800 636800 61000 637100
rect 61300 636800 61500 637100
rect 61800 636800 62200 637100
rect 57800 636600 62200 636800
rect 57800 636300 58000 636600
rect 58300 636300 58500 636600
rect 58800 636300 59000 636600
rect 59300 636300 59500 636600
rect 59800 636300 60000 636600
rect 60300 636300 60500 636600
rect 60800 636300 61000 636600
rect 61300 636300 61500 636600
rect 61800 636300 62200 636600
rect 57800 636100 62200 636300
rect 57800 635800 58000 636100
rect 58300 635800 58500 636100
rect 58800 635800 59000 636100
rect 59300 635800 59500 636100
rect 59800 635800 60000 636100
rect 60300 635800 60500 636100
rect 60800 635800 61000 636100
rect 61300 635800 61500 636100
rect 61800 635800 62200 636100
rect 57800 635600 62200 635800
rect 57800 635300 58000 635600
rect 58300 635300 58500 635600
rect 58800 635300 59000 635600
rect 59300 635300 59500 635600
rect 59800 635300 60000 635600
rect 60300 635300 60500 635600
rect 60800 635300 61000 635600
rect 61300 635300 61500 635600
rect 61800 635300 62200 635600
rect 57800 635100 62200 635300
rect 57800 634800 58000 635100
rect 58300 634800 58500 635100
rect 58800 634800 59000 635100
rect 59300 634800 59500 635100
rect 59800 634800 60000 635100
rect 60300 634800 60500 635100
rect 60800 634800 61000 635100
rect 61300 634800 61500 635100
rect 61800 634800 62200 635100
rect 57800 634600 62200 634800
rect 57800 634300 58000 634600
rect 58300 634300 58500 634600
rect 58800 634300 59000 634600
rect 59300 634300 59500 634600
rect 59800 634300 60000 634600
rect 60300 634300 60500 634600
rect 60800 634300 61000 634600
rect 61300 634300 61500 634600
rect 61800 634300 62200 634600
rect 57800 633800 62200 634300
rect 549700 644600 553100 680800
rect 549700 644400 550000 644600
rect 550200 644400 550400 644600
rect 550600 644400 550800 644600
rect 551000 644400 551200 644600
rect 551400 644400 551600 644600
rect 551800 644400 552000 644600
rect 552200 644400 552400 644600
rect 552600 644400 552800 644600
rect 553000 644400 553100 644600
rect 549700 644200 553100 644400
rect 549700 644000 550000 644200
rect 550200 644000 550400 644200
rect 550600 644000 550800 644200
rect 551000 644000 551200 644200
rect 551400 644000 551600 644200
rect 551800 644000 552000 644200
rect 552200 644000 552400 644200
rect 552600 644000 552800 644200
rect 553000 644000 553100 644200
rect 549700 643800 553100 644000
rect 549700 643600 550000 643800
rect 550200 643600 550400 643800
rect 550600 643600 550800 643800
rect 551000 643600 551200 643800
rect 551400 643600 551600 643800
rect 551800 643600 552000 643800
rect 552200 643600 552400 643800
rect 552600 643600 552800 643800
rect 553000 643600 553100 643800
rect 549700 643400 553100 643600
rect 549700 643200 550000 643400
rect 550200 643200 550400 643400
rect 550600 643200 550800 643400
rect 551000 643200 551200 643400
rect 551400 643200 551600 643400
rect 551800 643200 552000 643400
rect 552200 643200 552400 643400
rect 552600 643200 552800 643400
rect 553000 643200 553100 643400
rect 549700 643000 553100 643200
rect 549700 642800 550000 643000
rect 550200 642800 550400 643000
rect 550600 642800 550800 643000
rect 551000 642800 551200 643000
rect 551400 642800 551600 643000
rect 551800 642800 552000 643000
rect 552200 642800 552400 643000
rect 552600 642800 552800 643000
rect 553000 642800 553100 643000
rect 549700 642600 553100 642800
rect 549700 642400 550000 642600
rect 550200 642400 550400 642600
rect 550600 642400 550800 642600
rect 551000 642400 551200 642600
rect 551400 642400 551600 642600
rect 551800 642400 552000 642600
rect 552200 642400 552400 642600
rect 552600 642400 552800 642600
rect 553000 642400 553100 642600
rect 549700 642200 553100 642400
rect 549700 642000 550000 642200
rect 550200 642000 550400 642200
rect 550600 642000 550800 642200
rect 551000 642000 551200 642200
rect 551400 642000 551600 642200
rect 551800 642000 552000 642200
rect 552200 642000 552400 642200
rect 552600 642000 552800 642200
rect 553000 642000 553100 642200
rect 549700 641800 553100 642000
rect 549700 641600 550000 641800
rect 550200 641600 550400 641800
rect 550600 641600 550800 641800
rect 551000 641600 551200 641800
rect 551400 641600 551600 641800
rect 551800 641600 552000 641800
rect 552200 641600 552400 641800
rect 552600 641600 552800 641800
rect 553000 641600 553100 641800
rect 549700 641400 553100 641600
rect 549700 641200 550000 641400
rect 550200 641200 550400 641400
rect 550600 641200 550800 641400
rect 551000 641200 551200 641400
rect 551400 641200 551600 641400
rect 551800 641200 552000 641400
rect 552200 641200 552400 641400
rect 552600 641200 552800 641400
rect 553000 641200 553100 641400
rect 549700 641000 553100 641200
rect 549700 640800 550000 641000
rect 550200 640800 550400 641000
rect 550600 640800 550800 641000
rect 551000 640800 551200 641000
rect 551400 640800 551600 641000
rect 551800 640800 552000 641000
rect 552200 640800 552400 641000
rect 552600 640800 552800 641000
rect 553000 640800 553100 641000
rect 549700 640600 553100 640800
rect 549700 640400 550000 640600
rect 550200 640400 550400 640600
rect 550600 640400 550800 640600
rect 551000 640400 551200 640600
rect 551400 640400 551600 640600
rect 551800 640400 552000 640600
rect 552200 640400 552400 640600
rect 552600 640400 552800 640600
rect 553000 640400 553100 640600
rect 549700 640200 553100 640400
rect 549700 640000 550000 640200
rect 550200 640000 550400 640200
rect 550600 640000 550800 640200
rect 551000 640000 551200 640200
rect 551400 640000 551600 640200
rect 551800 640000 552000 640200
rect 552200 640000 552400 640200
rect 552600 640000 552800 640200
rect 553000 640000 553100 640200
rect 549700 639800 553100 640000
rect 549700 639600 550000 639800
rect 550200 639600 550400 639800
rect 550600 639600 550800 639800
rect 551000 639600 551200 639800
rect 551400 639600 551600 639800
rect 551800 639600 552000 639800
rect 552200 639600 552400 639800
rect 552600 639600 552800 639800
rect 553000 639600 553100 639800
rect 549700 639400 553100 639600
rect 549700 639200 550000 639400
rect 550200 639200 550400 639400
rect 550600 639200 550800 639400
rect 551000 639200 551200 639400
rect 551400 639200 551600 639400
rect 551800 639200 552000 639400
rect 552200 639200 552400 639400
rect 552600 639200 552800 639400
rect 553000 639200 553100 639400
rect 549700 639000 553100 639200
rect 549700 638800 550000 639000
rect 550200 638800 550400 639000
rect 550600 638800 550800 639000
rect 551000 638800 551200 639000
rect 551400 638800 551600 639000
rect 551800 638800 552000 639000
rect 552200 638800 552400 639000
rect 552600 638800 552800 639000
rect 553000 638800 553100 639000
rect 549700 638600 553100 638800
rect 549700 638400 550000 638600
rect 550200 638400 550400 638600
rect 550600 638400 550800 638600
rect 551000 638400 551200 638600
rect 551400 638400 551600 638600
rect 551800 638400 552000 638600
rect 552200 638400 552400 638600
rect 552600 638400 552800 638600
rect 553000 638400 553100 638600
rect 549700 638200 553100 638400
rect 549700 638000 550000 638200
rect 550200 638000 550400 638200
rect 550600 638000 550800 638200
rect 551000 638000 551200 638200
rect 551400 638000 551600 638200
rect 551800 638000 552000 638200
rect 552200 638000 552400 638200
rect 552600 638000 552800 638200
rect 553000 638000 553100 638200
rect 549700 637800 553100 638000
rect 549700 637600 550000 637800
rect 550200 637600 550400 637800
rect 550600 637600 550800 637800
rect 551000 637600 551200 637800
rect 551400 637600 551600 637800
rect 551800 637600 552000 637800
rect 552200 637600 552400 637800
rect 552600 637600 552800 637800
rect 553000 637600 553100 637800
rect 549700 637400 553100 637600
rect 549700 637200 550000 637400
rect 550200 637200 550400 637400
rect 550600 637200 550800 637400
rect 551000 637200 551200 637400
rect 551400 637200 551600 637400
rect 551800 637200 552000 637400
rect 552200 637200 552400 637400
rect 552600 637200 552800 637400
rect 553000 637200 553100 637400
rect 549700 637000 553100 637200
rect 549700 636800 550000 637000
rect 550200 636800 550400 637000
rect 550600 636800 550800 637000
rect 551000 636800 551200 637000
rect 551400 636800 551600 637000
rect 551800 636800 552000 637000
rect 552200 636800 552400 637000
rect 552600 636800 552800 637000
rect 553000 636800 553100 637000
rect 549700 636600 553100 636800
rect 549700 636400 550000 636600
rect 550200 636400 550400 636600
rect 550600 636400 550800 636600
rect 551000 636400 551200 636600
rect 551400 636400 551600 636600
rect 551800 636400 552000 636600
rect 552200 636400 552400 636600
rect 552600 636400 552800 636600
rect 553000 636400 553100 636600
rect 549700 636200 553100 636400
rect 549700 636000 550000 636200
rect 550200 636000 550400 636200
rect 550600 636000 550800 636200
rect 551000 636000 551200 636200
rect 551400 636000 551600 636200
rect 551800 636000 552000 636200
rect 552200 636000 552400 636200
rect 552600 636000 552800 636200
rect 553000 636000 553100 636200
rect 549700 635800 553100 636000
rect 549700 635600 550000 635800
rect 550200 635600 550400 635800
rect 550600 635600 550800 635800
rect 551000 635600 551200 635800
rect 551400 635600 551600 635800
rect 551800 635600 552000 635800
rect 552200 635600 552400 635800
rect 552600 635600 552800 635800
rect 553000 635600 553100 635800
rect 549700 635400 553100 635600
rect 549700 635200 550000 635400
rect 550200 635200 550400 635400
rect 550600 635200 550800 635400
rect 551000 635200 551200 635400
rect 551400 635200 551600 635400
rect 551800 635200 552000 635400
rect 552200 635200 552400 635400
rect 552600 635200 552800 635400
rect 553000 635200 553100 635400
rect 549700 635000 553100 635200
rect 549700 634800 550000 635000
rect 550200 634800 550400 635000
rect 550600 634800 550800 635000
rect 551000 634800 551200 635000
rect 551400 634800 551600 635000
rect 551800 634800 552000 635000
rect 552200 634800 552400 635000
rect 552600 634800 552800 635000
rect 553000 634800 553100 635000
rect 549700 634600 553100 634800
rect 549700 634400 550000 634600
rect 550200 634400 550400 634600
rect 550600 634400 550800 634600
rect 551000 634400 551200 634600
rect 551400 634400 551600 634600
rect 551800 634400 552000 634600
rect 552200 634400 552400 634600
rect 552600 634400 552800 634600
rect 553000 634400 553100 634600
rect 549700 634200 553100 634400
rect 549700 634000 550000 634200
rect 550200 634000 550400 634200
rect 550600 634000 550800 634200
rect 551000 634000 551200 634200
rect 551400 634000 551600 634200
rect 551800 634000 552000 634200
rect 552200 634000 552400 634200
rect 552600 634000 552800 634200
rect 553000 634000 553100 634200
rect 549700 633800 553100 634000
rect 549700 633600 550000 633800
rect 550200 633600 550400 633800
rect 550600 633600 550800 633800
rect 551000 633600 551200 633800
rect 551400 633600 551600 633800
rect 551800 633600 552000 633800
rect 552200 633600 552400 633800
rect 552600 633600 552800 633800
rect 553000 633600 553100 633800
rect 549700 633400 553100 633600
rect 549700 633200 550000 633400
rect 550200 633200 550400 633400
rect 550600 633200 550800 633400
rect 551000 633200 551200 633400
rect 551400 633200 551600 633400
rect 551800 633200 552000 633400
rect 552200 633200 552400 633400
rect 552600 633200 552800 633400
rect 553000 633200 553100 633400
rect 549700 633000 553100 633200
rect 549700 632800 550000 633000
rect 550200 632800 550400 633000
rect 550600 632800 550800 633000
rect 551000 632800 551200 633000
rect 551400 632800 551600 633000
rect 551800 632800 552000 633000
rect 552200 632800 552400 633000
rect 552600 632800 552800 633000
rect 553000 632800 553100 633000
rect 549700 632600 553100 632800
rect 549700 632400 550000 632600
rect 550200 632400 550400 632600
rect 550600 632400 550800 632600
rect 551000 632400 551200 632600
rect 551400 632400 551600 632600
rect 551800 632400 552000 632600
rect 552200 632400 552400 632600
rect 552600 632400 552800 632600
rect 553000 632400 553100 632600
rect 549700 632200 553100 632400
rect 549700 632000 550000 632200
rect 550200 632000 550400 632200
rect 550600 632000 550800 632200
rect 551000 632000 551200 632200
rect 551400 632000 551600 632200
rect 551800 632000 552000 632200
rect 552200 632000 552400 632200
rect 552600 632000 552800 632200
rect 553000 632000 553100 632200
rect 549700 631800 553100 632000
rect 549700 631600 550000 631800
rect 550200 631600 550400 631800
rect 550600 631600 550800 631800
rect 551000 631600 551200 631800
rect 551400 631600 551600 631800
rect 551800 631600 552000 631800
rect 552200 631600 552400 631800
rect 552600 631600 552800 631800
rect 553000 631600 553100 631800
rect 549700 631400 553100 631600
rect 549700 631200 550000 631400
rect 550200 631200 550400 631400
rect 550600 631200 550800 631400
rect 551000 631200 551200 631400
rect 551400 631200 551600 631400
rect 551800 631200 552000 631400
rect 552200 631200 552400 631400
rect 552600 631200 552800 631400
rect 553000 631200 553100 631400
rect 549700 631000 553100 631200
rect 549700 630800 550000 631000
rect 550200 630800 550400 631000
rect 550600 630800 550800 631000
rect 551000 630800 551200 631000
rect 551400 630800 551600 631000
rect 551800 630800 552000 631000
rect 552200 630800 552400 631000
rect 552600 630800 552800 631000
rect 553000 630800 553100 631000
rect 549700 630700 553100 630800
rect 549700 630500 550000 630700
rect 550200 630500 550400 630700
rect 550600 630500 550800 630700
rect 551000 630500 551200 630700
rect 551400 630500 551600 630700
rect 551800 630500 552000 630700
rect 552200 630500 552400 630700
rect 552600 630500 552800 630700
rect 553000 630500 553100 630700
rect 549700 630400 553100 630500
rect 549700 630200 550000 630400
rect 550200 630200 550400 630400
rect 550600 630200 550800 630400
rect 551000 630200 551200 630400
rect 551400 630200 551600 630400
rect 551800 630200 552000 630400
rect 552200 630200 552400 630400
rect 552600 630200 552800 630400
rect 553000 630200 553100 630400
rect 549700 630000 553100 630200
rect 549700 629800 550000 630000
rect 550200 629800 550400 630000
rect 550600 629800 550800 630000
rect 551000 629800 551200 630000
rect 551400 629800 551600 630000
rect 551800 629800 552000 630000
rect 552200 629800 552400 630000
rect 552600 629800 552800 630000
rect 553000 629800 553100 630000
rect 549700 629700 553100 629800
rect 32600 563900 32800 564100
rect 33000 563900 33200 564100
rect 33400 563900 33600 564100
rect 33800 563900 34000 564100
rect 34200 563900 34400 564100
rect 34600 563900 34800 564100
rect 35000 563900 35200 564100
rect 35400 563900 35600 564100
rect 35800 563900 36000 564100
rect 36200 563900 36400 564100
rect 36600 563900 36800 564100
rect 37000 563900 37200 564100
rect 37400 563900 37600 564100
rect 37800 563900 38000 564100
rect 38200 563900 38400 564100
rect 38600 563900 38800 564100
rect 39000 563900 39200 564100
rect 39400 563900 39600 564100
rect 39800 563900 40000 564100
rect 40200 563900 40400 564100
rect 40600 563900 40800 564100
rect 32600 563700 40800 563900
rect 32600 563500 32800 563700
rect 33000 563500 33200 563700
rect 33400 563500 33600 563700
rect 33800 563500 34000 563700
rect 34200 563500 34400 563700
rect 34600 563500 34800 563700
rect 35000 563500 35200 563700
rect 35400 563500 35600 563700
rect 35800 563500 36000 563700
rect 36200 563500 36400 563700
rect 36600 563500 36800 563700
rect 37000 563500 37200 563700
rect 37400 563500 37600 563700
rect 37800 563500 38000 563700
rect 38200 563500 38400 563700
rect 38600 563500 38800 563700
rect 39000 563500 39200 563700
rect 39400 563500 39600 563700
rect 39800 563500 40000 563700
rect 40200 563500 40400 563700
rect 40600 563500 40800 563700
rect 32600 563300 40800 563500
rect 32600 563100 32800 563300
rect 33000 563100 33200 563300
rect 33400 563100 33600 563300
rect 33800 563100 34000 563300
rect 34200 563100 34400 563300
rect 34600 563100 34800 563300
rect 35000 563100 35200 563300
rect 35400 563100 35600 563300
rect 35800 563100 36000 563300
rect 36200 563100 36400 563300
rect 36600 563100 36800 563300
rect 37000 563100 37200 563300
rect 37400 563100 37600 563300
rect 37800 563100 38000 563300
rect 38200 563100 38400 563300
rect 38600 563100 38800 563300
rect 39000 563100 39200 563300
rect 39400 563100 39600 563300
rect 39800 563100 40000 563300
rect 40200 563100 40400 563300
rect 40600 563100 40800 563300
rect 32600 562900 40800 563100
rect 32600 562700 32800 562900
rect 33000 562700 33200 562900
rect 33400 562700 33600 562900
rect 33800 562700 34000 562900
rect 34200 562700 34400 562900
rect 34600 562700 34800 562900
rect 35000 562700 35200 562900
rect 35400 562700 35600 562900
rect 35800 562700 36000 562900
rect 36200 562700 36400 562900
rect 36600 562700 36800 562900
rect 37000 562700 37200 562900
rect 37400 562700 37600 562900
rect 37800 562700 38000 562900
rect 38200 562700 38400 562900
rect 38600 562700 38800 562900
rect 39000 562700 39200 562900
rect 39400 562700 39600 562900
rect 39800 562700 40000 562900
rect 40200 562700 40400 562900
rect 40600 562700 40800 562900
rect 32600 562500 40800 562700
rect 32600 562300 32800 562500
rect 33000 562300 33200 562500
rect 33400 562300 33600 562500
rect 33800 562300 34000 562500
rect 34200 562300 34400 562500
rect 34600 562300 34800 562500
rect 35000 562300 35200 562500
rect 35400 562300 35600 562500
rect 35800 562300 36000 562500
rect 36200 562300 36400 562500
rect 36600 562300 36800 562500
rect 37000 562300 37200 562500
rect 37400 562300 37600 562500
rect 37800 562300 38000 562500
rect 38200 562300 38400 562500
rect 38600 562300 38800 562500
rect 39000 562300 39200 562500
rect 39400 562300 39600 562500
rect 39800 562300 40000 562500
rect 40200 562300 40400 562500
rect 40600 562300 40800 562500
rect 32600 562100 40800 562300
rect 32600 561900 32800 562100
rect 33000 561900 33200 562100
rect 33400 561900 33600 562100
rect 33800 561900 34000 562100
rect 34200 561900 34400 562100
rect 34600 561900 34800 562100
rect 35000 561900 35200 562100
rect 35400 561900 35600 562100
rect 35800 561900 36000 562100
rect 36200 561900 36400 562100
rect 36600 561900 36800 562100
rect 37000 561900 37200 562100
rect 37400 561900 37600 562100
rect 37800 561900 38000 562100
rect 38200 561900 38400 562100
rect 38600 561900 38800 562100
rect 39000 561900 39200 562100
rect 39400 561900 39600 562100
rect 39800 561900 40000 562100
rect 40200 561900 40400 562100
rect 40600 561900 40800 562100
rect 32600 561700 40800 561900
rect 32600 561500 32800 561700
rect 33000 561500 33200 561700
rect 33400 561500 33600 561700
rect 33800 561500 34000 561700
rect 34200 561500 34400 561700
rect 34600 561500 34800 561700
rect 35000 561500 35200 561700
rect 35400 561500 35600 561700
rect 35800 561500 36000 561700
rect 36200 561500 36400 561700
rect 36600 561500 36800 561700
rect 37000 561500 37200 561700
rect 37400 561500 37600 561700
rect 37800 561500 38000 561700
rect 38200 561500 38400 561700
rect 38600 561500 38800 561700
rect 39000 561500 39200 561700
rect 39400 561500 39600 561700
rect 39800 561500 40000 561700
rect 40200 561500 40400 561700
rect 40600 561500 40800 561700
rect 32600 561300 40800 561500
rect 32600 561100 32800 561300
rect 33000 561100 33200 561300
rect 33400 561100 33600 561300
rect 33800 561100 34000 561300
rect 34200 561100 34400 561300
rect 34600 561100 34800 561300
rect 35000 561100 35200 561300
rect 35400 561100 35600 561300
rect 35800 561100 36000 561300
rect 36200 561100 36400 561300
rect 36600 561100 36800 561300
rect 37000 561100 37200 561300
rect 37400 561100 37600 561300
rect 37800 561100 38000 561300
rect 38200 561100 38400 561300
rect 38600 561100 38800 561300
rect 39000 561100 39200 561300
rect 39400 561100 39600 561300
rect 39800 561100 40000 561300
rect 40200 561100 40400 561300
rect 40600 561100 40800 561300
rect 32600 560900 40800 561100
rect 32600 560700 32800 560900
rect 33000 560700 33200 560900
rect 33400 560700 33600 560900
rect 33800 560700 34000 560900
rect 34200 560700 34400 560900
rect 34600 560700 34800 560900
rect 35000 560700 35200 560900
rect 35400 560700 35600 560900
rect 35800 560700 36000 560900
rect 36200 560700 36400 560900
rect 36600 560700 36800 560900
rect 37000 560700 37200 560900
rect 37400 560700 37600 560900
rect 37800 560700 38000 560900
rect 38200 560700 38400 560900
rect 38600 560700 38800 560900
rect 39000 560700 39200 560900
rect 39400 560700 39600 560900
rect 39800 560700 40000 560900
rect 40200 560700 40400 560900
rect 40600 560700 40800 560900
rect 32600 560500 40800 560700
rect 32600 560300 32800 560500
rect 33000 560300 33200 560500
rect 33400 560300 33600 560500
rect 33800 560300 34000 560500
rect 34200 560300 34400 560500
rect 34600 560300 34800 560500
rect 35000 560300 35200 560500
rect 35400 560300 35600 560500
rect 35800 560300 36000 560500
rect 36200 560300 36400 560500
rect 36600 560300 36800 560500
rect 37000 560300 37200 560500
rect 37400 560300 37600 560500
rect 37800 560300 38000 560500
rect 38200 560300 38400 560500
rect 38600 560300 38800 560500
rect 39000 560300 39200 560500
rect 39400 560300 39600 560500
rect 39800 560300 40000 560500
rect 40200 560300 40400 560500
rect 40600 560300 40800 560500
rect 32600 560100 40800 560300
rect 32600 559900 32800 560100
rect 33000 559900 33200 560100
rect 33400 559900 33600 560100
rect 33800 559900 34000 560100
rect 34200 559900 34400 560100
rect 34600 559900 34800 560100
rect 35000 559900 35200 560100
rect 35400 559900 35600 560100
rect 35800 559900 36000 560100
rect 36200 559900 36400 560100
rect 36600 559900 36800 560100
rect 37000 559900 37200 560100
rect 37400 559900 37600 560100
rect 37800 559900 38000 560100
rect 38200 559900 38400 560100
rect 38600 559900 38800 560100
rect 39000 559900 39200 560100
rect 39400 559900 39600 560100
rect 39800 559900 40000 560100
rect 40200 559900 40400 560100
rect 40600 559900 40800 560100
rect 32600 559700 40800 559900
rect 32600 559500 32800 559700
rect 33000 559500 33200 559700
rect 33400 559500 33600 559700
rect 33800 559500 34000 559700
rect 34200 559500 34400 559700
rect 34600 559500 34800 559700
rect 35000 559500 35200 559700
rect 35400 559500 35600 559700
rect 35800 559500 36000 559700
rect 36200 559500 36400 559700
rect 36600 559500 36800 559700
rect 37000 559500 37200 559700
rect 37400 559500 37600 559700
rect 37800 559500 38000 559700
rect 38200 559500 38400 559700
rect 38600 559500 38800 559700
rect 39000 559500 39200 559700
rect 39400 559500 39600 559700
rect 39800 559500 40000 559700
rect 40200 559500 40400 559700
rect 40600 559500 40800 559700
rect 32600 559300 40800 559500
rect 32600 559100 32800 559300
rect 33000 559100 33200 559300
rect 33400 559100 33600 559300
rect 33800 559100 34000 559300
rect 34200 559100 34400 559300
rect 34600 559100 34800 559300
rect 35000 559100 35200 559300
rect 35400 559100 35600 559300
rect 35800 559100 36000 559300
rect 36200 559100 36400 559300
rect 36600 559100 36800 559300
rect 37000 559100 37200 559300
rect 37400 559100 37600 559300
rect 37800 559100 38000 559300
rect 38200 559100 38400 559300
rect 38600 559100 38800 559300
rect 39000 559100 39200 559300
rect 39400 559100 39600 559300
rect 39800 559100 40000 559300
rect 40200 559100 40400 559300
rect 40600 559100 40800 559300
rect 32600 558900 40800 559100
rect 32600 558700 32800 558900
rect 33000 558700 33200 558900
rect 33400 558700 33600 558900
rect 33800 558700 34000 558900
rect 34200 558700 34400 558900
rect 34600 558700 34800 558900
rect 35000 558700 35200 558900
rect 35400 558700 35600 558900
rect 35800 558700 36000 558900
rect 36200 558700 36400 558900
rect 36600 558700 36800 558900
rect 37000 558700 37200 558900
rect 37400 558700 37600 558900
rect 37800 558700 38000 558900
rect 38200 558700 38400 558900
rect 38600 558700 38800 558900
rect 39000 558700 39200 558900
rect 39400 558700 39600 558900
rect 39800 558700 40000 558900
rect 40200 558700 40400 558900
rect 40600 558700 40800 558900
rect 32600 558500 40800 558700
rect 32600 558300 32800 558500
rect 33000 558300 33200 558500
rect 33400 558300 33600 558500
rect 33800 558300 34000 558500
rect 34200 558300 34400 558500
rect 34600 558300 34800 558500
rect 35000 558300 35200 558500
rect 35400 558300 35600 558500
rect 35800 558300 36000 558500
rect 36200 558300 36400 558500
rect 36600 558300 36800 558500
rect 37000 558300 37200 558500
rect 37400 558300 37600 558500
rect 37800 558300 38000 558500
rect 38200 558300 38400 558500
rect 38600 558300 38800 558500
rect 39000 558300 39200 558500
rect 39400 558300 39600 558500
rect 39800 558300 40000 558500
rect 40200 558300 40400 558500
rect 40600 558300 40800 558500
rect 32600 558100 40800 558300
rect 32600 557900 32800 558100
rect 33000 557900 33200 558100
rect 33400 557900 33600 558100
rect 33800 557900 34000 558100
rect 34200 557900 34400 558100
rect 34600 557900 34800 558100
rect 35000 557900 35200 558100
rect 35400 557900 35600 558100
rect 35800 557900 36000 558100
rect 36200 557900 36400 558100
rect 36600 557900 36800 558100
rect 37000 557900 37200 558100
rect 37400 557900 37600 558100
rect 37800 557900 38000 558100
rect 38200 557900 38400 558100
rect 38600 557900 38800 558100
rect 39000 557900 39200 558100
rect 39400 557900 39600 558100
rect 39800 557900 40000 558100
rect 40200 557900 40400 558100
rect 40600 557900 40800 558100
rect 32600 557700 40800 557900
rect 32600 557500 32800 557700
rect 33000 557500 33200 557700
rect 33400 557500 33600 557700
rect 33800 557500 34000 557700
rect 34200 557500 34400 557700
rect 34600 557500 34800 557700
rect 35000 557500 35200 557700
rect 35400 557500 35600 557700
rect 35800 557500 36000 557700
rect 36200 557500 36400 557700
rect 36600 557500 36800 557700
rect 37000 557500 37200 557700
rect 37400 557500 37600 557700
rect 37800 557500 38000 557700
rect 38200 557500 38400 557700
rect 38600 557500 38800 557700
rect 39000 557500 39200 557700
rect 39400 557500 39600 557700
rect 39800 557500 40000 557700
rect 40200 557500 40400 557700
rect 40600 557500 40800 557700
rect 32600 557300 40800 557500
rect 32600 557100 32800 557300
rect 33000 557100 33200 557300
rect 33400 557100 33600 557300
rect 33800 557100 34000 557300
rect 34200 557100 34400 557300
rect 34600 557100 34800 557300
rect 35000 557100 35200 557300
rect 35400 557100 35600 557300
rect 35800 557100 36000 557300
rect 36200 557100 36400 557300
rect 36600 557100 36800 557300
rect 37000 557100 37200 557300
rect 37400 557100 37600 557300
rect 37800 557100 38000 557300
rect 38200 557100 38400 557300
rect 38600 557100 38800 557300
rect 39000 557100 39200 557300
rect 39400 557100 39600 557300
rect 39800 557100 40000 557300
rect 40200 557100 40400 557300
rect 40600 557100 40800 557300
rect 32600 556900 40800 557100
rect 32600 556700 32800 556900
rect 33000 556700 33200 556900
rect 33400 556700 33600 556900
rect 33800 556700 34000 556900
rect 34200 556700 34400 556900
rect 34600 556700 34800 556900
rect 35000 556700 35200 556900
rect 35400 556700 35600 556900
rect 35800 556700 36000 556900
rect 36200 556700 36400 556900
rect 36600 556700 36800 556900
rect 37000 556700 37200 556900
rect 37400 556700 37600 556900
rect 37800 556700 38000 556900
rect 38200 556700 38400 556900
rect 38600 556700 38800 556900
rect 39000 556700 39200 556900
rect 39400 556700 39600 556900
rect 39800 556700 40000 556900
rect 40200 556700 40400 556900
rect 40600 556700 40800 556900
rect 32600 556500 40800 556700
rect 32600 556300 32800 556500
rect 33000 556300 33200 556500
rect 33400 556300 33600 556500
rect 33800 556300 34000 556500
rect 34200 556300 34400 556500
rect 34600 556300 34800 556500
rect 35000 556300 35200 556500
rect 35400 556300 35600 556500
rect 35800 556300 36000 556500
rect 36200 556300 36400 556500
rect 36600 556300 36800 556500
rect 37000 556300 37200 556500
rect 37400 556300 37600 556500
rect 37800 556300 38000 556500
rect 38200 556300 38400 556500
rect 38600 556300 38800 556500
rect 39000 556300 39200 556500
rect 39400 556300 39600 556500
rect 39800 556300 40000 556500
rect 40200 556300 40400 556500
rect 40600 556300 40800 556500
rect 32600 556100 40800 556300
rect 32600 555900 32800 556100
rect 33000 555900 33200 556100
rect 33400 555900 33600 556100
rect 33800 555900 34000 556100
rect 34200 555900 34400 556100
rect 34600 555900 34800 556100
rect 35000 555900 35200 556100
rect 35400 555900 35600 556100
rect 35800 555900 36000 556100
rect 36200 555900 36400 556100
rect 36600 555900 36800 556100
rect 37000 555900 37200 556100
rect 37400 555900 37600 556100
rect 37800 555900 38000 556100
rect 38200 555900 38400 556100
rect 38600 555900 38800 556100
rect 39000 555900 39200 556100
rect 39400 555900 39600 556100
rect 39800 555900 40000 556100
rect 40200 555900 40400 556100
rect 40600 555900 40800 556100
rect 32600 555700 40800 555900
rect 32600 555500 32800 555700
rect 33000 555500 33200 555700
rect 33400 555500 33600 555700
rect 33800 555500 34000 555700
rect 34200 555500 34400 555700
rect 34600 555500 34800 555700
rect 35000 555500 35200 555700
rect 35400 555500 35600 555700
rect 35800 555500 36000 555700
rect 36200 555500 36400 555700
rect 36600 555500 36800 555700
rect 37000 555500 37200 555700
rect 37400 555500 37600 555700
rect 37800 555500 38000 555700
rect 38200 555500 38400 555700
rect 38600 555500 38800 555700
rect 39000 555500 39200 555700
rect 39400 555500 39600 555700
rect 39800 555500 40000 555700
rect 40200 555500 40400 555700
rect 40600 555500 40800 555700
rect 32600 555300 40800 555500
rect 32600 555100 32800 555300
rect 33000 555100 33200 555300
rect 33400 555100 33600 555300
rect 33800 555100 34000 555300
rect 34200 555100 34400 555300
rect 34600 555100 34800 555300
rect 35000 555100 35200 555300
rect 35400 555100 35600 555300
rect 35800 555100 36000 555300
rect 36200 555100 36400 555300
rect 36600 555100 36800 555300
rect 37000 555100 37200 555300
rect 37400 555100 37600 555300
rect 37800 555100 38000 555300
rect 38200 555100 38400 555300
rect 38600 555100 38800 555300
rect 39000 555100 39200 555300
rect 39400 555100 39600 555300
rect 39800 555100 40000 555300
rect 40200 555100 40400 555300
rect 40600 555100 40800 555300
rect 32600 554900 40800 555100
rect 32600 554700 32800 554900
rect 33000 554700 33200 554900
rect 33400 554700 33600 554900
rect 33800 554700 34000 554900
rect 34200 554700 34400 554900
rect 34600 554700 34800 554900
rect 35000 554700 35200 554900
rect 35400 554700 35600 554900
rect 35800 554700 36000 554900
rect 36200 554700 36400 554900
rect 36600 554700 36800 554900
rect 37000 554700 37200 554900
rect 37400 554700 37600 554900
rect 37800 554700 38000 554900
rect 38200 554700 38400 554900
rect 38600 554700 38800 554900
rect 39000 554700 39200 554900
rect 39400 554700 39600 554900
rect 39800 554700 40000 554900
rect 40200 554700 40400 554900
rect 40600 554700 40800 554900
rect 32600 554500 40800 554700
rect 32600 554300 32800 554500
rect 33000 554300 33200 554500
rect 33400 554300 33600 554500
rect 33800 554300 34000 554500
rect 34200 554300 34400 554500
rect 34600 554300 34800 554500
rect 35000 554300 35200 554500
rect 35400 554300 35600 554500
rect 35800 554300 36000 554500
rect 36200 554300 36400 554500
rect 36600 554300 36800 554500
rect 37000 554300 37200 554500
rect 37400 554300 37600 554500
rect 37800 554300 38000 554500
rect 38200 554300 38400 554500
rect 38600 554300 38800 554500
rect 39000 554300 39200 554500
rect 39400 554300 39600 554500
rect 39800 554300 40000 554500
rect 40200 554300 40400 554500
rect 40600 554300 40800 554500
rect 32600 554100 40800 554300
rect 32600 553900 32800 554100
rect 33000 553900 33200 554100
rect 33400 553900 33600 554100
rect 33800 553900 34000 554100
rect 34200 553900 34400 554100
rect 34600 553900 34800 554100
rect 35000 553900 35200 554100
rect 35400 553900 35600 554100
rect 35800 553900 36000 554100
rect 36200 553900 36400 554100
rect 36600 553900 36800 554100
rect 37000 553900 37200 554100
rect 37400 553900 37600 554100
rect 37800 553900 38000 554100
rect 38200 553900 38400 554100
rect 38600 553900 38800 554100
rect 39000 553900 39200 554100
rect 39400 553900 39600 554100
rect 39800 553900 40000 554100
rect 40200 553900 40400 554100
rect 40600 553900 40800 554100
rect 32600 553700 40800 553900
rect 32600 553500 32800 553700
rect 33000 553500 33200 553700
rect 33400 553500 33600 553700
rect 33800 553500 34000 553700
rect 34200 553500 34400 553700
rect 34600 553500 34800 553700
rect 35000 553500 35200 553700
rect 35400 553500 35600 553700
rect 35800 553500 36000 553700
rect 36200 553500 36400 553700
rect 36600 553500 36800 553700
rect 37000 553500 37200 553700
rect 37400 553500 37600 553700
rect 37800 553500 38000 553700
rect 38200 553500 38400 553700
rect 38600 553500 38800 553700
rect 39000 553500 39200 553700
rect 39400 553500 39600 553700
rect 39800 553500 40000 553700
rect 40200 553500 40400 553700
rect 40600 553500 40800 553700
rect 32600 553300 40800 553500
rect 32600 553100 32800 553300
rect 33000 553100 33200 553300
rect 33400 553100 33600 553300
rect 33800 553100 34000 553300
rect 34200 553100 34400 553300
rect 34600 553100 34800 553300
rect 35000 553100 35200 553300
rect 35400 553100 35600 553300
rect 35800 553100 36000 553300
rect 36200 553100 36400 553300
rect 36600 553100 36800 553300
rect 37000 553100 37200 553300
rect 37400 553100 37600 553300
rect 37800 553100 38000 553300
rect 38200 553100 38400 553300
rect 38600 553100 38800 553300
rect 39000 553100 39200 553300
rect 39400 553100 39600 553300
rect 39800 553100 40000 553300
rect 40200 553100 40400 553300
rect 40600 553100 40800 553300
rect 32600 552900 40800 553100
rect 32600 552700 32800 552900
rect 33000 552700 33200 552900
rect 33400 552700 33600 552900
rect 33800 552700 34000 552900
rect 34200 552700 34400 552900
rect 34600 552700 34800 552900
rect 35000 552700 35200 552900
rect 35400 552700 35600 552900
rect 35800 552700 36000 552900
rect 36200 552700 36400 552900
rect 36600 552700 36800 552900
rect 37000 552700 37200 552900
rect 37400 552700 37600 552900
rect 37800 552700 38000 552900
rect 38200 552700 38400 552900
rect 38600 552700 38800 552900
rect 39000 552700 39200 552900
rect 39400 552700 39600 552900
rect 39800 552700 40000 552900
rect 40200 552700 40400 552900
rect 40600 552700 40800 552900
rect 32600 552500 40800 552700
rect 32600 552300 32800 552500
rect 33000 552300 33200 552500
rect 33400 552300 33600 552500
rect 33800 552300 34000 552500
rect 34200 552300 34400 552500
rect 34600 552300 34800 552500
rect 35000 552300 35200 552500
rect 35400 552300 35600 552500
rect 35800 552300 36000 552500
rect 36200 552300 36400 552500
rect 36600 552300 36800 552500
rect 37000 552300 37200 552500
rect 37400 552300 37600 552500
rect 37800 552300 38000 552500
rect 38200 552300 38400 552500
rect 38600 552300 38800 552500
rect 39000 552300 39200 552500
rect 39400 552300 39600 552500
rect 39800 552300 40000 552500
rect 40200 552300 40400 552500
rect 40600 552300 40800 552500
rect 32600 552100 40800 552300
rect 32600 551900 32800 552100
rect 33000 551900 33200 552100
rect 33400 551900 33600 552100
rect 33800 551900 34000 552100
rect 34200 551900 34400 552100
rect 34600 551900 34800 552100
rect 35000 551900 35200 552100
rect 35400 551900 35600 552100
rect 35800 551900 36000 552100
rect 36200 551900 36400 552100
rect 36600 551900 36800 552100
rect 37000 551900 37200 552100
rect 37400 551900 37600 552100
rect 37800 551900 38000 552100
rect 38200 551900 38400 552100
rect 38600 551900 38800 552100
rect 39000 551900 39200 552100
rect 39400 551900 39600 552100
rect 39800 551900 40000 552100
rect 40200 551900 40400 552100
rect 40600 551900 40800 552100
rect 32600 551700 40800 551900
rect 32600 551500 32800 551700
rect 33000 551500 33200 551700
rect 33400 551500 33600 551700
rect 33800 551500 34000 551700
rect 34200 551500 34400 551700
rect 34600 551500 34800 551700
rect 35000 551500 35200 551700
rect 35400 551500 35600 551700
rect 35800 551500 36000 551700
rect 36200 551500 36400 551700
rect 36600 551500 36800 551700
rect 37000 551500 37200 551700
rect 37400 551500 37600 551700
rect 37800 551500 38000 551700
rect 38200 551500 38400 551700
rect 38600 551500 38800 551700
rect 39000 551500 39200 551700
rect 39400 551500 39600 551700
rect 39800 551500 40000 551700
rect 40200 551500 40400 551700
rect 40600 551500 40800 551700
rect 32600 551300 40800 551500
rect 32600 551100 32800 551300
rect 33000 551100 33200 551300
rect 33400 551100 33600 551300
rect 33800 551100 34000 551300
rect 34200 551100 34400 551300
rect 34600 551100 34800 551300
rect 35000 551100 35200 551300
rect 35400 551100 35600 551300
rect 35800 551100 36000 551300
rect 36200 551100 36400 551300
rect 36600 551100 36800 551300
rect 37000 551100 37200 551300
rect 37400 551100 37600 551300
rect 37800 551100 38000 551300
rect 38200 551100 38400 551300
rect 38600 551100 38800 551300
rect 39000 551100 39200 551300
rect 39400 551100 39600 551300
rect 39800 551100 40000 551300
rect 40200 551100 40400 551300
rect 40600 551100 40800 551300
rect 32600 550900 40800 551100
rect 32600 550700 32800 550900
rect 33000 550700 33200 550900
rect 33400 550700 33600 550900
rect 33800 550700 34000 550900
rect 34200 550700 34400 550900
rect 34600 550700 34800 550900
rect 35000 550700 35200 550900
rect 35400 550700 35600 550900
rect 35800 550700 36000 550900
rect 36200 550700 36400 550900
rect 36600 550700 36800 550900
rect 37000 550700 37200 550900
rect 37400 550700 37600 550900
rect 37800 550700 38000 550900
rect 38200 550700 38400 550900
rect 38600 550700 38800 550900
rect 39000 550700 39200 550900
rect 39400 550700 39600 550900
rect 39800 550700 40000 550900
rect 40200 550700 40400 550900
rect 40600 550700 40800 550900
rect 32600 550500 40800 550700
rect 32600 550300 32800 550500
rect 33000 550300 33200 550500
rect 33400 550300 33600 550500
rect 33800 550300 34000 550500
rect 34200 550300 34400 550500
rect 34600 550300 34800 550500
rect 35000 550300 35200 550500
rect 35400 550300 35600 550500
rect 35800 550300 36000 550500
rect 36200 550300 36400 550500
rect 36600 550300 36800 550500
rect 37000 550300 37200 550500
rect 37400 550300 37600 550500
rect 37800 550300 38000 550500
rect 38200 550300 38400 550500
rect 38600 550300 38800 550500
rect 39000 550300 39200 550500
rect 39400 550300 39600 550500
rect 39800 550300 40000 550500
rect 40200 550300 40400 550500
rect 40600 550300 40800 550500
rect 32600 550100 40800 550300
rect 32600 549900 32800 550100
rect 33000 549900 33200 550100
rect 33400 549900 33600 550100
rect 33800 549900 34000 550100
rect 34200 549900 34400 550100
rect 34600 549900 34800 550100
rect 35000 549900 35200 550100
rect 35400 549900 35600 550100
rect 35800 549900 36000 550100
rect 36200 549900 36400 550100
rect 36600 549900 36800 550100
rect 37000 549900 37200 550100
rect 37400 549900 37600 550100
rect 37800 549900 38000 550100
rect 38200 549900 38400 550100
rect 38600 549900 38800 550100
rect 39000 549900 39200 550100
rect 39400 549900 39600 550100
rect 39800 549900 40000 550100
rect 40200 549900 40400 550100
rect 40600 549900 40800 550100
rect 32600 549700 40800 549900
rect 32600 549500 32800 549700
rect 33000 549500 33200 549700
rect 33400 549500 33600 549700
rect 33800 549500 34000 549700
rect 34200 549500 34400 549700
rect 34600 549500 34800 549700
rect 35000 549500 35200 549700
rect 35400 549500 35600 549700
rect 35800 549500 36000 549700
rect 36200 549500 36400 549700
rect 36600 549500 36800 549700
rect 37000 549500 37200 549700
rect 37400 549500 37600 549700
rect 37800 549500 38000 549700
rect 38200 549500 38400 549700
rect 38600 549500 38800 549700
rect 39000 549500 39200 549700
rect 39400 549500 39600 549700
rect 39800 549500 40000 549700
rect 40200 549500 40400 549700
rect 40600 549500 40800 549700
rect 32600 549400 40800 549500
<< rmetal4 >>
rect 515500 697940 521000 698500
<< via4 >>
rect 12900 673800 13200 674100
rect 13700 673800 14000 674100
rect 12900 673300 13200 673600
rect 13700 673300 14000 673600
rect 12900 672800 13200 673100
rect 13700 672800 14000 673100
rect 2500 648300 2800 648600
rect 3000 648300 3300 648600
rect 3500 648300 3800 648600
rect 23400 648200 23700 648500
rect 24100 648200 24400 648500
rect 2500 647800 2800 648100
rect 3000 647800 3300 648100
rect 3500 647800 3800 648100
rect 2500 647300 2800 647600
rect 3000 647300 3300 647600
rect 3500 647300 3800 647600
rect 23400 647600 23700 647900
rect 24100 647600 24400 647900
rect 2500 646800 2800 647100
rect 3000 646800 3300 647100
rect 3500 646800 3800 647100
rect 23400 647000 23700 647300
rect 24100 647000 24400 647300
rect 2500 646300 2800 646600
rect 3000 646300 3300 646600
rect 3500 646300 3800 646600
rect 23400 646300 23700 646600
rect 24100 646300 24400 646600
rect 2500 645800 2800 646100
rect 3000 645800 3300 646100
rect 3500 645800 3800 646100
rect 23400 645700 23700 646000
rect 24100 645700 24400 646000
rect 2500 645300 2800 645600
rect 3000 645300 3300 645600
rect 3500 645300 3800 645600
rect 2500 644800 2800 645100
rect 3000 644800 3300 645100
rect 3500 644800 3800 645100
rect 23400 645100 23700 645400
rect 24100 645100 24400 645400
rect 2500 644300 2800 644600
rect 3000 644300 3300 644600
rect 3500 644300 3800 644600
rect 23400 644500 23700 644800
rect 24100 644500 24400 644800
rect 2500 643800 2800 644100
rect 3000 643800 3300 644100
rect 3500 643800 3800 644100
rect 23400 643900 23700 644200
rect 24100 643900 24400 644200
rect 2500 643300 2800 643600
rect 3000 643300 3300 643600
rect 3500 643300 3800 643600
rect 23400 643300 23700 643600
rect 24100 643300 24400 643600
rect 2500 642800 2800 643100
rect 3000 642800 3300 643100
rect 3500 642800 3800 643100
rect 2500 642300 2800 642600
rect 3000 642300 3300 642600
rect 3500 642300 3800 642600
rect 23400 642600 23700 642900
rect 24100 642600 24400 642900
rect 2500 641800 2800 642100
rect 3000 641800 3300 642100
rect 3500 641800 3800 642100
rect 23400 642000 23700 642300
rect 24100 642000 24400 642300
rect 2500 641300 2800 641600
rect 3000 641300 3300 641600
rect 3500 641300 3800 641600
rect 23400 641400 23700 641700
rect 24100 641400 24400 641700
rect 2500 640800 2800 641100
rect 3000 640800 3300 641100
rect 3500 640800 3800 641100
rect 23400 640800 23700 641100
rect 24100 640800 24400 641100
rect 2500 640300 2800 640600
rect 3000 640300 3300 640600
rect 3500 640300 3800 640600
rect 23400 640200 23700 640500
rect 24100 640200 24400 640500
rect 2500 639800 2800 640100
rect 3000 639800 3300 640100
rect 3500 639800 3800 640100
rect 2500 639300 2800 639600
rect 3000 639300 3300 639600
rect 3500 639300 3800 639600
rect 23400 639600 23700 639900
rect 24100 639600 24400 639900
rect 2500 638800 2800 639100
rect 3000 638800 3300 639100
rect 3500 638800 3800 639100
rect 23400 639000 23700 639300
rect 24100 639000 24400 639300
rect 2500 638300 2800 638600
rect 3000 638300 3300 638600
rect 3500 638300 3800 638600
rect 23400 638400 23700 638700
rect 24100 638400 24400 638700
rect 2500 637800 2800 638100
rect 3000 637800 3300 638100
rect 3500 637800 3800 638100
rect 23400 637800 23700 638100
rect 24100 637800 24400 638100
rect 2500 637300 2800 637600
rect 3000 637300 3300 637600
rect 3500 637300 3800 637600
rect 2500 636800 2800 637100
rect 3000 636800 3300 637100
rect 3500 636800 3800 637100
rect 23400 637100 23700 637400
rect 24100 637100 24400 637400
rect 2500 636300 2800 636600
rect 3000 636300 3300 636600
rect 3500 636300 3800 636600
rect 23400 636400 23700 636700
rect 24100 636400 24400 636700
rect 2500 635800 2800 636100
rect 3000 635800 3300 636100
rect 3500 635800 3800 636100
rect 23400 635700 23700 636000
rect 24100 635700 24400 636000
rect 2500 635300 2800 635600
rect 3000 635300 3300 635600
rect 3500 635300 3800 635600
rect 2500 634800 2800 635100
rect 3000 634800 3300 635100
rect 3500 634800 3800 635100
rect 23400 634900 23700 635200
rect 24100 634900 24400 635200
rect 2500 634300 2800 634600
rect 3000 634300 3300 634600
rect 3500 634300 3800 634600
rect 23400 634200 23700 634500
rect 24100 634200 24400 634500
rect 32800 673700 33100 674000
rect 33300 673700 33600 674000
rect 33800 673700 34100 674000
rect 34300 673700 34600 674000
rect 34800 673700 35100 674000
rect 35300 673700 35600 674000
rect 35800 673700 36100 674000
rect 36300 673700 36600 674000
rect 36800 673700 37100 674000
rect 37300 673700 37600 674000
rect 37800 673700 38100 674000
rect 38300 673700 38600 674000
rect 38800 673700 39100 674000
rect 39300 673700 39600 674000
rect 39800 673700 40100 674000
rect 40300 673700 40600 674000
rect 32800 672900 33100 673200
rect 33300 672900 33600 673200
rect 33800 672900 34100 673200
rect 34300 672900 34600 673200
rect 34800 672900 35100 673200
rect 35300 672900 35600 673200
rect 35800 672900 36100 673200
rect 36300 672900 36600 673200
rect 36800 672900 37100 673200
rect 37300 672900 37600 673200
rect 37800 672900 38100 673200
rect 38300 672900 38600 673200
rect 38800 672900 39100 673200
rect 39300 672900 39600 673200
rect 39800 672900 40100 673200
rect 40300 672900 40600 673200
rect 50100 673700 50400 674000
rect 50100 673300 50400 673600
rect 50100 672900 50400 673200
rect 32800 670400 33100 670700
rect 33300 670400 33600 670700
rect 33800 670400 34100 670700
rect 34300 670400 34600 670700
rect 34800 670400 35100 670700
rect 35300 670400 35600 670700
rect 35800 670400 36100 670700
rect 36300 670400 36600 670700
rect 36800 670400 37100 670700
rect 37300 670400 37600 670700
rect 37800 670400 38100 670700
rect 38300 670400 38600 670700
rect 38800 670400 39100 670700
rect 39300 670400 39600 670700
rect 39800 670400 40100 670700
rect 40300 670400 40600 670700
rect 32800 669700 33100 670000
rect 33300 669700 33600 670000
rect 33800 669700 34100 670000
rect 34300 669700 34600 670000
rect 34800 669700 35100 670000
rect 35300 669700 35600 670000
rect 35800 669700 36100 670000
rect 36300 669700 36600 670000
rect 36800 669700 37100 670000
rect 37300 669700 37600 670000
rect 37800 669700 38100 670000
rect 38300 669700 38600 670000
rect 38800 669700 39100 670000
rect 39300 669700 39600 670000
rect 39800 669700 40100 670000
rect 40300 669700 40600 670000
rect 32800 667100 33100 667400
rect 33300 667100 33600 667400
rect 33800 667100 34100 667400
rect 34300 667100 34600 667400
rect 34800 667100 35100 667400
rect 35300 667100 35600 667400
rect 35800 667100 36100 667400
rect 36300 667100 36600 667400
rect 36800 667100 37100 667400
rect 37300 667100 37600 667400
rect 37800 667100 38100 667400
rect 38300 667100 38600 667400
rect 38800 667100 39100 667400
rect 39300 667100 39600 667400
rect 39800 667100 40100 667400
rect 40300 667100 40600 667400
rect 32800 666400 33100 666700
rect 33300 666400 33600 666700
rect 33800 666400 34100 666700
rect 34300 666400 34600 666700
rect 34800 666400 35100 666700
rect 35300 666400 35600 666700
rect 35800 666400 36100 666700
rect 36300 666400 36600 666700
rect 36800 666400 37100 666700
rect 37300 666400 37600 666700
rect 37800 666400 38100 666700
rect 38300 666400 38600 666700
rect 38800 666400 39100 666700
rect 39300 666400 39600 666700
rect 39800 666400 40100 666700
rect 40300 666400 40600 666700
rect 549900 684600 550200 684900
rect 550400 684600 550700 684900
rect 550900 684600 551200 684900
rect 551400 684600 551700 684900
rect 551900 684600 552200 684900
rect 552400 684600 552700 684900
rect 549900 684100 550200 684400
rect 550400 684100 550700 684400
rect 550900 684100 551200 684400
rect 551400 684100 551700 684400
rect 551900 684100 552200 684400
rect 552400 684100 552700 684400
rect 549900 683600 550200 683900
rect 550400 683600 550700 683900
rect 550900 683600 551200 683900
rect 551400 683600 551700 683900
rect 551900 683600 552200 683900
rect 552400 683600 552700 683900
rect 573200 684600 573500 684900
rect 573800 684600 574100 684900
rect 573200 684100 573500 684400
rect 573800 684100 574100 684400
rect 576800 684400 577100 684700
rect 577300 684400 577600 684700
rect 577800 684400 578100 684700
rect 578300 684400 578600 684700
rect 573200 683600 573500 683900
rect 573800 683600 574100 683900
rect 576800 683900 577100 684200
rect 577300 683900 577600 684200
rect 577800 683900 578100 684200
rect 578300 683900 578600 684200
rect 58000 648300 58300 648600
rect 58500 648300 58800 648600
rect 59000 648300 59300 648600
rect 59500 648300 59800 648600
rect 60000 648300 60300 648600
rect 60500 648300 60800 648600
rect 61000 648300 61300 648600
rect 61500 648300 61800 648600
rect 58000 647800 58300 648100
rect 58500 647800 58800 648100
rect 59000 647800 59300 648100
rect 59500 647800 59800 648100
rect 60000 647800 60300 648100
rect 60500 647800 60800 648100
rect 61000 647800 61300 648100
rect 61500 647800 61800 648100
rect 58000 647300 58300 647600
rect 58500 647300 58800 647600
rect 59000 647300 59300 647600
rect 59500 647300 59800 647600
rect 60000 647300 60300 647600
rect 60500 647300 60800 647600
rect 61000 647300 61300 647600
rect 61500 647300 61800 647600
rect 58000 646800 58300 647100
rect 58500 646800 58800 647100
rect 59000 646800 59300 647100
rect 59500 646800 59800 647100
rect 60000 646800 60300 647100
rect 60500 646800 60800 647100
rect 61000 646800 61300 647100
rect 61500 646800 61800 647100
rect 58000 646300 58300 646600
rect 58500 646300 58800 646600
rect 59000 646300 59300 646600
rect 59500 646300 59800 646600
rect 60000 646300 60300 646600
rect 60500 646300 60800 646600
rect 61000 646300 61300 646600
rect 61500 646300 61800 646600
rect 58000 645800 58300 646100
rect 58500 645800 58800 646100
rect 59000 645800 59300 646100
rect 59500 645800 59800 646100
rect 60000 645800 60300 646100
rect 60500 645800 60800 646100
rect 61000 645800 61300 646100
rect 61500 645800 61800 646100
rect 58000 645300 58300 645600
rect 58500 645300 58800 645600
rect 59000 645300 59300 645600
rect 59500 645300 59800 645600
rect 60000 645300 60300 645600
rect 60500 645300 60800 645600
rect 61000 645300 61300 645600
rect 61500 645300 61800 645600
rect 58000 644800 58300 645100
rect 58500 644800 58800 645100
rect 59000 644800 59300 645100
rect 59500 644800 59800 645100
rect 60000 644800 60300 645100
rect 60500 644800 60800 645100
rect 61000 644800 61300 645100
rect 61500 644800 61800 645100
rect 58000 644300 58300 644600
rect 58500 644300 58800 644600
rect 59000 644300 59300 644600
rect 59500 644300 59800 644600
rect 60000 644300 60300 644600
rect 60500 644300 60800 644600
rect 61000 644300 61300 644600
rect 61500 644300 61800 644600
rect 58000 643800 58300 644100
rect 58500 643800 58800 644100
rect 59000 643800 59300 644100
rect 59500 643800 59800 644100
rect 60000 643800 60300 644100
rect 60500 643800 60800 644100
rect 61000 643800 61300 644100
rect 61500 643800 61800 644100
rect 58000 643300 58300 643600
rect 58500 643300 58800 643600
rect 59000 643300 59300 643600
rect 59500 643300 59800 643600
rect 60000 643300 60300 643600
rect 60500 643300 60800 643600
rect 61000 643300 61300 643600
rect 61500 643300 61800 643600
rect 58000 642800 58300 643100
rect 58500 642800 58800 643100
rect 59000 642800 59300 643100
rect 59500 642800 59800 643100
rect 60000 642800 60300 643100
rect 60500 642800 60800 643100
rect 61000 642800 61300 643100
rect 61500 642800 61800 643100
rect 58000 642300 58300 642600
rect 58500 642300 58800 642600
rect 59000 642300 59300 642600
rect 59500 642300 59800 642600
rect 60000 642300 60300 642600
rect 60500 642300 60800 642600
rect 61000 642300 61300 642600
rect 61500 642300 61800 642600
rect 58000 641800 58300 642100
rect 58500 641800 58800 642100
rect 59000 641800 59300 642100
rect 59500 641800 59800 642100
rect 60000 641800 60300 642100
rect 60500 641800 60800 642100
rect 61000 641800 61300 642100
rect 61500 641800 61800 642100
rect 58000 641300 58300 641600
rect 58500 641300 58800 641600
rect 59000 641300 59300 641600
rect 59500 641300 59800 641600
rect 60000 641300 60300 641600
rect 60500 641300 60800 641600
rect 61000 641300 61300 641600
rect 61500 641300 61800 641600
rect 58000 640800 58300 641100
rect 58500 640800 58800 641100
rect 59000 640800 59300 641100
rect 59500 640800 59800 641100
rect 60000 640800 60300 641100
rect 60500 640800 60800 641100
rect 61000 640800 61300 641100
rect 61500 640800 61800 641100
rect 58000 640300 58300 640600
rect 58500 640300 58800 640600
rect 59000 640300 59300 640600
rect 59500 640300 59800 640600
rect 60000 640300 60300 640600
rect 60500 640300 60800 640600
rect 61000 640300 61300 640600
rect 61500 640300 61800 640600
rect 58000 639800 58300 640100
rect 58500 639800 58800 640100
rect 59000 639800 59300 640100
rect 59500 639800 59800 640100
rect 60000 639800 60300 640100
rect 60500 639800 60800 640100
rect 61000 639800 61300 640100
rect 61500 639800 61800 640100
rect 58000 639300 58300 639600
rect 58500 639300 58800 639600
rect 59000 639300 59300 639600
rect 59500 639300 59800 639600
rect 60000 639300 60300 639600
rect 60500 639300 60800 639600
rect 61000 639300 61300 639600
rect 61500 639300 61800 639600
rect 58000 638800 58300 639100
rect 58500 638800 58800 639100
rect 59000 638800 59300 639100
rect 59500 638800 59800 639100
rect 60000 638800 60300 639100
rect 60500 638800 60800 639100
rect 61000 638800 61300 639100
rect 61500 638800 61800 639100
rect 58000 638300 58300 638600
rect 58500 638300 58800 638600
rect 59000 638300 59300 638600
rect 59500 638300 59800 638600
rect 60000 638300 60300 638600
rect 60500 638300 60800 638600
rect 61000 638300 61300 638600
rect 61500 638300 61800 638600
rect 58000 637800 58300 638100
rect 58500 637800 58800 638100
rect 59000 637800 59300 638100
rect 59500 637800 59800 638100
rect 60000 637800 60300 638100
rect 60500 637800 60800 638100
rect 61000 637800 61300 638100
rect 61500 637800 61800 638100
rect 58000 637300 58300 637600
rect 58500 637300 58800 637600
rect 59000 637300 59300 637600
rect 59500 637300 59800 637600
rect 60000 637300 60300 637600
rect 60500 637300 60800 637600
rect 61000 637300 61300 637600
rect 61500 637300 61800 637600
rect 58000 636800 58300 637100
rect 58500 636800 58800 637100
rect 59000 636800 59300 637100
rect 59500 636800 59800 637100
rect 60000 636800 60300 637100
rect 60500 636800 60800 637100
rect 61000 636800 61300 637100
rect 61500 636800 61800 637100
rect 58000 636300 58300 636600
rect 58500 636300 58800 636600
rect 59000 636300 59300 636600
rect 59500 636300 59800 636600
rect 60000 636300 60300 636600
rect 60500 636300 60800 636600
rect 61000 636300 61300 636600
rect 61500 636300 61800 636600
rect 58000 635800 58300 636100
rect 58500 635800 58800 636100
rect 59000 635800 59300 636100
rect 59500 635800 59800 636100
rect 60000 635800 60300 636100
rect 60500 635800 60800 636100
rect 61000 635800 61300 636100
rect 61500 635800 61800 636100
rect 58000 635300 58300 635600
rect 58500 635300 58800 635600
rect 59000 635300 59300 635600
rect 59500 635300 59800 635600
rect 60000 635300 60300 635600
rect 60500 635300 60800 635600
rect 61000 635300 61300 635600
rect 61500 635300 61800 635600
rect 58000 634800 58300 635100
rect 58500 634800 58800 635100
rect 59000 634800 59300 635100
rect 59500 634800 59800 635100
rect 60000 634800 60300 635100
rect 60500 634800 60800 635100
rect 61000 634800 61300 635100
rect 61500 634800 61800 635100
rect 58000 634300 58300 634600
rect 58500 634300 58800 634600
rect 59000 634300 59300 634600
rect 59500 634300 59800 634600
rect 60000 634300 60300 634600
rect 60500 634300 60800 634600
rect 61000 634300 61300 634600
rect 61500 634300 61800 634600
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 549700 684900 578640 685100
rect 549700 684600 549900 684900
rect 550200 684600 550400 684900
rect 550700 684600 550900 684900
rect 551200 684600 551400 684900
rect 551700 684600 551900 684900
rect 552200 684600 552400 684900
rect 552700 684600 573200 684900
rect 573500 684600 573800 684900
rect 574100 684700 578640 684900
rect 574100 684600 576800 684700
rect 549700 684400 576800 684600
rect 577100 684400 577300 684700
rect 577600 684400 577800 684700
rect 578100 684400 578300 684700
rect 578600 684400 578640 684700
rect 549700 684100 549900 684400
rect 550200 684100 550400 684400
rect 550700 684100 550900 684400
rect 551200 684100 551400 684400
rect 551700 684100 551900 684400
rect 552200 684100 552400 684400
rect 552700 684100 573200 684400
rect 573500 684100 573800 684400
rect 574100 684200 578640 684400
rect 574100 684100 576800 684200
rect 549700 683900 576800 684100
rect 577100 683900 577300 684200
rect 577600 683900 577800 684200
rect 578100 683900 578300 684200
rect 578600 683900 578640 684200
rect 549700 683600 549900 683900
rect 550200 683600 550400 683900
rect 550700 683600 550900 683900
rect 551200 683600 551400 683900
rect 551700 683600 551900 683900
rect 552200 683600 552400 683900
rect 552700 683600 573200 683900
rect 573500 683600 573800 683900
rect 574100 683600 578640 683900
rect 549700 683400 578640 683600
rect 12800 674100 51300 674200
rect 12800 673800 12900 674100
rect 13200 673800 13700 674100
rect 14000 674000 51300 674100
rect 14000 673800 32800 674000
rect 12800 673700 32800 673800
rect 33100 673700 33300 674000
rect 33600 673700 33800 674000
rect 34100 673700 34300 674000
rect 34600 673700 34800 674000
rect 35100 673700 35300 674000
rect 35600 673700 35800 674000
rect 36100 673700 36300 674000
rect 36600 673700 36800 674000
rect 37100 673700 37300 674000
rect 37600 673700 37800 674000
rect 38100 673700 38300 674000
rect 38600 673700 38800 674000
rect 39100 673700 39300 674000
rect 39600 673700 39800 674000
rect 40100 673700 40300 674000
rect 40600 673700 50100 674000
rect 50400 673700 51300 674000
rect 12800 673600 51300 673700
rect 12800 673300 12900 673600
rect 13200 673300 13700 673600
rect 14000 673300 50100 673600
rect 50400 673300 51300 673600
rect 12800 673200 51300 673300
rect 12800 673100 32800 673200
rect 12800 672800 12900 673100
rect 13200 672800 13700 673100
rect 14000 672900 32800 673100
rect 33100 672900 33300 673200
rect 33600 672900 33800 673200
rect 34100 672900 34300 673200
rect 34600 672900 34800 673200
rect 35100 672900 35300 673200
rect 35600 672900 35800 673200
rect 36100 672900 36300 673200
rect 36600 672900 36800 673200
rect 37100 672900 37300 673200
rect 37600 672900 37800 673200
rect 38100 672900 38300 673200
rect 38600 672900 38800 673200
rect 39100 672900 39300 673200
rect 39600 672900 39800 673200
rect 40100 672900 40300 673200
rect 40600 672900 50100 673200
rect 50400 672900 51300 673200
rect 14000 672800 51300 672900
rect 12800 672700 51300 672800
rect 32600 670700 48300 670900
rect 32600 670400 32800 670700
rect 33100 670400 33300 670700
rect 33600 670400 33800 670700
rect 34100 670400 34300 670700
rect 34600 670400 34800 670700
rect 35100 670400 35300 670700
rect 35600 670400 35800 670700
rect 36100 670400 36300 670700
rect 36600 670400 36800 670700
rect 37100 670400 37300 670700
rect 37600 670400 37800 670700
rect 38100 670400 38300 670700
rect 38600 670400 38800 670700
rect 39100 670400 39300 670700
rect 39600 670400 39800 670700
rect 40100 670400 40300 670700
rect 40600 670400 48300 670700
rect 32600 670000 48300 670400
rect 32600 669700 32800 670000
rect 33100 669700 33300 670000
rect 33600 669700 33800 670000
rect 34100 669700 34300 670000
rect 34600 669700 34800 670000
rect 35100 669700 35300 670000
rect 35600 669700 35800 670000
rect 36100 669700 36300 670000
rect 36600 669700 36800 670000
rect 37100 669700 37300 670000
rect 37600 669700 37800 670000
rect 38100 669700 38300 670000
rect 38600 669700 38800 670000
rect 39100 669700 39300 670000
rect 39600 669700 39800 670000
rect 40100 669700 40300 670000
rect 40600 669700 48300 670000
rect 32600 669500 48300 669700
rect 32600 667400 48300 667600
rect 32600 667100 32800 667400
rect 33100 667100 33300 667400
rect 33600 667100 33800 667400
rect 34100 667100 34300 667400
rect 34600 667100 34800 667400
rect 35100 667100 35300 667400
rect 35600 667100 35800 667400
rect 36100 667100 36300 667400
rect 36600 667100 36800 667400
rect 37100 667100 37300 667400
rect 37600 667100 37800 667400
rect 38100 667100 38300 667400
rect 38600 667100 38800 667400
rect 39100 667100 39300 667400
rect 39600 667100 39800 667400
rect 40100 667100 40300 667400
rect 40600 667100 48300 667400
rect 32600 666700 48300 667100
rect 32600 666400 32800 666700
rect 33100 666400 33300 666700
rect 33600 666400 33800 666700
rect 34100 666400 34300 666700
rect 34600 666400 34800 666700
rect 35100 666400 35300 666700
rect 35600 666400 35800 666700
rect 36100 666400 36300 666700
rect 36600 666400 36800 666700
rect 37100 666400 37300 666700
rect 37600 666400 37800 666700
rect 38100 666400 38300 666700
rect 38600 666400 38800 666700
rect 39100 666400 39300 666700
rect 39600 666400 39800 666700
rect 40100 666400 40300 666700
rect 40600 666400 48300 666700
rect 32600 666200 48300 666400
rect 2300 648600 62200 648800
rect 2300 648300 2500 648600
rect 2800 648300 3000 648600
rect 3300 648300 3500 648600
rect 3800 648500 58000 648600
rect 3800 648300 23400 648500
rect 2300 648200 23400 648300
rect 23700 648200 24100 648500
rect 24400 648300 58000 648500
rect 58300 648300 58500 648600
rect 58800 648300 59000 648600
rect 59300 648300 59500 648600
rect 59800 648300 60000 648600
rect 60300 648300 60500 648600
rect 60800 648300 61000 648600
rect 61300 648300 61500 648600
rect 61800 648300 62200 648600
rect 24400 648200 62200 648300
rect 2300 648100 62200 648200
rect 2300 647800 2500 648100
rect 2800 647800 3000 648100
rect 3300 647800 3500 648100
rect 3800 647900 58000 648100
rect 3800 647800 23400 647900
rect 2300 647600 23400 647800
rect 23700 647600 24100 647900
rect 24400 647800 58000 647900
rect 58300 647800 58500 648100
rect 58800 647800 59000 648100
rect 59300 647800 59500 648100
rect 59800 647800 60000 648100
rect 60300 647800 60500 648100
rect 60800 647800 61000 648100
rect 61300 647800 61500 648100
rect 61800 647800 62200 648100
rect 24400 647600 62200 647800
rect 2300 647300 2500 647600
rect 2800 647300 3000 647600
rect 3300 647300 3500 647600
rect 3800 647300 58000 647600
rect 58300 647300 58500 647600
rect 58800 647300 59000 647600
rect 59300 647300 59500 647600
rect 59800 647300 60000 647600
rect 60300 647300 60500 647600
rect 60800 647300 61000 647600
rect 61300 647300 61500 647600
rect 61800 647300 62200 647600
rect 2300 647100 23400 647300
rect 2300 646800 2500 647100
rect 2800 646800 3000 647100
rect 3300 646800 3500 647100
rect 3800 647000 23400 647100
rect 23700 647000 24100 647300
rect 24400 647100 62200 647300
rect 24400 647000 58000 647100
rect 3800 646800 58000 647000
rect 58300 646800 58500 647100
rect 58800 646800 59000 647100
rect 59300 646800 59500 647100
rect 59800 646800 60000 647100
rect 60300 646800 60500 647100
rect 60800 646800 61000 647100
rect 61300 646800 61500 647100
rect 61800 646800 62200 647100
rect 2300 646600 62200 646800
rect 2300 646300 2500 646600
rect 2800 646300 3000 646600
rect 3300 646300 3500 646600
rect 3800 646300 23400 646600
rect 23700 646300 24100 646600
rect 24400 646300 58000 646600
rect 58300 646300 58500 646600
rect 58800 646300 59000 646600
rect 59300 646300 59500 646600
rect 59800 646300 60000 646600
rect 60300 646300 60500 646600
rect 60800 646300 61000 646600
rect 61300 646300 61500 646600
rect 61800 646300 62200 646600
rect 2300 646100 62200 646300
rect 2300 645800 2500 646100
rect 2800 645800 3000 646100
rect 3300 645800 3500 646100
rect 3800 646000 58000 646100
rect 3800 645800 23400 646000
rect 2300 645700 23400 645800
rect 23700 645700 24100 646000
rect 24400 645800 58000 646000
rect 58300 645800 58500 646100
rect 58800 645800 59000 646100
rect 59300 645800 59500 646100
rect 59800 645800 60000 646100
rect 60300 645800 60500 646100
rect 60800 645800 61000 646100
rect 61300 645800 61500 646100
rect 61800 645800 62200 646100
rect 24400 645700 62200 645800
rect 2300 645600 62200 645700
rect 2300 645300 2500 645600
rect 2800 645300 3000 645600
rect 3300 645300 3500 645600
rect 3800 645400 58000 645600
rect 3800 645300 23400 645400
rect 2300 645100 23400 645300
rect 23700 645100 24100 645400
rect 24400 645300 58000 645400
rect 58300 645300 58500 645600
rect 58800 645300 59000 645600
rect 59300 645300 59500 645600
rect 59800 645300 60000 645600
rect 60300 645300 60500 645600
rect 60800 645300 61000 645600
rect 61300 645300 61500 645600
rect 61800 645300 62200 645600
rect 24400 645100 62200 645300
rect 2300 644800 2500 645100
rect 2800 644800 3000 645100
rect 3300 644800 3500 645100
rect 3800 644800 58000 645100
rect 58300 644800 58500 645100
rect 58800 644800 59000 645100
rect 59300 644800 59500 645100
rect 59800 644800 60000 645100
rect 60300 644800 60500 645100
rect 60800 644800 61000 645100
rect 61300 644800 61500 645100
rect 61800 644800 62200 645100
rect 2300 644600 23400 644800
rect 2300 644300 2500 644600
rect 2800 644300 3000 644600
rect 3300 644300 3500 644600
rect 3800 644500 23400 644600
rect 23700 644500 24100 644800
rect 24400 644600 62200 644800
rect 24400 644500 58000 644600
rect 3800 644300 58000 644500
rect 58300 644300 58500 644600
rect 58800 644300 59000 644600
rect 59300 644300 59500 644600
rect 59800 644300 60000 644600
rect 60300 644300 60500 644600
rect 60800 644300 61000 644600
rect 61300 644300 61500 644600
rect 61800 644300 62200 644600
rect 2300 644200 62200 644300
rect 2300 644100 23400 644200
rect 2300 643800 2500 644100
rect 2800 643800 3000 644100
rect 3300 643800 3500 644100
rect 3800 643900 23400 644100
rect 23700 643900 24100 644200
rect 24400 644100 62200 644200
rect 24400 643900 58000 644100
rect 3800 643800 58000 643900
rect 58300 643800 58500 644100
rect 58800 643800 59000 644100
rect 59300 643800 59500 644100
rect 59800 643800 60000 644100
rect 60300 643800 60500 644100
rect 60800 643800 61000 644100
rect 61300 643800 61500 644100
rect 61800 643800 62200 644100
rect 2300 643600 62200 643800
rect 2300 643300 2500 643600
rect 2800 643300 3000 643600
rect 3300 643300 3500 643600
rect 3800 643300 23400 643600
rect 23700 643300 24100 643600
rect 24400 643300 58000 643600
rect 58300 643300 58500 643600
rect 58800 643300 59000 643600
rect 59300 643300 59500 643600
rect 59800 643300 60000 643600
rect 60300 643300 60500 643600
rect 60800 643300 61000 643600
rect 61300 643300 61500 643600
rect 61800 643300 62200 643600
rect 2300 643100 62200 643300
rect 2300 642800 2500 643100
rect 2800 642800 3000 643100
rect 3300 642800 3500 643100
rect 3800 642900 58000 643100
rect 3800 642800 23400 642900
rect 2300 642600 23400 642800
rect 23700 642600 24100 642900
rect 24400 642800 58000 642900
rect 58300 642800 58500 643100
rect 58800 642800 59000 643100
rect 59300 642800 59500 643100
rect 59800 642800 60000 643100
rect 60300 642800 60500 643100
rect 60800 642800 61000 643100
rect 61300 642800 61500 643100
rect 61800 642800 62200 643100
rect 24400 642600 62200 642800
rect 2300 642300 2500 642600
rect 2800 642300 3000 642600
rect 3300 642300 3500 642600
rect 3800 642300 58000 642600
rect 58300 642300 58500 642600
rect 58800 642300 59000 642600
rect 59300 642300 59500 642600
rect 59800 642300 60000 642600
rect 60300 642300 60500 642600
rect 60800 642300 61000 642600
rect 61300 642300 61500 642600
rect 61800 642300 62200 642600
rect 2300 642100 23400 642300
rect 2300 641800 2500 642100
rect 2800 641800 3000 642100
rect 3300 641800 3500 642100
rect 3800 642000 23400 642100
rect 23700 642000 24100 642300
rect 24400 642100 62200 642300
rect 24400 642000 58000 642100
rect 3800 641800 58000 642000
rect 58300 641800 58500 642100
rect 58800 641800 59000 642100
rect 59300 641800 59500 642100
rect 59800 641800 60000 642100
rect 60300 641800 60500 642100
rect 60800 641800 61000 642100
rect 61300 641800 61500 642100
rect 61800 641800 62200 642100
rect 2300 641700 62200 641800
rect 2300 641600 23400 641700
rect 2300 641300 2500 641600
rect 2800 641300 3000 641600
rect 3300 641300 3500 641600
rect 3800 641400 23400 641600
rect 23700 641400 24100 641700
rect 24400 641600 62200 641700
rect 24400 641400 58000 641600
rect 3800 641300 58000 641400
rect 58300 641300 58500 641600
rect 58800 641300 59000 641600
rect 59300 641300 59500 641600
rect 59800 641300 60000 641600
rect 60300 641300 60500 641600
rect 60800 641300 61000 641600
rect 61300 641300 61500 641600
rect 61800 641300 62200 641600
rect 2300 641100 62200 641300
rect 2300 640800 2500 641100
rect 2800 640800 3000 641100
rect 3300 640800 3500 641100
rect 3800 640800 23400 641100
rect 23700 640800 24100 641100
rect 24400 640800 58000 641100
rect 58300 640800 58500 641100
rect 58800 640800 59000 641100
rect 59300 640800 59500 641100
rect 59800 640800 60000 641100
rect 60300 640800 60500 641100
rect 60800 640800 61000 641100
rect 61300 640800 61500 641100
rect 61800 640800 62200 641100
rect 2300 640600 62200 640800
rect 2300 640300 2500 640600
rect 2800 640300 3000 640600
rect 3300 640300 3500 640600
rect 3800 640500 58000 640600
rect 3800 640300 23400 640500
rect 2300 640200 23400 640300
rect 23700 640200 24100 640500
rect 24400 640300 58000 640500
rect 58300 640300 58500 640600
rect 58800 640300 59000 640600
rect 59300 640300 59500 640600
rect 59800 640300 60000 640600
rect 60300 640300 60500 640600
rect 60800 640300 61000 640600
rect 61300 640300 61500 640600
rect 61800 640300 62200 640600
rect 24400 640200 62200 640300
rect 2300 640100 62200 640200
rect 2300 639800 2500 640100
rect 2800 639800 3000 640100
rect 3300 639800 3500 640100
rect 3800 639900 58000 640100
rect 3800 639800 23400 639900
rect 2300 639600 23400 639800
rect 23700 639600 24100 639900
rect 24400 639800 58000 639900
rect 58300 639800 58500 640100
rect 58800 639800 59000 640100
rect 59300 639800 59500 640100
rect 59800 639800 60000 640100
rect 60300 639800 60500 640100
rect 60800 639800 61000 640100
rect 61300 639800 61500 640100
rect 61800 639800 62200 640100
rect 24400 639600 62200 639800
rect 2300 639300 2500 639600
rect 2800 639300 3000 639600
rect 3300 639300 3500 639600
rect 3800 639300 58000 639600
rect 58300 639300 58500 639600
rect 58800 639300 59000 639600
rect 59300 639300 59500 639600
rect 59800 639300 60000 639600
rect 60300 639300 60500 639600
rect 60800 639300 61000 639600
rect 61300 639300 61500 639600
rect 61800 639300 62200 639600
rect 2300 639100 23400 639300
rect 2300 638800 2500 639100
rect 2800 638800 3000 639100
rect 3300 638800 3500 639100
rect 3800 639000 23400 639100
rect 23700 639000 24100 639300
rect 24400 639100 62200 639300
rect 24400 639000 58000 639100
rect 3800 638800 58000 639000
rect 58300 638800 58500 639100
rect 58800 638800 59000 639100
rect 59300 638800 59500 639100
rect 59800 638800 60000 639100
rect 60300 638800 60500 639100
rect 60800 638800 61000 639100
rect 61300 638800 61500 639100
rect 61800 638800 62200 639100
rect 2300 638700 62200 638800
rect 2300 638600 23400 638700
rect 2300 638300 2500 638600
rect 2800 638300 3000 638600
rect 3300 638300 3500 638600
rect 3800 638400 23400 638600
rect 23700 638400 24100 638700
rect 24400 638600 62200 638700
rect 24400 638400 58000 638600
rect 3800 638300 58000 638400
rect 58300 638300 58500 638600
rect 58800 638300 59000 638600
rect 59300 638300 59500 638600
rect 59800 638300 60000 638600
rect 60300 638300 60500 638600
rect 60800 638300 61000 638600
rect 61300 638300 61500 638600
rect 61800 638300 62200 638600
rect 2300 638100 62200 638300
rect 2300 637800 2500 638100
rect 2800 637800 3000 638100
rect 3300 637800 3500 638100
rect 3800 637800 23400 638100
rect 23700 637800 24100 638100
rect 24400 637800 58000 638100
rect 58300 637800 58500 638100
rect 58800 637800 59000 638100
rect 59300 637800 59500 638100
rect 59800 637800 60000 638100
rect 60300 637800 60500 638100
rect 60800 637800 61000 638100
rect 61300 637800 61500 638100
rect 61800 637800 62200 638100
rect 2300 637600 62200 637800
rect 2300 637300 2500 637600
rect 2800 637300 3000 637600
rect 3300 637300 3500 637600
rect 3800 637400 58000 637600
rect 3800 637300 23400 637400
rect 2300 637100 23400 637300
rect 23700 637100 24100 637400
rect 24400 637300 58000 637400
rect 58300 637300 58500 637600
rect 58800 637300 59000 637600
rect 59300 637300 59500 637600
rect 59800 637300 60000 637600
rect 60300 637300 60500 637600
rect 60800 637300 61000 637600
rect 61300 637300 61500 637600
rect 61800 637300 62200 637600
rect 24400 637100 62200 637300
rect 2300 636800 2500 637100
rect 2800 636800 3000 637100
rect 3300 636800 3500 637100
rect 3800 636800 58000 637100
rect 58300 636800 58500 637100
rect 58800 636800 59000 637100
rect 59300 636800 59500 637100
rect 59800 636800 60000 637100
rect 60300 636800 60500 637100
rect 60800 636800 61000 637100
rect 61300 636800 61500 637100
rect 61800 636800 62200 637100
rect 2300 636700 62200 636800
rect 2300 636600 23400 636700
rect 2300 636300 2500 636600
rect 2800 636300 3000 636600
rect 3300 636300 3500 636600
rect 3800 636400 23400 636600
rect 23700 636400 24100 636700
rect 24400 636600 62200 636700
rect 24400 636400 58000 636600
rect 3800 636300 58000 636400
rect 58300 636300 58500 636600
rect 58800 636300 59000 636600
rect 59300 636300 59500 636600
rect 59800 636300 60000 636600
rect 60300 636300 60500 636600
rect 60800 636300 61000 636600
rect 61300 636300 61500 636600
rect 61800 636300 62200 636600
rect 2300 636100 62200 636300
rect 2300 635800 2500 636100
rect 2800 635800 3000 636100
rect 3300 635800 3500 636100
rect 3800 636000 58000 636100
rect 3800 635800 23400 636000
rect 2300 635700 23400 635800
rect 23700 635700 24100 636000
rect 24400 635800 58000 636000
rect 58300 635800 58500 636100
rect 58800 635800 59000 636100
rect 59300 635800 59500 636100
rect 59800 635800 60000 636100
rect 60300 635800 60500 636100
rect 60800 635800 61000 636100
rect 61300 635800 61500 636100
rect 61800 635800 62200 636100
rect 24400 635700 62200 635800
rect 2300 635600 62200 635700
rect 2300 635300 2500 635600
rect 2800 635300 3000 635600
rect 3300 635300 3500 635600
rect 3800 635300 58000 635600
rect 58300 635300 58500 635600
rect 58800 635300 59000 635600
rect 59300 635300 59500 635600
rect 59800 635300 60000 635600
rect 60300 635300 60500 635600
rect 60800 635300 61000 635600
rect 61300 635300 61500 635600
rect 61800 635300 62200 635600
rect 2300 635200 62200 635300
rect 2300 635100 23400 635200
rect 2300 634800 2500 635100
rect 2800 634800 3000 635100
rect 3300 634800 3500 635100
rect 3800 634900 23400 635100
rect 23700 634900 24100 635200
rect 24400 635100 62200 635200
rect 24400 634900 58000 635100
rect 3800 634800 58000 634900
rect 58300 634800 58500 635100
rect 58800 634800 59000 635100
rect 59300 634800 59500 635100
rect 59800 634800 60000 635100
rect 60300 634800 60500 635100
rect 60800 634800 61000 635100
rect 61300 634800 61500 635100
rect 61800 634800 62200 635100
rect 2300 634600 62200 634800
rect 2300 634300 2500 634600
rect 2800 634300 3000 634600
rect 3300 634300 3500 634600
rect 3800 634500 58000 634600
rect 3800 634300 23400 634500
rect 2300 634200 23400 634300
rect 23700 634200 24100 634500
rect 24400 634300 58000 634500
rect 58300 634300 58500 634600
rect 58800 634300 59000 634600
rect 59300 634300 59500 634600
rect 59800 634300 60000 634600
rect 60300 634300 60500 634600
rect 60800 634300 61000 634600
rect 61300 634300 61500 634600
rect 61800 634300 62200 634600
rect 24400 634200 62200 634300
rect 2300 633800 62200 634200
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use OTA_MULT_GM  OTA_MULT_GM_0
timestamp 1683391037
transform 1 0 544600 0 1 677936
box -10044 -14658 10212 17116
use OTA_fingers_031123_NON_FLAT  OTA_fingers_031123_NON_FLAT_0
timestamp 1683391037
transform 1 0 42740 0 1 684710
box -5940 -310 9780 16550
use constant_gm_fingers  constant_gm_fingers_0
timestamp 1683407140
transform 1 0 43810 0 1 682900
box -2700 -20100 4420 1140
use diode_connected_nmos  diode_connected_nmos_0
timestamp 1683391037
transform 1 0 23260 0 1 691860
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_1
timestamp 1683391037
transform 1 0 12860 0 1 691860
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_2
timestamp 1683391037
transform 1 0 75260 0 1 691860
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_3
timestamp 1683391037
transform 1 0 64860 0 1 691860
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_4
timestamp 1683391037
transform 1 0 563860 0 1 691660
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_5
timestamp 1683391037
transform 1 0 573060 0 1 691660
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_6
timestamp 1683391037
transform 0 1 572140 -1 0 684834
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_7
timestamp 1683391037
transform 0 1 572160 -1 0 677354
box -60 -60 1254 10360
<< labels >>
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
